-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Aug 25 2019 21:32:08

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    USBPU : out std_logic;
    PIN_9 : in std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : in std_logic;
    PIN_5 : in std_logic;
    PIN_4 : in std_logic;
    PIN_3 : out std_logic;
    PIN_24 : in std_logic;
    PIN_23 : in std_logic;
    PIN_22 : in std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : in std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : in std_logic;
    PIN_10 : in std_logic;
    PIN_1 : out std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17357\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \CLK_ibuf_gb_io_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \PIN_2_c\ : std_logic;
signal \c0.rx.r_Rx_Data_RZ0\ : std_logic;
signal \c0.rx.rx_data_ready\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_c2_cascade_\ : std_logic;
signal \c0.rx.g0_i_o4_0_1_cascade_\ : std_logic;
signal \c0.rx.g0_i_o2_2_3_cascade_\ : std_logic;
signal \c0.rx.g0_i_a4_1_1\ : std_logic;
signal \PIN_1_c\ : std_logic;
signal \c0.rx.un1_r_Rx_DV7_0\ : std_logic;
signal \c0.rx.g0_i_o2_5\ : std_logic;
signal \c0.rx.g0_i_o2_4\ : std_logic;
signal \c0.rx.g0_i_o2_6\ : std_logic;
signal \c0.rx.g0_i_a4_1_3\ : std_logic;
signal \c0.rx.N_7_cascade_\ : std_logic;
signal \c0.rx.r_SM_Main_RNICMJF6_0Z0Z_1\ : std_logic;
signal \c0.rx.N_10_0\ : std_logic;
signal \c0.rx.N_13_0\ : std_logic;
signal \c0.rx.N_12_1_cascade_\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_c2\ : std_logic;
signal \c0.rx.N_6_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count_2_sqmuxa_0\ : std_logic;
signal \c0.rx.r_Clock_Count_2_sqmuxa_0_cascade_\ : std_logic;
signal \c0.rx.g1_4\ : std_logic;
signal \c0.rx.g1_5_cascade_\ : std_logic;
signal \c0.rx.g1\ : std_logic;
signal \c0.rx.g0_0_1_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count14_cascade_\ : std_logic;
signal \c0.rx.m6_ns_1\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_m_0_cascade_\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_2_sqmuxa_0\ : std_logic;
signal \c0.rx.r_Clock_Count_1_sqmuxa_0\ : std_logic;
signal \c0.rx.un1_r_Clock_Count_5_m_1_cascade_\ : std_logic;
signal \N_12\ : std_logic;
signal \N_8_0\ : std_logic;
signal \LED_c\ : std_logic;
signal \c0.rx.CO1_cascade_\ : std_logic;
signal \c0.rx.g0_i_o3_0_4_cascade_\ : std_logic;
signal \c0.rx.N_10\ : std_logic;
signal \c0.rx.N_12_0\ : std_logic;
signal \c0.rx.N_9_0_cascade_\ : std_logic;
signal \c0.rx.N_11_i\ : std_logic;
signal \c0.rx.r_Clock_CountZ0Z_6\ : std_logic;
signal \c0.rx.r_Clock_CountZ0Z_5\ : std_logic;
signal \c0.rx.r_Clock_CountZ0Z_7\ : std_logic;
signal \c0.rx.r_Clock_CountZ0Z_4\ : std_logic;
signal \c0.rx.r_Clock_Count14_3_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count26_cascade_\ : std_logic;
signal \c0.rx.r_Clock_CountZ0Z_2\ : std_logic;
signal \c0.rx.r_Clock_CountZ0Z_3\ : std_logic;
signal \c0.rx.g0_i_a4_0_3_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count14_3\ : std_logic;
signal \c0.rx.N_13\ : std_logic;
signal \c0.rx.r_Clock_Count26\ : std_logic;
signal \c0.rx.r_SM_MainZ0Z_2\ : std_logic;
signal \c0.rx.r_Rx_DV_1_sqmuxa_cascade_\ : std_logic;
signal \c0.rx.r_SM_MainZ0Z_1\ : std_logic;
signal \c0.rx.r_SM_MainZ0Z_0\ : std_logic;
signal \c0.rx.r_Clock_Count14\ : std_logic;
signal \c0.rx.N_9\ : std_logic;
signal \c0.rx.r_Clock_CountZ0Z_0\ : std_logic;
signal \c0.rx.r_Clock_CountZ0Z_1\ : std_logic;
signal \c0.rx.r_Clock_Count14_1\ : std_logic;
signal \bfn_5_25_0_\ : std_logic;
signal \c0.tx.un1_r_Clock_Count_cry_0\ : std_logic;
signal \c0.tx.r_Clock_Count_RNO_0Z0Z_2\ : std_logic;
signal \c0.tx.un1_r_Clock_Count_cry_1\ : std_logic;
signal \c0.tx.un1_r_Clock_Count_cry_2\ : std_logic;
signal \c0.tx.r_Clock_Count_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \c0.tx.r_Clock_Count_RNO_0Z0Z_0\ : std_logic;
signal \c0.tx.r_Clock_CountZ0Z_0\ : std_logic;
signal \c0.tx.r_Clock_Count_0_sqmuxa\ : std_logic;
signal \c0.tx.r_Clock_Count_RNO_0Z0Z_1\ : std_logic;
signal \blink_counterZ0Z_0\ : std_logic;
signal \bfn_6_20_0_\ : std_logic;
signal \blink_counterZ0Z_1\ : std_logic;
signal blink_counter_cry_0 : std_logic;
signal \blink_counterZ0Z_2\ : std_logic;
signal blink_counter_cry_1 : std_logic;
signal \blink_counterZ0Z_3\ : std_logic;
signal blink_counter_cry_2 : std_logic;
signal \blink_counterZ0Z_4\ : std_logic;
signal blink_counter_cry_3 : std_logic;
signal \blink_counterZ0Z_5\ : std_logic;
signal blink_counter_cry_4 : std_logic;
signal \blink_counterZ0Z_6\ : std_logic;
signal blink_counter_cry_5 : std_logic;
signal \blink_counterZ0Z_7\ : std_logic;
signal blink_counter_cry_6 : std_logic;
signal blink_counter_cry_7 : std_logic;
signal \blink_counterZ0Z_8\ : std_logic;
signal \bfn_6_21_0_\ : std_logic;
signal \blink_counterZ0Z_9\ : std_logic;
signal blink_counter_cry_8 : std_logic;
signal \blink_counterZ0Z_10\ : std_logic;
signal blink_counter_cry_9 : std_logic;
signal \blink_counterZ0Z_11\ : std_logic;
signal blink_counter_cry_10 : std_logic;
signal \blink_counterZ0Z_12\ : std_logic;
signal blink_counter_cry_11 : std_logic;
signal \blink_counterZ0Z_13\ : std_logic;
signal blink_counter_cry_12 : std_logic;
signal \blink_counterZ0Z_14\ : std_logic;
signal blink_counter_cry_13 : std_logic;
signal \blink_counterZ0Z_15\ : std_logic;
signal blink_counter_cry_14 : std_logic;
signal blink_counter_cry_15 : std_logic;
signal \blink_counterZ0Z_16\ : std_logic;
signal \bfn_6_22_0_\ : std_logic;
signal \blink_counterZ0Z_17\ : std_logic;
signal blink_counter_cry_16 : std_logic;
signal \blink_counterZ0Z_18\ : std_logic;
signal blink_counter_cry_17 : std_logic;
signal \blink_counterZ0Z_19\ : std_logic;
signal blink_counter_cry_18 : std_logic;
signal \blink_counterZ0Z_20\ : std_logic;
signal blink_counter_cry_19 : std_logic;
signal \blink_counterZ0Z_21\ : std_logic;
signal blink_counter_cry_20 : std_logic;
signal \blink_counterZ0Z_22\ : std_logic;
signal blink_counter_cry_21 : std_logic;
signal \blink_counterZ0Z_23\ : std_logic;
signal blink_counter_cry_22 : std_logic;
signal blink_counter_cry_23 : std_logic;
signal \blink_counterZ0Z_24\ : std_logic;
signal \bfn_6_23_0_\ : std_logic;
signal blink_counter_cry_24 : std_logic;
signal \blink_counterZ0Z_25\ : std_logic;
signal \c0.tx.N_287_cascade_\ : std_logic;
signal \c0.tx.N_294\ : std_logic;
signal \c0.tx.o_Tx_Serial12\ : std_logic;
signal \c0.tx.N_294_cascade_\ : std_logic;
signal \c0.tx.m5_0_0\ : std_logic;
signal \c0.tx.N_287\ : std_logic;
signal \c0.tx.N_288_cascade_\ : std_logic;
signal \c0.tx.r_Clock_Count_i_0\ : std_logic;
signal \bfn_6_25_0_\ : std_logic;
signal \c0.tx.r_Clock_CountZ0Z_1\ : std_logic;
signal \c0.tx.r_Clock_Count_i_1\ : std_logic;
signal \c0.tx.r_Clock_Count12_cry_0\ : std_logic;
signal \c0.tx.r_Clock_CountZ0Z_2\ : std_logic;
signal \c0.tx.r_Clock_Count_i_2\ : std_logic;
signal \c0.tx.r_Clock_Count12_cry_1\ : std_logic;
signal \c0.tx.r_Clock_CountZ0Z_3\ : std_logic;
signal \c0.tx.r_Clock_Count_i_3\ : std_logic;
signal \c0.tx.r_Clock_Count12_cry_2\ : std_logic;
signal \c0.tx.r_Clock_Count12\ : std_logic;
signal \c0.rx.r_Rx_Bytece_1_1_cascade_\ : std_logic;
signal \c0.rx.r_Rx_Bytece_1_5\ : std_logic;
signal \c0.rx.r_Rx_DV6\ : std_logic;
signal \c0.tx.r_Tx_Active_1_sqmuxa_cascade_\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_1\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_1\ : std_logic;
signal \c0.tx.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_3_cascade_\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_3\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_5\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_5\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_3\ : std_logic;
signal \c0.tx.r_Bit_IndexZ0Z_2\ : std_logic;
signal \c0.tx.r_Bit_IndexZ0Z_1\ : std_logic;
signal \c0.tx.r_Tx_Data_pmux_3_i_m2_ns_1_cascade_\ : std_logic;
signal \c0.tx.N_354\ : std_logic;
signal \c0.tx.r_Bit_IndexZ0Z_0\ : std_logic;
signal \c0.tx.N_357_cascade_\ : std_logic;
signal \c0.tx.N_320\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_5_cascade_\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_5\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_0\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_4\ : std_logic;
signal \c0.data_out_7_Z0Z_5\ : std_logic;
signal \c0.rx.r_Rx_Bytece_0_3_cascade_\ : std_logic;
signal \c0.rx_data_3\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_2_cascade_\ : std_logic;
signal \c0.tx.r_SM_MainZ0Z_0\ : std_logic;
signal \c0.tx.r_SM_MainZ0Z_1\ : std_logic;
signal \c0.tx.r_Clock_Count12_THRU_CO\ : std_logic;
signal \c0.tx.r_SM_MainZ0Z_2\ : std_logic;
signal \c0.nextCRC16_3_3_12_cascade_\ : std_logic;
signal \c0.nextCRC16_3_4_12\ : std_logic;
signal \c0.data_out_6_Z0Z_4\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_4\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_1_cascade_\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_1\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_3\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_11_cascade_\ : std_logic;
signal \c0.data_out_6_Z0Z_3\ : std_logic;
signal \c0.d_2_7\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_7_cascade_\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_7\ : std_logic;
signal \c0.N_74\ : std_logic;
signal \c0.N_74_cascade_\ : std_logic;
signal \c0.d_2_19\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \c0.dataZ0Z_1\ : std_logic;
signal \c0.data_cry_0\ : std_logic;
signal \c0.data_cry_1\ : std_logic;
signal \c0.data_cry_2\ : std_logic;
signal \c0.data_cry_3\ : std_logic;
signal \c0.data_cry_4\ : std_logic;
signal \c0.data_cry_5\ : std_logic;
signal \c0.data_cry_6\ : std_logic;
signal \c0.data_cry_7\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \c0.data_cry_8\ : std_logic;
signal \c0.data_cry_9\ : std_logic;
signal \c0.dataZ0Z_11\ : std_logic;
signal \c0.data_cry_10\ : std_logic;
signal \c0.dataZ0Z_12\ : std_logic;
signal \c0.data_cry_11\ : std_logic;
signal \c0.data_cry_12\ : std_logic;
signal \c0.dataZ0Z_14\ : std_logic;
signal \c0.data_cry_13\ : std_logic;
signal \c0.data_cry_14\ : std_logic;
signal \c0.i12_0_and\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \c0.i12_0\ : std_logic;
signal \c0.i12_2_and\ : std_logic;
signal \c0.i12_1\ : std_logic;
signal \c0.i12_2\ : std_logic;
signal \c0.i12_3\ : std_logic;
signal \c0.i12_5_and\ : std_logic;
signal \c0.i12_4\ : std_logic;
signal \c0.i12_5\ : std_logic;
signal \c0.i12_6\ : std_logic;
signal \c0.i12\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \c0.i12_1_and\ : std_logic;
signal \c0.i12_3_and\ : std_logic;
signal \c0.i12_4_and\ : std_logic;
signal \c0.i12_6_and\ : std_logic;
signal \c0.rx_data_5\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_2\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_2\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \c0.tx2_data_1_0_i_ns_1_2\ : std_logic;
signal \c0.tx2_data_1_iv_4_3\ : std_logic;
signal \c0.rx.un1_r_Rx_Byte_7\ : std_logic;
signal \c0.tx2.o_Tx_Serial12_cascade_\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_3\ : std_logic;
signal \c0.d_2_38\ : std_logic;
signal \c0.m115_amcf1\ : std_logic;
signal \c0.N_293_cascade_\ : std_logic;
signal \c0.tx_data_1_0_i_1_6\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_6\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_2\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_7\ : std_logic;
signal \c0.tx.r_Tx_DataZ0Z_7\ : std_logic;
signal \c0.tx.r_Tx_Data_0_sqmuxa\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_4\ : std_logic;
signal \c0.data_out_6_Z0Z_1\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_5\ : std_logic;
signal \c0.d_2_23\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_7\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_1\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_2\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_15_cascade_\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_4_cascade_\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_4\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_4\ : std_logic;
signal \c0.data_out_7_Z0Z_4\ : std_logic;
signal \c0.dataZ0Z_7\ : std_logic;
signal \c0.dataZ0Z_3\ : std_logic;
signal \c0.dataZ0Z_10\ : std_logic;
signal \c0.dataZ0Z_6\ : std_logic;
signal \c0.dataZ0Z_2\ : std_logic;
signal \c0.data_out_7_Z0Z_2\ : std_logic;
signal \c0.dataZ0Z_5\ : std_logic;
signal \c0.dataZ0Z_13\ : std_logic;
signal \c0.d_2_37\ : std_logic;
signal \c0.dataZ0Z_4\ : std_logic;
signal \c0.dataZ0Z_9\ : std_logic;
signal \c0.i12_7_and\ : std_logic;
signal \c0.g1_1_cascade_\ : std_logic;
signal \c0.N_72_mux\ : std_logic;
signal \c0.N_249_cascade_\ : std_logic;
signal \c0.data_in_4_Z0Z_0\ : std_logic;
signal \c0.g1_cascade_\ : std_logic;
signal \c0.g0_3\ : std_logic;
signal \c0.byte_transmit_counter2_0_sqmuxa_0\ : std_logic;
signal \c0.g3_2_0_cascade_\ : std_logic;
signal \c0.g0_2\ : std_logic;
signal \c0.rx_data_1\ : std_logic;
signal \c0.data_in_3_Z0Z_4\ : std_logic;
signal \c0.data_in_1_Z0Z_6\ : std_logic;
signal \c0.data_in_3_Z0Z_5\ : std_logic;
signal \c0.data_in_5_Z0Z_2\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \c0.tx2.un1_r_Clock_Count_cry_0\ : std_logic;
signal \c0.tx2.r_Clock_Count_RNO_0_0_2\ : std_logic;
signal \c0.tx2.un1_r_Clock_Count_cry_1\ : std_logic;
signal \c0.tx2.un1_r_Clock_Count_cry_2\ : std_logic;
signal \c0.tx2.r_Clock_Count_RNO_0_0_3\ : std_logic;
signal \c0.tx2.r_Clock_Count_0_sqmuxa\ : std_logic;
signal \c0.tx2.r_Clock_Count_RNO_0_0_0\ : std_logic;
signal \c0.tx2.r_Clock_CountZ0Z_0\ : std_logic;
signal \c0.tx2.r_Clock_Count_RNO_0_0_1\ : std_logic;
signal \c0.tx2.r_Clock_Count_i_0\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \c0.tx2.r_Clock_CountZ0Z_1\ : std_logic;
signal \c0.tx2.r_Clock_Count_i_1\ : std_logic;
signal \c0.tx2.r_Clock_Count12_cry_0\ : std_logic;
signal \c0.tx2.r_Clock_CountZ0Z_2\ : std_logic;
signal \c0.tx2.r_Clock_Count_i_2\ : std_logic;
signal \c0.tx2.r_Clock_Count12_cry_1\ : std_logic;
signal \c0.tx2.r_Clock_CountZ0Z_3\ : std_logic;
signal \c0.tx2.r_Clock_Count_i_3\ : std_logic;
signal \c0.tx2.r_Clock_Count12_cry_2\ : std_logic;
signal \c0.tx2.r_Clock_Count12\ : std_logic;
signal \c0.N_76\ : std_logic;
signal \c0.data_out_6_Z0Z_2\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_2\ : std_logic;
signal \c0.d_2_21\ : std_logic;
signal \c0.tx_data_1_iv_i_m2_0_ns_1_0_cascade_\ : std_logic;
signal \c0.N_304_cascade_\ : std_logic;
signal \c0.tx_data_1_iv_i_1_0\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_8\ : std_logic;
signal \c0.N_77\ : std_logic;
signal \c0.data_out_6_Z0Z_0\ : std_logic;
signal \c0.dataZ0Z_0\ : std_logic;
signal \c0.data_out_7_Z0Z_0\ : std_logic;
signal \c0.d_2_8\ : std_logic;
signal \c0.tx_data_RNO_0Z0Z_0\ : std_logic;
signal \c0.N_93\ : std_logic;
signal \c0.nextCRC16_3_0_a2_0_10\ : std_logic;
signal \c0.d_2_22\ : std_logic;
signal \c0.d_2_6\ : std_logic;
signal \c0.nextCRC16_3_9\ : std_logic;
signal \c0.nextCRC16_3_0_a2_6_0_15_cascade_\ : std_logic;
signal \c0.N_92\ : std_logic;
signal \c0.d_2_41\ : std_logic;
signal \c0.d_2_12\ : std_logic;
signal \c0.d_2_40\ : std_logic;
signal \c0.nextCRC16_3_0_a2_2_2\ : std_logic;
signal \c0.d_2_3\ : std_logic;
signal \c0.N_75\ : std_logic;
signal \c0.N_75_cascade_\ : std_logic;
signal \c0.d_2_44\ : std_logic;
signal \c0.N_95\ : std_logic;
signal \c0.d_2_14\ : std_logic;
signal \c0.N_95_cascade_\ : std_logic;
signal \c0.d_2_25\ : std_logic;
signal \c0.d_2_11\ : std_logic;
signal \c0.dataZ0Z_8\ : std_logic;
signal \c0.dataZ0Z_15\ : std_logic;
signal \c0.tx2_active\ : std_logic;
signal \c0.tx2_data_1_iv_5_1_0_7\ : std_logic;
signal \c0.tx2_data_1_iv_5_1_7_cascade_\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_7\ : std_logic;
signal \c0.tx2_data_1_iv_3_1_3\ : std_logic;
signal \c0.tx2_data_1_iv_3_3\ : std_logic;
signal \c0.data_in_0_Z0Z_3\ : std_logic;
signal \c0.N_247_0\ : std_logic;
signal \c0.un1_data_in_6__0_0_a2_5_a2_2_cascade_\ : std_logic;
signal \c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_\ : std_logic;
signal \c0.un1_data_in_7__4_i_cascade_\ : std_logic;
signal \c0.un1_data_in_6__0\ : std_logic;
signal \c0.d_4_RNIF73E2Z0Z_14_cascade_\ : std_logic;
signal \c0.d_4_RNIMKFE3Z0Z_14_cascade_\ : std_logic;
signal \c0.un1_data_in_6__7_cascade_\ : std_logic;
signal \c0.wait_for_transmission4_12\ : std_logic;
signal \c0.data_in_frame_0__0_sqmuxa\ : std_logic;
signal \c0.wait_for_transmission4_12_cascade_\ : std_logic;
signal \c0.un1_data_in_7__4_0_a2_0_a2_4\ : std_logic;
signal \c0.data_in_0_Z0Z_2\ : std_logic;
signal \c0.d_4_RNID6K21_0Z0Z_15\ : std_logic;
signal \c0.d_4_RNID6K21Z0Z_15\ : std_logic;
signal \c0.data_in_0_Z0Z_1\ : std_logic;
signal \c0.data_in_1_Z0Z_7\ : std_logic;
signal \c0.data_in_3_Z0Z_7\ : std_logic;
signal \c0.un1_data_in_7__1_0_a2_24_a2_2_cascade_\ : std_logic;
signal \c0.d_4_2\ : std_logic;
signal \c0.N_103\ : std_logic;
signal \c0.wait_for_transmission4_13_1_1\ : std_logic;
signal \c0.un1_data_in_7__1_0_a2_24_a2_6_cascade_\ : std_logic;
signal \c0.un1_data_in_7__1_0_a2_24_a2_1_cascade_\ : std_logic;
signal \c0.un1_data_in_7__1_0_a2_24_a2_5\ : std_logic;
signal \c0.d_4_RNITCRCZ0Z_29\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_0_cascade_\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_0\ : std_logic;
signal \c0.tx2_data_1_0_i_ns_1_0_cascade_\ : std_logic;
signal \c0.d_4_1\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_1_cascade_\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_1\ : std_logic;
signal \c0.tx2_data_1_0_i_ns_1_1_cascade_\ : std_logic;
signal \c0.tx2_data_RNO_0Z0Z_1\ : std_logic;
signal \c0.tx2_data_RNO_4Z0Z_1\ : std_logic;
signal \c0.tx2_data_RNO_1Z0Z_0\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_2\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_0\ : std_logic;
signal \c0.tx2.r_Tx_Data_pmux_3_i_m2_ns_1\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_1\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_3\ : std_logic;
signal \c0.tx2.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_\ : std_logic;
signal \c0.tx2.N_349\ : std_logic;
signal \c0.tx2.N_346_cascade_\ : std_logic;
signal \c0.tx2.N_279_cascade_\ : std_logic;
signal \PIN_3_c\ : std_logic;
signal \c0.tx2.r_Tx_Active_1_sqmuxa\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_1\ : std_logic;
signal \c0.tx2.m5_0_0_cascade_\ : std_logic;
signal \c0.d_2_9\ : std_logic;
signal \c0.N_94\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_5\ : std_logic;
signal \c0.d_2_45\ : std_logic;
signal \c0.nextCRC16_3_0_a2_0_0\ : std_logic;
signal \c0.nextCRC16_3_0_a2_4_0\ : std_logic;
signal \c0.d_2_28\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_2\ : std_logic;
signal \c0.d_2_0\ : std_logic;
signal \c0.nextCRC16_3_4_0\ : std_logic;
signal \c0.d_2_13\ : std_logic;
signal \c0.d_2_26\ : std_logic;
signal \c0.nextCRC16_3_4_0_cascade_\ : std_logic;
signal \c0.N_99\ : std_logic;
signal \c0.nextCRC16_3_0_a2_3_0\ : std_logic;
signal \c0.d_2_39\ : std_logic;
signal \c0.data_out_6_Z0Z_5\ : std_logic;
signal \c0.nextCRC16_3_0_a2_4_15\ : std_logic;
signal \c0.nextCRC16_3_0_a2_3_15\ : std_logic;
signal \c0.data_out_6_Z0Z_7\ : std_logic;
signal \c0.d_2_16\ : std_logic;
signal \c0.d_2_24\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \c0.N_105\ : std_logic;
signal \c0.nextCRC16_3_2_1\ : std_logic;
signal \c0.N_106\ : std_logic;
signal \c0.data_out_7_Z0Z_1\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_5\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_7\ : std_logic;
signal \c0.wait_for_transmission_RNOZ0Z_10_cascade_\ : std_logic;
signal \c0.g0_5_4\ : std_logic;
signal \c0.d_4_3\ : std_logic;
signal \c0.d_4_45\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_2\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_3_cascade_\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_5\ : std_logic;
signal \c0.g3_2_1\ : std_logic;
signal \c0.g0_3_0\ : std_logic;
signal \c0.un1_data_in_7__0_0_a2_1_a2_3_cascade_\ : std_logic;
signal \c0.un1_data_in_7__0_0_a2_1_a2_5_0_cascade_\ : std_logic;
signal \c0.tx2_transmit_0_sqmuxa_1\ : std_logic;
signal \c0.un1_data_in_7__3_0_a2_0_a2_3_cascade_\ : std_logic;
signal \c0.N_129\ : std_logic;
signal \c0.data_in_2_Z0Z_1\ : std_logic;
signal \c0.d_4_17\ : std_logic;
signal \c0.data_in_3_Z0Z_6\ : std_logic;
signal \c0.data_in_0_Z0Z_0\ : std_logic;
signal \c0.data_in_2_Z0Z_0\ : std_logic;
signal \c0.d_4_16\ : std_logic;
signal \c0.d_4_0\ : std_logic;
signal \c0.tx2_data_RNO_3Z0Z_0\ : std_logic;
signal \c0.data_in_0_Z0Z_4\ : std_logic;
signal \c0.data_in_4_Z0Z_2\ : std_logic;
signal \c0.data_in_1_Z0Z_3\ : std_logic;
signal \c0.data_in_1_Z0Z_5\ : std_logic;
signal \c0.data_in_2_Z0Z_5\ : std_logic;
signal \c0.data_in_3_Z0Z_1\ : std_logic;
signal \c0.data_in_5_Z0Z_1\ : std_logic;
signal \c0.data_in_3_Z0Z_3\ : std_logic;
signal \c0.tx2_data_1_iv_3_1_6_cascade_\ : std_logic;
signal \c0.d_4_34\ : std_logic;
signal \c0.un1_data_in_7__7_i\ : std_logic;
signal \c0.tx2_data_1_0_i_1_3\ : std_logic;
signal \c0.tx2_data_1_iv_4_1_0_3\ : std_logic;
signal \c0.data_in_1_Z0Z_4\ : std_logic;
signal \c0.data_in_7_Z0Z_3\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_3\ : std_logic;
signal \c0.d_4_14\ : std_logic;
signal \c0.d_4_30\ : std_logic;
signal \c0.tx2_data_1_iv_4_1_6_cascade_\ : std_logic;
signal \c0.data_in_5_Z0Z_3\ : std_logic;
signal \c0.tx2.r_SM_MainZ0Z_2\ : std_logic;
signal \c0.tx2.r_SM_MainZ0Z_0\ : std_logic;
signal \c0.tx2.N_257_cascade_\ : std_logic;
signal \c0.tx2.N_261\ : std_logic;
signal \c0.tx2.o_Tx_Serial12\ : std_logic;
signal \c0.tx2.N_261_cascade_\ : std_logic;
signal \c0.tx2.r_Bit_IndexZ0Z_2\ : std_logic;
signal \c0.tx_transmitZ0\ : std_logic;
signal \c0.tx_active\ : std_logic;
signal \c0.tx2_data_1_iv_4_6\ : std_logic;
signal \c0.tx2_data_1_iv_3_6\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_6\ : std_logic;
signal \c0.d_2_27\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_3\ : std_logic;
signal \c0.data_out_7_Z0Z_7\ : std_logic;
signal \c0.tx_data_RNO_1Z0Z_7\ : std_logic;
signal \c0.tx_data_RNO_3Z0Z_2_cascade_\ : std_logic;
signal \c0.tx_data_1_0_i_ns_1_2\ : std_logic;
signal \c0.d_2_10\ : std_logic;
signal \c0.d_2_42\ : std_logic;
signal \c0.tx_data_RNO_4Z0Z_2\ : std_logic;
signal \c0.N_81\ : std_logic;
signal \c0.d_2_29\ : std_logic;
signal \c0.d_2_30\ : std_logic;
signal \c0.data_out_7_Z0Z_3\ : std_logic;
signal \c0.d_2_31\ : std_logic;
signal \c0.d_2_43\ : std_logic;
signal \c0.d_2_15\ : std_logic;
signal \c0.d_2_2\ : std_logic;
signal \c0.d_2_47\ : std_logic;
signal \c0.un105_newcrc_0_a2_3_cascade_\ : std_logic;
signal \c0.un105_newcrc_0_a2_4\ : std_logic;
signal \c0.d_2_5\ : std_logic;
signal \c0.d_2_32\ : std_logic;
signal \c0.d_2_18\ : std_logic;
signal \c0.d_2_46\ : std_logic;
signal \c0.d_2_20\ : std_logic;
signal \c0.nextCRC16_3_3_1\ : std_logic;
signal \c0.d_2_17\ : std_logic;
signal \c0.d_2_1\ : std_logic;
signal \c0.d_2_4\ : std_logic;
signal \c0.nextCRC16_3_0_a2_1_1\ : std_logic;
signal \c0.un1_data_in_6__4_0_a2_5_a2_1\ : std_logic;
signal \c0.N_133\ : std_logic;
signal \c0.un1_data_in_7__2_0_a2_0_a2_5\ : std_logic;
signal \c0.un1_data_in_6__4\ : std_logic;
signal \c0.wait_for_transmission4_12_5_1_cascade_\ : std_logic;
signal \c0.N_108\ : std_logic;
signal \c0.d_4_32\ : std_logic;
signal \c0.un1_data_in_7__6_0_a2_5_a2_2\ : std_logic;
signal \c0.wait_for_transmission_RNOZ0Z_11\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_4_1\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_4_1_cascade_\ : std_logic;
signal \c0.d_4_47\ : std_logic;
signal \c0.N_125\ : std_logic;
signal \c0.data_in_0_Z0Z_6\ : std_logic;
signal \c0.d_4_6\ : std_logic;
signal \c0.data_in_2_Z0Z_3\ : std_logic;
signal \c0.d_4_19\ : std_logic;
signal \c0.un1_data_in_6__7_0_a2_17_a2_4_1_0\ : std_logic;
signal \c0.data_in_4_Z0Z_3\ : std_logic;
signal \c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_\ : std_logic;
signal \c0.g3_2\ : std_logic;
signal \c0.un1_data_in_6__6_0_a2_0_a2_3_cascade_\ : std_logic;
signal \c0.N_128\ : std_logic;
signal \c0.d_4_41\ : std_logic;
signal \c0.un1_data_in_6__5_0_a2_5_a2_2_cascade_\ : std_logic;
signal \c0.N_132\ : std_logic;
signal \c0.un1_data_in_6__6_0_a2_0_a2_3\ : std_logic;
signal \c0.un1_data_in_6__5_cascade_\ : std_logic;
signal \c0.g0_2_0\ : std_logic;
signal \c0.d_4_43\ : std_logic;
signal \c0.un1_data_in_7__0_0_a2_1_a2_2\ : std_logic;
signal \c0.un1_data_in_6__3_0_a2_5_a2_2_cascade_\ : std_logic;
signal \c0.d_4_25\ : std_logic;
signal \c0.un1_data_in_6__3\ : std_logic;
signal \c0.un1_data_in_6__3_0_a2_5_a2_1\ : std_logic;
signal \c0.data_in_1_Z0Z_1\ : std_logic;
signal \c0.data_in_2_Z0Z_7\ : std_logic;
signal \c0.data_in_5_Z0Z_0\ : std_logic;
signal \c0.d_4_40\ : std_logic;
signal \c0.un1_data_in_7__7_0_a2_0_a2_2\ : std_logic;
signal \c0.data_in_0_Z0Z_5\ : std_logic;
signal \c0.wait_for_transmission_RNOZ0Z_9\ : std_logic;
signal \c0.data_in_2_Z0Z_2\ : std_logic;
signal \c0.data_in_2_Z0Z_4\ : std_logic;
signal \c0.d_4_18\ : std_logic;
signal \c0.N_124\ : std_logic;
signal \c0.N_124_cascade_\ : std_logic;
signal \c0.d_4_RNI21N6Z0Z_11\ : std_logic;
signal \c0.d_4_RNIPF9J2Z0Z_37\ : std_logic;
signal \c0.data_in_4_Z0Z_1\ : std_logic;
signal \c0.d_4_33\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_0\ : std_logic;
signal \c0.data_in_3_Z0Z_2\ : std_logic;
signal \c0.d_4_26\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_1\ : std_logic;
signal \c0.data_in_1_Z0Z_2\ : std_logic;
signal \c0.d_4_10\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_0\ : std_logic;
signal \c0.d_2_36\ : std_logic;
signal \c0.d_2_35\ : std_logic;
signal \c0.N_71\ : std_logic;
signal \c0.tx2.r_Bit_IndexZ0Z_0\ : std_logic;
signal \c0.tx2.r_Clock_Count12_THRU_CO\ : std_logic;
signal \c0.tx2.N_257\ : std_logic;
signal \c0.tx2.N_258_cascade_\ : std_logic;
signal \c0.tx2.r_SM_MainZ0Z_1\ : std_logic;
signal \c0.tx2.r_Bit_IndexZ0Z_1\ : std_logic;
signal \c0.data_out_6_Z0Z_6\ : std_logic;
signal \c0.N_4_0_cascade_\ : std_logic;
signal \c0.N_197\ : std_logic;
signal \c0.data_out_0__1_sqmuxa\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_6\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_3\ : std_logic;
signal \c0.m2_e_1_cascade_\ : std_logic;
signal \c0.N_129_mux_cascade_\ : std_logic;
signal \c0.N_86\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_1\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_4\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_0\ : std_logic;
signal \c0.un144_newcrc_3\ : std_logic;
signal \c0.d_2_34\ : std_logic;
signal \c0.un144_newcrc_4\ : std_logic;
signal \c0.d_2_33\ : std_logic;
signal \c0.data_out_7_Z0Z_6\ : std_logic;
signal \c0.data_out_0__1_sqmuxa_g\ : std_logic;
signal \c0.d_4_12\ : std_logic;
signal \c0.d_4_44\ : std_logic;
signal \c0.tx2_data_1_iv_5_7\ : std_logic;
signal \c0.tx2_data_1_0_i_1_7\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_7\ : std_logic;
signal \c0.d_4_13\ : std_logic;
signal \c0.d_4_29\ : std_logic;
signal \c0.data_in_frame_1__m_5_cascade_\ : std_logic;
signal \c0.tx2_data_1_0_i_1_5\ : std_logic;
signal \c0.tx2_data_1_iv_1_5_cascade_\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_5\ : std_logic;
signal \c0.d_4_15\ : std_logic;
signal \c0.data_in_frame_1__m_7_cascade_\ : std_logic;
signal \c0.d_4_31\ : std_logic;
signal \c0.tx2_data_1_iv_1_7\ : std_logic;
signal \c0.N_205\ : std_logic;
signal \c0.d_4_27\ : std_logic;
signal \c0.N_205_cascade_\ : std_logic;
signal \c0.d_4_11\ : std_logic;
signal \c0.tx2_data_1_iv_4_1_3\ : std_logic;
signal \c0.un1_data_in_6__5\ : std_logic;
signal \c0.i12_THRU_CO\ : std_logic;
signal \c0.N_136\ : std_logic;
signal \c0.wait_for_transmission4_13_1\ : std_logic;
signal \c0.g1_3_cascade_\ : std_logic;
signal \c0.un1_data_in_7__0_0_a2_1_a2_5_0\ : std_logic;
signal \c0.i12_7_c_RNIP740G_cascade_\ : std_logic;
signal \c0.g1_2\ : std_logic;
signal \c0.wait_for_transmission4_12_5\ : std_logic;
signal \c0.un1_data_in_7__3_i\ : std_logic;
signal \c0.g1_5_cascade_\ : std_logic;
signal \c0.wait_for_transmission4_12_4\ : std_logic;
signal \c0.d_4_RNI9LFUVZ0Z_43_cascade_\ : std_logic;
signal \c0.wait_for_transmission_RNI9PP5BZ0Z1_cascade_\ : std_logic;
signal \c0.un1_data_in_6__1_1\ : std_logic;
signal \c0.g0_2_3\ : std_logic;
signal \c0.d_4_23\ : std_logic;
signal \c0.N_126_cascade_\ : std_logic;
signal \c0.un1_data_in_6__1\ : std_logic;
signal \c0.d_4_35\ : std_logic;
signal \c0.data_in_0_Z0Z_7\ : std_logic;
signal \c0.d_4_7\ : std_logic;
signal \c0.data_in_1_Z0Z_0\ : std_logic;
signal \c0.d_4_8\ : std_logic;
signal \c0.d_4_9\ : std_logic;
signal \c0.d_4_39\ : std_logic;
signal \c0.un1_data_in_6__2_0\ : std_logic;
signal \c0.N_107\ : std_logic;
signal \c0.un1_data_in_6__2_0_a2_6_a2_2\ : std_logic;
signal \c0.N_107_cascade_\ : std_logic;
signal \c0.un1_data_in_6__2\ : std_logic;
signal \c0.data_in_2_Z0Z_6\ : std_logic;
signal \c0.d_4_22\ : std_logic;
signal \c0.d_4_RNIU6U8Z0Z_22\ : std_logic;
signal \c0.d_4_RNIU6U8_0Z0Z_22_cascade_\ : std_logic;
signal \c0.d_4_RNIMI4KZ0Z_37\ : std_logic;
signal \c0.data_in_3_Z0Z_0\ : std_logic;
signal \c0.d_4_24\ : std_logic;
signal \c0.N_126\ : std_logic;
signal \c0.un1_data_in_6__1_0_a2_4_a2_1\ : std_logic;
signal \c0.un1_data_in_6__1_0\ : std_logic;
signal \c0.data_in_4_Z0Z_4\ : std_logic;
signal \c0.d_4_36\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_4\ : std_logic;
signal \c0.tx2_data_1_iv_4_1_0_6\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_6\ : std_logic;
signal \c0.d_4_42\ : std_logic;
signal \c0.d_4_46\ : std_logic;
signal \c0.un1_data_in_7__2_0_a2_0_a2_4\ : std_logic;
signal \c0.data_in_4_Z0Z_7\ : std_logic;
signal \c0.rx_data_7\ : std_logic;
signal \c0.data_in_6_Z0Z_1\ : std_logic;
signal \c0.data_in_6_Z0Z_0\ : std_logic;
signal \c0.data_in_7_Z0Z_0\ : std_logic;
signal \c0.data_in_5_Z0Z_4\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_5\ : std_logic;
signal \c0.N_201\ : std_logic;
signal \c0.N_129_mux\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_2\ : std_logic;
signal \GNDG0\ : std_logic;
signal \c0.byte_transmit_counterZ0Z_7\ : std_logic;
signal \c0.byte_transmit_counter15\ : std_logic;
signal \c0.tx2_data_1_iv_5_1_0_4\ : std_logic;
signal \c0.N_207\ : std_logic;
signal \c0.N_207_cascade_\ : std_logic;
signal \c0.d_4_28\ : std_logic;
signal \c0.m2_e_0_2_cascade_\ : std_logic;
signal \c0.N_71_mux\ : std_logic;
signal \c0.d_4_RNII9QU3Z0Z_14\ : std_logic;
signal \c0.wait_for_transmission_RNI94LSZ0Z6\ : std_logic;
signal \c0.wait_for_transmissionZ0\ : std_logic;
signal \c0.d_4_RNI9LFUVZ0Z_43\ : std_logic;
signal \c0.tx2_transmitZ0\ : std_logic;
signal \c0.m2_e_0_2\ : std_logic;
signal \c0.d_4_20\ : std_logic;
signal \c0.N_203_cascade_\ : std_logic;
signal \c0.d_4_4\ : std_logic;
signal \c0.tx2_data_1_iv_5_1_4\ : std_logic;
signal \c0.un1_m4_0_a2_2_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_7\ : std_logic;
signal \c0.un1_m4_0_a2_1_0\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_6\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_5\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_0\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_ac0_3_out_cascade_\ : std_logic;
signal \c0.wait_for_transmission_RNI9PP5BZ0Z1\ : std_logic;
signal \c0.tx2_transmit_0_sqmuxa\ : std_logic;
signal \c0.data_in_4_Z0Z_5\ : std_logic;
signal \c0.data_in_5_Z0Z_5\ : std_logic;
signal \c0.data_in_7_Z0Z_5\ : std_logic;
signal \c0.data_in_6_Z0Z_5\ : std_logic;
signal \c0.data_in_5_Z0Z_6\ : std_logic;
signal \c0.data_in_7_Z0Z_6\ : std_logic;
signal \c0.data_in_6_Z0Z_3\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_3\ : std_logic;
signal \c0.tx2_data_1_0_i_1_6\ : std_logic;
signal \c0.data_in_6_Z0Z_6\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_6\ : std_logic;
signal \c0.data_in_4_Z0Z_6\ : std_logic;
signal \c0.d_4_38\ : std_logic;
signal \c0.d_4_5\ : std_logic;
signal \c0.d_4_21\ : std_logic;
signal \c0.N_203\ : std_logic;
signal \c0.tx2_data_1_iv_5_1_5_cascade_\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_2\ : std_logic;
signal \c0.tx2_data_1_iv_5_5\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_5\ : std_logic;
signal \c0.d_4_37\ : std_logic;
signal \c0.tx2_data_1_iv_5_1_0_5\ : std_logic;
signal \c0.rx.r_Rx_Bytece_1_6\ : std_logic;
signal \c0.rx_data_6\ : std_logic;
signal \c0.rx.r_Rx_Bytece_1_2\ : std_logic;
signal \c0.rx_data_2\ : std_logic;
signal \c0.rx.r_Rx_Bytece_1_4_cascade_\ : std_logic;
signal \c0.rx_data_4\ : std_logic;
signal \c0.rx.r_Bit_IndexZ0Z_2\ : std_logic;
signal \c0.rx.r_Bit_IndexZ0Z_1\ : std_logic;
signal \c0.rx.r_Bit_IndexZ0Z_0\ : std_logic;
signal \c0.rx.r_Rx_DataZ0\ : std_logic;
signal \c0.rx.r_Rx_Bytece_1_0_cascade_\ : std_logic;
signal \c0.rx.r_Rx_Byte_1_sqmuxa\ : std_logic;
signal \c0.rx_data_0\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_ac0_3_out\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_3\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_4\ : std_logic;
signal \c0.un1_byte_transmit_counter2_1_ac0_7_out_0\ : std_logic;
signal \c0.tx2_data_1_iv_5_4\ : std_logic;
signal \c0.tx2_data_1_0_i_1_4\ : std_logic;
signal \c0.tx2_data_1_0_i_1_0_4\ : std_logic;
signal \c0.byte_transmit_counter2Z0Z_1\ : std_logic;
signal \c0.tx2.r_Tx_DataZ0Z_4\ : std_logic;
signal \c0.tx2.r_Tx_Data_0_sqmuxa\ : std_logic;
signal \c0.data_in_5_Z0Z_7\ : std_logic;
signal \c0.data_in_6_Z0Z_4\ : std_logic;
signal \c0.data_in_7_Z0Z_7\ : std_logic;
signal \c0.data_in_6_Z0Z_7\ : std_logic;
signal \c0.rx_data_ready_g\ : std_logic;
signal \c0.data_in_6_Z0Z_2\ : std_logic;
signal \c0.data_in_frame_6_Z0Z_2\ : std_logic;
signal \c0.data_in_7_Z0Z_1\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_1\ : std_logic;
signal \c0.data_in_7_Z0Z_2\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_2\ : std_logic;
signal \c0.data_in_7_Z0Z_4\ : std_logic;
signal \c0.data_in_frame_7_Z0Z_4\ : std_logic;
signal \CLK_c_g\ : std_logic;
signal \c0.data_in_frame_0__0_sqmuxa_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \PIN_1_wire\ : std_logic;
signal \PIN_2_wire\ : std_logic;
signal \PIN_3_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    PIN_1 <= \PIN_1_wire\;
    \PIN_2_wire\ <= PIN_2;
    PIN_3 <= \PIN_3_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \LED_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22335\,
            DIN => \N__22334\,
            DOUT => \N__22333\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22335\,
            PADOUT => \N__22334\,
            PADIN => \N__22333\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8477\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22326\,
            DIN => \N__22325\,
            DOUT => \N__22324\,
            PACKAGEPIN => \PIN_1_wire\
        );

    \PIN_1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22326\,
            PADOUT => \N__22325\,
            PADIN => \N__22324\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__8336\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22317\,
            DIN => \N__22316\,
            DOUT => \N__22315\,
            PACKAGEPIN => \PIN_2_wire\
        );

    \PIN_2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22317\,
            PADOUT => \N__22316\,
            PADIN => \N__22315\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_2_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22308\,
            DIN => \N__22307\,
            DOUT => \N__22306\,
            PACKAGEPIN => \PIN_3_wire\
        );

    \PIN_3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22308\,
            PADOUT => \N__22307\,
            PADIN => \N__22306\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12668\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22299\,
            DIN => \N__22298\,
            DOUT => \N__22297\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22299\,
            PADOUT => \N__22298\,
            PADIN => \N__22297\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22290\,
            DIN => \N__22289\,
            DOUT => \N__22288\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22290\,
            PADOUT => \N__22289\,
            PADIN => \N__22288\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_ibuf_gb_io_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__5372\ : CascadeMux
    port map (
            O => \N__22271\,
            I => \N__22267\
        );

    \I__5371\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22264\
        );

    \I__5370\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22260\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__22264\,
            I => \N__22257\
        );

    \I__5368\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22254\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__22260\,
            I => \N__22251\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__22257\,
            I => \N__22246\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__22254\,
            I => \N__22246\
        );

    \I__5364\ : Span4Mux_h
    port map (
            O => \N__22251\,
            I => \N__22243\
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__22246\,
            I => \c0.data_in_6_Z0Z_4\
        );

    \I__5362\ : Odrv4
    port map (
            O => \N__22243\,
            I => \c0.data_in_6_Z0Z_4\
        );

    \I__5361\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22235\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__22235\,
            I => \N__22231\
        );

    \I__5359\ : InMux
    port map (
            O => \N__22234\,
            I => \N__22228\
        );

    \I__5358\ : Span4Mux_h
    port map (
            O => \N__22231\,
            I => \N__22224\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__22228\,
            I => \N__22221\
        );

    \I__5356\ : CascadeMux
    port map (
            O => \N__22227\,
            I => \N__22218\
        );

    \I__5355\ : Span4Mux_v
    port map (
            O => \N__22224\,
            I => \N__22213\
        );

    \I__5354\ : Span4Mux_h
    port map (
            O => \N__22221\,
            I => \N__22213\
        );

    \I__5353\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22210\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__22213\,
            I => \c0.data_in_7_Z0Z_7\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__22210\,
            I => \c0.data_in_7_Z0Z_7\
        );

    \I__5350\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__22202\,
            I => \N__22197\
        );

    \I__5348\ : InMux
    port map (
            O => \N__22201\,
            I => \N__22194\
        );

    \I__5347\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22191\
        );

    \I__5346\ : Span4Mux_h
    port map (
            O => \N__22197\,
            I => \N__22187\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__22194\,
            I => \N__22184\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__22191\,
            I => \N__22181\
        );

    \I__5343\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22178\
        );

    \I__5342\ : Span4Mux_v
    port map (
            O => \N__22187\,
            I => \N__22173\
        );

    \I__5341\ : Span4Mux_h
    port map (
            O => \N__22184\,
            I => \N__22173\
        );

    \I__5340\ : Span4Mux_h
    port map (
            O => \N__22181\,
            I => \N__22170\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__22178\,
            I => \c0.data_in_6_Z0Z_7\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__22173\,
            I => \c0.data_in_6_Z0Z_7\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__22170\,
            I => \c0.data_in_6_Z0Z_7\
        );

    \I__5336\ : CEMux
    port map (
            O => \N__22163\,
            I => \N__22121\
        );

    \I__5335\ : CEMux
    port map (
            O => \N__22162\,
            I => \N__22121\
        );

    \I__5334\ : CEMux
    port map (
            O => \N__22161\,
            I => \N__22121\
        );

    \I__5333\ : CEMux
    port map (
            O => \N__22160\,
            I => \N__22121\
        );

    \I__5332\ : CEMux
    port map (
            O => \N__22159\,
            I => \N__22121\
        );

    \I__5331\ : CEMux
    port map (
            O => \N__22158\,
            I => \N__22121\
        );

    \I__5330\ : CEMux
    port map (
            O => \N__22157\,
            I => \N__22121\
        );

    \I__5329\ : CEMux
    port map (
            O => \N__22156\,
            I => \N__22121\
        );

    \I__5328\ : CEMux
    port map (
            O => \N__22155\,
            I => \N__22121\
        );

    \I__5327\ : CEMux
    port map (
            O => \N__22154\,
            I => \N__22121\
        );

    \I__5326\ : CEMux
    port map (
            O => \N__22153\,
            I => \N__22121\
        );

    \I__5325\ : CEMux
    port map (
            O => \N__22152\,
            I => \N__22121\
        );

    \I__5324\ : CEMux
    port map (
            O => \N__22151\,
            I => \N__22121\
        );

    \I__5323\ : CEMux
    port map (
            O => \N__22150\,
            I => \N__22121\
        );

    \I__5322\ : GlobalMux
    port map (
            O => \N__22121\,
            I => \N__22118\
        );

    \I__5321\ : gio2CtrlBuf
    port map (
            O => \N__22118\,
            I => \c0.rx_data_ready_g\
        );

    \I__5320\ : InMux
    port map (
            O => \N__22115\,
            I => \N__22112\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__22112\,
            I => \N__22107\
        );

    \I__5318\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22104\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__22110\,
            I => \N__22101\
        );

    \I__5316\ : Span4Mux_h
    port map (
            O => \N__22107\,
            I => \N__22096\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__22104\,
            I => \N__22096\
        );

    \I__5314\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22093\
        );

    \I__5313\ : Odrv4
    port map (
            O => \N__22096\,
            I => \c0.data_in_6_Z0Z_2\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__22093\,
            I => \c0.data_in_6_Z0Z_2\
        );

    \I__5311\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22085\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__5309\ : Span4Mux_h
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__22079\,
            I => \N__22076\
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__22076\,
            I => \c0.data_in_frame_6_Z0Z_2\
        );

    \I__5306\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__22070\,
            I => \N__22066\
        );

    \I__5304\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22063\
        );

    \I__5303\ : Span4Mux_v
    port map (
            O => \N__22066\,
            I => \N__22060\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__22063\,
            I => \N__22057\
        );

    \I__5301\ : Span4Mux_h
    port map (
            O => \N__22060\,
            I => \N__22053\
        );

    \I__5300\ : Span4Mux_h
    port map (
            O => \N__22057\,
            I => \N__22050\
        );

    \I__5299\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22047\
        );

    \I__5298\ : Odrv4
    port map (
            O => \N__22053\,
            I => \c0.data_in_7_Z0Z_1\
        );

    \I__5297\ : Odrv4
    port map (
            O => \N__22050\,
            I => \c0.data_in_7_Z0Z_1\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__22047\,
            I => \c0.data_in_7_Z0Z_1\
        );

    \I__5295\ : CascadeMux
    port map (
            O => \N__22040\,
            I => \N__22037\
        );

    \I__5294\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22034\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__22034\,
            I => \N__22031\
        );

    \I__5292\ : Span4Mux_h
    port map (
            O => \N__22031\,
            I => \N__22028\
        );

    \I__5291\ : Span4Mux_h
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__5290\ : Odrv4
    port map (
            O => \N__22025\,
            I => \c0.data_in_frame_7_Z0Z_1\
        );

    \I__5289\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22019\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__22014\
        );

    \I__5287\ : InMux
    port map (
            O => \N__22018\,
            I => \N__22011\
        );

    \I__5286\ : InMux
    port map (
            O => \N__22017\,
            I => \N__22008\
        );

    \I__5285\ : Span4Mux_v
    port map (
            O => \N__22014\,
            I => \N__22005\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__22011\,
            I => \N__22002\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__22008\,
            I => \N__21999\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__22005\,
            I => \c0.data_in_7_Z0Z_2\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__22002\,
            I => \c0.data_in_7_Z0Z_2\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__21999\,
            I => \c0.data_in_7_Z0Z_2\
        );

    \I__5279\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21989\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__21989\,
            I => \N__21986\
        );

    \I__5277\ : Span12Mux_h
    port map (
            O => \N__21986\,
            I => \N__21983\
        );

    \I__5276\ : Odrv12
    port map (
            O => \N__21983\,
            I => \c0.data_in_frame_7_Z0Z_2\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__5274\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21972\
        );

    \I__5273\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21969\
        );

    \I__5272\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21966\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__21972\,
            I => \N__21963\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__21969\,
            I => \N__21958\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__21966\,
            I => \N__21958\
        );

    \I__5268\ : Span4Mux_h
    port map (
            O => \N__21963\,
            I => \N__21955\
        );

    \I__5267\ : Span4Mux_v
    port map (
            O => \N__21958\,
            I => \N__21952\
        );

    \I__5266\ : Span4Mux_h
    port map (
            O => \N__21955\,
            I => \N__21949\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__21952\,
            I => \c0.data_in_7_Z0Z_4\
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__21949\,
            I => \c0.data_in_7_Z0Z_4\
        );

    \I__5263\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__5261\ : Span4Mux_h
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__21935\,
            I => \c0.data_in_frame_7_Z0Z_4\
        );

    \I__5259\ : ClkMux
    port map (
            O => \N__21932\,
            I => \N__21605\
        );

    \I__5258\ : ClkMux
    port map (
            O => \N__21931\,
            I => \N__21605\
        );

    \I__5257\ : ClkMux
    port map (
            O => \N__21930\,
            I => \N__21605\
        );

    \I__5256\ : ClkMux
    port map (
            O => \N__21929\,
            I => \N__21605\
        );

    \I__5255\ : ClkMux
    port map (
            O => \N__21928\,
            I => \N__21605\
        );

    \I__5254\ : ClkMux
    port map (
            O => \N__21927\,
            I => \N__21605\
        );

    \I__5253\ : ClkMux
    port map (
            O => \N__21926\,
            I => \N__21605\
        );

    \I__5252\ : ClkMux
    port map (
            O => \N__21925\,
            I => \N__21605\
        );

    \I__5251\ : ClkMux
    port map (
            O => \N__21924\,
            I => \N__21605\
        );

    \I__5250\ : ClkMux
    port map (
            O => \N__21923\,
            I => \N__21605\
        );

    \I__5249\ : ClkMux
    port map (
            O => \N__21922\,
            I => \N__21605\
        );

    \I__5248\ : ClkMux
    port map (
            O => \N__21921\,
            I => \N__21605\
        );

    \I__5247\ : ClkMux
    port map (
            O => \N__21920\,
            I => \N__21605\
        );

    \I__5246\ : ClkMux
    port map (
            O => \N__21919\,
            I => \N__21605\
        );

    \I__5245\ : ClkMux
    port map (
            O => \N__21918\,
            I => \N__21605\
        );

    \I__5244\ : ClkMux
    port map (
            O => \N__21917\,
            I => \N__21605\
        );

    \I__5243\ : ClkMux
    port map (
            O => \N__21916\,
            I => \N__21605\
        );

    \I__5242\ : ClkMux
    port map (
            O => \N__21915\,
            I => \N__21605\
        );

    \I__5241\ : ClkMux
    port map (
            O => \N__21914\,
            I => \N__21605\
        );

    \I__5240\ : ClkMux
    port map (
            O => \N__21913\,
            I => \N__21605\
        );

    \I__5239\ : ClkMux
    port map (
            O => \N__21912\,
            I => \N__21605\
        );

    \I__5238\ : ClkMux
    port map (
            O => \N__21911\,
            I => \N__21605\
        );

    \I__5237\ : ClkMux
    port map (
            O => \N__21910\,
            I => \N__21605\
        );

    \I__5236\ : ClkMux
    port map (
            O => \N__21909\,
            I => \N__21605\
        );

    \I__5235\ : ClkMux
    port map (
            O => \N__21908\,
            I => \N__21605\
        );

    \I__5234\ : ClkMux
    port map (
            O => \N__21907\,
            I => \N__21605\
        );

    \I__5233\ : ClkMux
    port map (
            O => \N__21906\,
            I => \N__21605\
        );

    \I__5232\ : ClkMux
    port map (
            O => \N__21905\,
            I => \N__21605\
        );

    \I__5231\ : ClkMux
    port map (
            O => \N__21904\,
            I => \N__21605\
        );

    \I__5230\ : ClkMux
    port map (
            O => \N__21903\,
            I => \N__21605\
        );

    \I__5229\ : ClkMux
    port map (
            O => \N__21902\,
            I => \N__21605\
        );

    \I__5228\ : ClkMux
    port map (
            O => \N__21901\,
            I => \N__21605\
        );

    \I__5227\ : ClkMux
    port map (
            O => \N__21900\,
            I => \N__21605\
        );

    \I__5226\ : ClkMux
    port map (
            O => \N__21899\,
            I => \N__21605\
        );

    \I__5225\ : ClkMux
    port map (
            O => \N__21898\,
            I => \N__21605\
        );

    \I__5224\ : ClkMux
    port map (
            O => \N__21897\,
            I => \N__21605\
        );

    \I__5223\ : ClkMux
    port map (
            O => \N__21896\,
            I => \N__21605\
        );

    \I__5222\ : ClkMux
    port map (
            O => \N__21895\,
            I => \N__21605\
        );

    \I__5221\ : ClkMux
    port map (
            O => \N__21894\,
            I => \N__21605\
        );

    \I__5220\ : ClkMux
    port map (
            O => \N__21893\,
            I => \N__21605\
        );

    \I__5219\ : ClkMux
    port map (
            O => \N__21892\,
            I => \N__21605\
        );

    \I__5218\ : ClkMux
    port map (
            O => \N__21891\,
            I => \N__21605\
        );

    \I__5217\ : ClkMux
    port map (
            O => \N__21890\,
            I => \N__21605\
        );

    \I__5216\ : ClkMux
    port map (
            O => \N__21889\,
            I => \N__21605\
        );

    \I__5215\ : ClkMux
    port map (
            O => \N__21888\,
            I => \N__21605\
        );

    \I__5214\ : ClkMux
    port map (
            O => \N__21887\,
            I => \N__21605\
        );

    \I__5213\ : ClkMux
    port map (
            O => \N__21886\,
            I => \N__21605\
        );

    \I__5212\ : ClkMux
    port map (
            O => \N__21885\,
            I => \N__21605\
        );

    \I__5211\ : ClkMux
    port map (
            O => \N__21884\,
            I => \N__21605\
        );

    \I__5210\ : ClkMux
    port map (
            O => \N__21883\,
            I => \N__21605\
        );

    \I__5209\ : ClkMux
    port map (
            O => \N__21882\,
            I => \N__21605\
        );

    \I__5208\ : ClkMux
    port map (
            O => \N__21881\,
            I => \N__21605\
        );

    \I__5207\ : ClkMux
    port map (
            O => \N__21880\,
            I => \N__21605\
        );

    \I__5206\ : ClkMux
    port map (
            O => \N__21879\,
            I => \N__21605\
        );

    \I__5205\ : ClkMux
    port map (
            O => \N__21878\,
            I => \N__21605\
        );

    \I__5204\ : ClkMux
    port map (
            O => \N__21877\,
            I => \N__21605\
        );

    \I__5203\ : ClkMux
    port map (
            O => \N__21876\,
            I => \N__21605\
        );

    \I__5202\ : ClkMux
    port map (
            O => \N__21875\,
            I => \N__21605\
        );

    \I__5201\ : ClkMux
    port map (
            O => \N__21874\,
            I => \N__21605\
        );

    \I__5200\ : ClkMux
    port map (
            O => \N__21873\,
            I => \N__21605\
        );

    \I__5199\ : ClkMux
    port map (
            O => \N__21872\,
            I => \N__21605\
        );

    \I__5198\ : ClkMux
    port map (
            O => \N__21871\,
            I => \N__21605\
        );

    \I__5197\ : ClkMux
    port map (
            O => \N__21870\,
            I => \N__21605\
        );

    \I__5196\ : ClkMux
    port map (
            O => \N__21869\,
            I => \N__21605\
        );

    \I__5195\ : ClkMux
    port map (
            O => \N__21868\,
            I => \N__21605\
        );

    \I__5194\ : ClkMux
    port map (
            O => \N__21867\,
            I => \N__21605\
        );

    \I__5193\ : ClkMux
    port map (
            O => \N__21866\,
            I => \N__21605\
        );

    \I__5192\ : ClkMux
    port map (
            O => \N__21865\,
            I => \N__21605\
        );

    \I__5191\ : ClkMux
    port map (
            O => \N__21864\,
            I => \N__21605\
        );

    \I__5190\ : ClkMux
    port map (
            O => \N__21863\,
            I => \N__21605\
        );

    \I__5189\ : ClkMux
    port map (
            O => \N__21862\,
            I => \N__21605\
        );

    \I__5188\ : ClkMux
    port map (
            O => \N__21861\,
            I => \N__21605\
        );

    \I__5187\ : ClkMux
    port map (
            O => \N__21860\,
            I => \N__21605\
        );

    \I__5186\ : ClkMux
    port map (
            O => \N__21859\,
            I => \N__21605\
        );

    \I__5185\ : ClkMux
    port map (
            O => \N__21858\,
            I => \N__21605\
        );

    \I__5184\ : ClkMux
    port map (
            O => \N__21857\,
            I => \N__21605\
        );

    \I__5183\ : ClkMux
    port map (
            O => \N__21856\,
            I => \N__21605\
        );

    \I__5182\ : ClkMux
    port map (
            O => \N__21855\,
            I => \N__21605\
        );

    \I__5181\ : ClkMux
    port map (
            O => \N__21854\,
            I => \N__21605\
        );

    \I__5180\ : ClkMux
    port map (
            O => \N__21853\,
            I => \N__21605\
        );

    \I__5179\ : ClkMux
    port map (
            O => \N__21852\,
            I => \N__21605\
        );

    \I__5178\ : ClkMux
    port map (
            O => \N__21851\,
            I => \N__21605\
        );

    \I__5177\ : ClkMux
    port map (
            O => \N__21850\,
            I => \N__21605\
        );

    \I__5176\ : ClkMux
    port map (
            O => \N__21849\,
            I => \N__21605\
        );

    \I__5175\ : ClkMux
    port map (
            O => \N__21848\,
            I => \N__21605\
        );

    \I__5174\ : ClkMux
    port map (
            O => \N__21847\,
            I => \N__21605\
        );

    \I__5173\ : ClkMux
    port map (
            O => \N__21846\,
            I => \N__21605\
        );

    \I__5172\ : ClkMux
    port map (
            O => \N__21845\,
            I => \N__21605\
        );

    \I__5171\ : ClkMux
    port map (
            O => \N__21844\,
            I => \N__21605\
        );

    \I__5170\ : ClkMux
    port map (
            O => \N__21843\,
            I => \N__21605\
        );

    \I__5169\ : ClkMux
    port map (
            O => \N__21842\,
            I => \N__21605\
        );

    \I__5168\ : ClkMux
    port map (
            O => \N__21841\,
            I => \N__21605\
        );

    \I__5167\ : ClkMux
    port map (
            O => \N__21840\,
            I => \N__21605\
        );

    \I__5166\ : ClkMux
    port map (
            O => \N__21839\,
            I => \N__21605\
        );

    \I__5165\ : ClkMux
    port map (
            O => \N__21838\,
            I => \N__21605\
        );

    \I__5164\ : ClkMux
    port map (
            O => \N__21837\,
            I => \N__21605\
        );

    \I__5163\ : ClkMux
    port map (
            O => \N__21836\,
            I => \N__21605\
        );

    \I__5162\ : ClkMux
    port map (
            O => \N__21835\,
            I => \N__21605\
        );

    \I__5161\ : ClkMux
    port map (
            O => \N__21834\,
            I => \N__21605\
        );

    \I__5160\ : ClkMux
    port map (
            O => \N__21833\,
            I => \N__21605\
        );

    \I__5159\ : ClkMux
    port map (
            O => \N__21832\,
            I => \N__21605\
        );

    \I__5158\ : ClkMux
    port map (
            O => \N__21831\,
            I => \N__21605\
        );

    \I__5157\ : ClkMux
    port map (
            O => \N__21830\,
            I => \N__21605\
        );

    \I__5156\ : ClkMux
    port map (
            O => \N__21829\,
            I => \N__21605\
        );

    \I__5155\ : ClkMux
    port map (
            O => \N__21828\,
            I => \N__21605\
        );

    \I__5154\ : ClkMux
    port map (
            O => \N__21827\,
            I => \N__21605\
        );

    \I__5153\ : ClkMux
    port map (
            O => \N__21826\,
            I => \N__21605\
        );

    \I__5152\ : ClkMux
    port map (
            O => \N__21825\,
            I => \N__21605\
        );

    \I__5151\ : ClkMux
    port map (
            O => \N__21824\,
            I => \N__21605\
        );

    \I__5150\ : GlobalMux
    port map (
            O => \N__21605\,
            I => \N__21602\
        );

    \I__5149\ : gio2CtrlBuf
    port map (
            O => \N__21602\,
            I => \CLK_c_g\
        );

    \I__5148\ : CEMux
    port map (
            O => \N__21599\,
            I => \N__21542\
        );

    \I__5147\ : CEMux
    port map (
            O => \N__21598\,
            I => \N__21542\
        );

    \I__5146\ : CEMux
    port map (
            O => \N__21597\,
            I => \N__21542\
        );

    \I__5145\ : CEMux
    port map (
            O => \N__21596\,
            I => \N__21542\
        );

    \I__5144\ : CEMux
    port map (
            O => \N__21595\,
            I => \N__21542\
        );

    \I__5143\ : CEMux
    port map (
            O => \N__21594\,
            I => \N__21542\
        );

    \I__5142\ : CEMux
    port map (
            O => \N__21593\,
            I => \N__21542\
        );

    \I__5141\ : CEMux
    port map (
            O => \N__21592\,
            I => \N__21542\
        );

    \I__5140\ : CEMux
    port map (
            O => \N__21591\,
            I => \N__21542\
        );

    \I__5139\ : CEMux
    port map (
            O => \N__21590\,
            I => \N__21542\
        );

    \I__5138\ : CEMux
    port map (
            O => \N__21589\,
            I => \N__21542\
        );

    \I__5137\ : CEMux
    port map (
            O => \N__21588\,
            I => \N__21542\
        );

    \I__5136\ : CEMux
    port map (
            O => \N__21587\,
            I => \N__21542\
        );

    \I__5135\ : CEMux
    port map (
            O => \N__21586\,
            I => \N__21542\
        );

    \I__5134\ : CEMux
    port map (
            O => \N__21585\,
            I => \N__21542\
        );

    \I__5133\ : CEMux
    port map (
            O => \N__21584\,
            I => \N__21542\
        );

    \I__5132\ : CEMux
    port map (
            O => \N__21583\,
            I => \N__21542\
        );

    \I__5131\ : CEMux
    port map (
            O => \N__21582\,
            I => \N__21542\
        );

    \I__5130\ : CEMux
    port map (
            O => \N__21581\,
            I => \N__21542\
        );

    \I__5129\ : GlobalMux
    port map (
            O => \N__21542\,
            I => \N__21539\
        );

    \I__5128\ : gio2CtrlBuf
    port map (
            O => \N__21539\,
            I => \c0.data_in_frame_0__0_sqmuxa_g\
        );

    \I__5127\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21533\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__21533\,
            I => \N__21530\
        );

    \I__5125\ : Odrv12
    port map (
            O => \N__21530\,
            I => \c0.rx.r_Rx_Bytece_1_2\
        );

    \I__5124\ : CascadeMux
    port map (
            O => \N__21527\,
            I => \N__21523\
        );

    \I__5123\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21520\
        );

    \I__5122\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21517\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__21520\,
            I => \c0.rx_data_2\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__21517\,
            I => \c0.rx_data_2\
        );

    \I__5119\ : CascadeMux
    port map (
            O => \N__21512\,
            I => \c0.rx.r_Rx_Bytece_1_4_cascade_\
        );

    \I__5118\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21505\
        );

    \I__5117\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21502\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__21505\,
            I => \c0.rx_data_4\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__21502\,
            I => \c0.rx_data_4\
        );

    \I__5114\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21491\
        );

    \I__5113\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21486\
        );

    \I__5112\ : InMux
    port map (
            O => \N__21495\,
            I => \N__21486\
        );

    \I__5111\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21482\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21478\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__21486\,
            I => \N__21475\
        );

    \I__5108\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21472\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__21482\,
            I => \N__21468\
        );

    \I__5106\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21465\
        );

    \I__5105\ : Span4Mux_v
    port map (
            O => \N__21478\,
            I => \N__21462\
        );

    \I__5104\ : Span4Mux_h
    port map (
            O => \N__21475\,
            I => \N__21456\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__21472\,
            I => \N__21456\
        );

    \I__5102\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21453\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__21468\,
            I => \N__21447\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21465\,
            I => \N__21447\
        );

    \I__5099\ : Span4Mux_h
    port map (
            O => \N__21462\,
            I => \N__21444\
        );

    \I__5098\ : InMux
    port map (
            O => \N__21461\,
            I => \N__21441\
        );

    \I__5097\ : Span4Mux_h
    port map (
            O => \N__21456\,
            I => \N__21436\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__21453\,
            I => \N__21436\
        );

    \I__5095\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21433\
        );

    \I__5094\ : Span4Mux_h
    port map (
            O => \N__21447\,
            I => \N__21430\
        );

    \I__5093\ : Span4Mux_h
    port map (
            O => \N__21444\,
            I => \N__21425\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__21441\,
            I => \N__21425\
        );

    \I__5091\ : Span4Mux_h
    port map (
            O => \N__21436\,
            I => \N__21422\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__21433\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__21430\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__21425\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__5087\ : Odrv4
    port map (
            O => \N__21422\,
            I => \c0.rx.r_Bit_IndexZ0Z_2\
        );

    \I__5086\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21407\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__21412\,
            I => \N__21404\
        );

    \I__5084\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21400\
        );

    \I__5083\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21397\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__21407\,
            I => \N__21392\
        );

    \I__5081\ : InMux
    port map (
            O => \N__21404\,
            I => \N__21385\
        );

    \I__5080\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21385\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__21400\,
            I => \N__21382\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__21397\,
            I => \N__21379\
        );

    \I__5077\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21376\
        );

    \I__5076\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21373\
        );

    \I__5075\ : Span4Mux_v
    port map (
            O => \N__21392\,
            I => \N__21370\
        );

    \I__5074\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21367\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__21390\,
            I => \N__21364\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__21385\,
            I => \N__21360\
        );

    \I__5071\ : Span4Mux_h
    port map (
            O => \N__21382\,
            I => \N__21357\
        );

    \I__5070\ : Span4Mux_h
    port map (
            O => \N__21379\,
            I => \N__21354\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__21376\,
            I => \N__21349\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__21373\,
            I => \N__21349\
        );

    \I__5067\ : Span4Mux_h
    port map (
            O => \N__21370\,
            I => \N__21344\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__21367\,
            I => \N__21344\
        );

    \I__5065\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21339\
        );

    \I__5064\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21339\
        );

    \I__5063\ : Odrv12
    port map (
            O => \N__21360\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__21357\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__21354\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__21349\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__21344\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__21339\,
            I => \c0.rx.r_Bit_IndexZ0Z_1\
        );

    \I__5057\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21319\
        );

    \I__5056\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21319\
        );

    \I__5055\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21316\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21319\,
            I => \N__21312\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21309\
        );

    \I__5052\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21305\
        );

    \I__5051\ : Span4Mux_h
    port map (
            O => \N__21312\,
            I => \N__21299\
        );

    \I__5050\ : Span4Mux_v
    port map (
            O => \N__21309\,
            I => \N__21299\
        );

    \I__5049\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21296\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21290\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21287\
        );

    \I__5046\ : Span4Mux_h
    port map (
            O => \N__21299\,
            I => \N__21282\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__21296\,
            I => \N__21282\
        );

    \I__5044\ : InMux
    port map (
            O => \N__21295\,
            I => \N__21279\
        );

    \I__5043\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21274\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21271\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__21290\,
            I => \N__21266\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__21287\,
            I => \N__21266\
        );

    \I__5039\ : Span4Mux_h
    port map (
            O => \N__21282\,
            I => \N__21261\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__21279\,
            I => \N__21261\
        );

    \I__5037\ : InMux
    port map (
            O => \N__21278\,
            I => \N__21256\
        );

    \I__5036\ : InMux
    port map (
            O => \N__21277\,
            I => \N__21256\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__21274\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__21271\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__5033\ : Odrv4
    port map (
            O => \N__21266\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__5032\ : Odrv4
    port map (
            O => \N__21261\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__21256\,
            I => \c0.rx.r_Bit_IndexZ0Z_0\
        );

    \I__5030\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21232\
        );

    \I__5029\ : InMux
    port map (
            O => \N__21244\,
            I => \N__21232\
        );

    \I__5028\ : InMux
    port map (
            O => \N__21243\,
            I => \N__21232\
        );

    \I__5027\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21232\
        );

    \I__5026\ : CascadeMux
    port map (
            O => \N__21241\,
            I => \N__21229\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21224\
        );

    \I__5024\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21219\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21219\
        );

    \I__5022\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21215\
        );

    \I__5021\ : Span4Mux_v
    port map (
            O => \N__21224\,
            I => \N__21210\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__21219\,
            I => \N__21207\
        );

    \I__5019\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21204\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21201\
        );

    \I__5017\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21198\
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__21213\,
            I => \N__21195\
        );

    \I__5015\ : Sp12to4
    port map (
            O => \N__21210\,
            I => \N__21190\
        );

    \I__5014\ : Span4Mux_v
    port map (
            O => \N__21207\,
            I => \N__21187\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__21204\,
            I => \N__21184\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__21201\,
            I => \N__21179\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__21198\,
            I => \N__21179\
        );

    \I__5010\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21174\
        );

    \I__5009\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21174\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__21193\,
            I => \N__21171\
        );

    \I__5007\ : Span12Mux_h
    port map (
            O => \N__21190\,
            I => \N__21164\
        );

    \I__5006\ : Sp12to4
    port map (
            O => \N__21187\,
            I => \N__21164\
        );

    \I__5005\ : Span12Mux_v
    port map (
            O => \N__21184\,
            I => \N__21164\
        );

    \I__5004\ : Span4Mux_h
    port map (
            O => \N__21179\,
            I => \N__21159\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__21174\,
            I => \N__21159\
        );

    \I__5002\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21156\
        );

    \I__5001\ : Odrv12
    port map (
            O => \N__21164\,
            I => \c0.rx.r_Rx_DataZ0\
        );

    \I__5000\ : Odrv4
    port map (
            O => \N__21159\,
            I => \c0.rx.r_Rx_DataZ0\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__21156\,
            I => \c0.rx.r_Rx_DataZ0\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__21149\,
            I => \c0.rx.r_Rx_Bytece_1_0_cascade_\
        );

    \I__4997\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21138\
        );

    \I__4996\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21133\
        );

    \I__4995\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21123\
        );

    \I__4994\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21123\
        );

    \I__4993\ : InMux
    port map (
            O => \N__21142\,
            I => \N__21123\
        );

    \I__4992\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21123\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__21138\,
            I => \N__21119\
        );

    \I__4990\ : InMux
    port map (
            O => \N__21137\,
            I => \N__21114\
        );

    \I__4989\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21114\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__21133\,
            I => \N__21111\
        );

    \I__4987\ : InMux
    port map (
            O => \N__21132\,
            I => \N__21108\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__21123\,
            I => \N__21105\
        );

    \I__4985\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21102\
        );

    \I__4984\ : Span4Mux_h
    port map (
            O => \N__21119\,
            I => \N__21097\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__21114\,
            I => \N__21097\
        );

    \I__4982\ : Span4Mux_h
    port map (
            O => \N__21111\,
            I => \N__21093\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__21108\,
            I => \N__21086\
        );

    \I__4980\ : Span12Mux_h
    port map (
            O => \N__21105\,
            I => \N__21086\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__21102\,
            I => \N__21086\
        );

    \I__4978\ : Span4Mux_h
    port map (
            O => \N__21097\,
            I => \N__21083\
        );

    \I__4977\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21080\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__21093\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa\
        );

    \I__4975\ : Odrv12
    port map (
            O => \N__21086\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa\
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__21083\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__21080\,
            I => \c0.rx.r_Rx_Byte_1_sqmuxa\
        );

    \I__4972\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21067\
        );

    \I__4971\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21064\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__21067\,
            I => \c0.rx_data_0\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__21064\,
            I => \c0.rx_data_0\
        );

    \I__4968\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21055\
        );

    \I__4967\ : InMux
    port map (
            O => \N__21058\,
            I => \N__21052\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__21055\,
            I => \N__21049\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__21052\,
            I => \N__21046\
        );

    \I__4964\ : Odrv12
    port map (
            O => \N__21049\,
            I => \c0.un1_byte_transmit_counter2_1_ac0_3_out\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__21046\,
            I => \c0.un1_byte_transmit_counter2_1_ac0_3_out\
        );

    \I__4962\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21034\
        );

    \I__4961\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21034\
        );

    \I__4960\ : InMux
    port map (
            O => \N__21039\,
            I => \N__21029\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__21034\,
            I => \N__21026\
        );

    \I__4958\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21023\
        );

    \I__4957\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21020\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__21029\,
            I => \c0.byte_transmit_counter2Z0Z_3\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__21026\,
            I => \c0.byte_transmit_counter2Z0Z_3\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__21023\,
            I => \c0.byte_transmit_counter2Z0Z_3\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__21020\,
            I => \c0.byte_transmit_counter2Z0Z_3\
        );

    \I__4952\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21006\
        );

    \I__4951\ : InMux
    port map (
            O => \N__21010\,
            I => \N__21002\
        );

    \I__4950\ : InMux
    port map (
            O => \N__21009\,
            I => \N__20999\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__21006\,
            I => \N__20996\
        );

    \I__4948\ : InMux
    port map (
            O => \N__21005\,
            I => \N__20993\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__21002\,
            I => \c0.byte_transmit_counter2Z0Z_4\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__20999\,
            I => \c0.byte_transmit_counter2Z0Z_4\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__20996\,
            I => \c0.byte_transmit_counter2Z0Z_4\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__20993\,
            I => \c0.byte_transmit_counter2Z0Z_4\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__20984\,
            I => \N__20980\
        );

    \I__4942\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20975\
        );

    \I__4941\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20975\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20972\
        );

    \I__4939\ : Odrv4
    port map (
            O => \N__20972\,
            I => \c0.un1_byte_transmit_counter2_1_ac0_7_out_0\
        );

    \I__4938\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__20966\,
            I => \c0.tx2_data_1_iv_5_4\
        );

    \I__4936\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__20960\,
            I => \c0.tx2_data_1_0_i_1_4\
        );

    \I__4934\ : CascadeMux
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__4933\ : InMux
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__20951\,
            I => \N__20948\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__20948\,
            I => \N__20945\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__20945\,
            I => \c0.tx2_data_1_0_i_1_0_4\
        );

    \I__4929\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20934\
        );

    \I__4928\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20934\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__20940\,
            I => \N__20929\
        );

    \I__4926\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20916\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__20934\,
            I => \N__20913\
        );

    \I__4924\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20908\
        );

    \I__4923\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20908\
        );

    \I__4922\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20903\
        );

    \I__4921\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20903\
        );

    \I__4920\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20896\
        );

    \I__4919\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20896\
        );

    \I__4918\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20891\
        );

    \I__4917\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20891\
        );

    \I__4916\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20884\
        );

    \I__4915\ : InMux
    port map (
            O => \N__20922\,
            I => \N__20884\
        );

    \I__4914\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20884\
        );

    \I__4913\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20879\
        );

    \I__4912\ : InMux
    port map (
            O => \N__20919\,
            I => \N__20879\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20875\
        );

    \I__4910\ : Span4Mux_h
    port map (
            O => \N__20913\,
            I => \N__20868\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__20908\,
            I => \N__20868\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__20903\,
            I => \N__20868\
        );

    \I__4907\ : InMux
    port map (
            O => \N__20902\,
            I => \N__20865\
        );

    \I__4906\ : CascadeMux
    port map (
            O => \N__20901\,
            I => \N__20862\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__20896\,
            I => \N__20853\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__20891\,
            I => \N__20853\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__20884\,
            I => \N__20850\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20847\
        );

    \I__4901\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20840\
        );

    \I__4900\ : Span4Mux_v
    port map (
            O => \N__20875\,
            I => \N__20833\
        );

    \I__4899\ : Span4Mux_v
    port map (
            O => \N__20868\,
            I => \N__20833\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__20865\,
            I => \N__20833\
        );

    \I__4897\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20826\
        );

    \I__4896\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20826\
        );

    \I__4895\ : InMux
    port map (
            O => \N__20860\,
            I => \N__20821\
        );

    \I__4894\ : InMux
    port map (
            O => \N__20859\,
            I => \N__20821\
        );

    \I__4893\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20818\
        );

    \I__4892\ : Span4Mux_v
    port map (
            O => \N__20853\,
            I => \N__20813\
        );

    \I__4891\ : Span4Mux_v
    port map (
            O => \N__20850\,
            I => \N__20813\
        );

    \I__4890\ : Span4Mux_v
    port map (
            O => \N__20847\,
            I => \N__20810\
        );

    \I__4889\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20803\
        );

    \I__4888\ : InMux
    port map (
            O => \N__20845\,
            I => \N__20803\
        );

    \I__4887\ : InMux
    port map (
            O => \N__20844\,
            I => \N__20803\
        );

    \I__4886\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20800\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__20840\,
            I => \N__20795\
        );

    \I__4884\ : Span4Mux_h
    port map (
            O => \N__20833\,
            I => \N__20795\
        );

    \I__4883\ : InMux
    port map (
            O => \N__20832\,
            I => \N__20790\
        );

    \I__4882\ : InMux
    port map (
            O => \N__20831\,
            I => \N__20790\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__20826\,
            I => \N__20787\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__20821\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__20818\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4878\ : Odrv4
    port map (
            O => \N__20813\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4877\ : Odrv4
    port map (
            O => \N__20810\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__20803\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__20800\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__20795\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__20790\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4872\ : Odrv12
    port map (
            O => \N__20787\,
            I => \c0.byte_transmit_counter2Z0Z_1\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__4870\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20762\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__20762\,
            I => \N__20759\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__4867\ : Span4Mux_h
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__4866\ : Odrv4
    port map (
            O => \N__20753\,
            I => \c0.tx2.r_Tx_DataZ0Z_4\
        );

    \I__4865\ : CEMux
    port map (
            O => \N__20750\,
            I => \N__20746\
        );

    \I__4864\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20742\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__20746\,
            I => \N__20738\
        );

    \I__4862\ : CEMux
    port map (
            O => \N__20745\,
            I => \N__20735\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__20742\,
            I => \N__20730\
        );

    \I__4860\ : CEMux
    port map (
            O => \N__20741\,
            I => \N__20727\
        );

    \I__4859\ : Span4Mux_v
    port map (
            O => \N__20738\,
            I => \N__20722\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__20735\,
            I => \N__20722\
        );

    \I__4857\ : CEMux
    port map (
            O => \N__20734\,
            I => \N__20719\
        );

    \I__4856\ : CEMux
    port map (
            O => \N__20733\,
            I => \N__20716\
        );

    \I__4855\ : Span4Mux_v
    port map (
            O => \N__20730\,
            I => \N__20710\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__20727\,
            I => \N__20710\
        );

    \I__4853\ : Span4Mux_h
    port map (
            O => \N__20722\,
            I => \N__20707\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__20719\,
            I => \N__20704\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20701\
        );

    \I__4850\ : CascadeMux
    port map (
            O => \N__20715\,
            I => \N__20698\
        );

    \I__4849\ : Span4Mux_v
    port map (
            O => \N__20710\,
            I => \N__20695\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__20707\,
            I => \N__20690\
        );

    \I__4847\ : Span4Mux_h
    port map (
            O => \N__20704\,
            I => \N__20690\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__20701\,
            I => \N__20687\
        );

    \I__4845\ : InMux
    port map (
            O => \N__20698\,
            I => \N__20684\
        );

    \I__4844\ : Span4Mux_h
    port map (
            O => \N__20695\,
            I => \N__20681\
        );

    \I__4843\ : Sp12to4
    port map (
            O => \N__20690\,
            I => \N__20678\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__20687\,
            I => \N__20675\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__20684\,
            I => \c0.tx2.r_Tx_Data_0_sqmuxa\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__20681\,
            I => \c0.tx2.r_Tx_Data_0_sqmuxa\
        );

    \I__4839\ : Odrv12
    port map (
            O => \N__20678\,
            I => \c0.tx2.r_Tx_Data_0_sqmuxa\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__20675\,
            I => \c0.tx2.r_Tx_Data_0_sqmuxa\
        );

    \I__4837\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20662\
        );

    \I__4836\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20659\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__20662\,
            I => \N__20656\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__20659\,
            I => \N__20653\
        );

    \I__4833\ : Span12Mux_v
    port map (
            O => \N__20656\,
            I => \N__20650\
        );

    \I__4832\ : Span4Mux_h
    port map (
            O => \N__20653\,
            I => \N__20647\
        );

    \I__4831\ : Odrv12
    port map (
            O => \N__20650\,
            I => \c0.data_in_5_Z0Z_7\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__20647\,
            I => \c0.data_in_5_Z0Z_7\
        );

    \I__4829\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20638\
        );

    \I__4828\ : CascadeMux
    port map (
            O => \N__20641\,
            I => \N__20635\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__20638\,
            I => \N__20632\
        );

    \I__4826\ : InMux
    port map (
            O => \N__20635\,
            I => \N__20628\
        );

    \I__4825\ : Span12Mux_h
    port map (
            O => \N__20632\,
            I => \N__20625\
        );

    \I__4824\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20622\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__20628\,
            I => \N__20619\
        );

    \I__4822\ : Odrv12
    port map (
            O => \N__20625\,
            I => \c0.data_in_6_Z0Z_3\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__20622\,
            I => \c0.data_in_6_Z0Z_3\
        );

    \I__4820\ : Odrv12
    port map (
            O => \N__20619\,
            I => \c0.data_in_6_Z0Z_3\
        );

    \I__4819\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20606\
        );

    \I__4817\ : Span4Mux_h
    port map (
            O => \N__20606\,
            I => \N__20603\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__20603\,
            I => \c0.data_in_frame_6_Z0Z_3\
        );

    \I__4815\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20597\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__20597\,
            I => \N__20594\
        );

    \I__4813\ : Span4Mux_h
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__20591\,
            I => \c0.tx2_data_1_0_i_1_6\
        );

    \I__4811\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20585\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__20585\,
            I => \N__20580\
        );

    \I__4809\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20577\
        );

    \I__4808\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20574\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__20580\,
            I => \N__20571\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__20577\,
            I => \c0.data_in_6_Z0Z_6\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__20574\,
            I => \c0.data_in_6_Z0Z_6\
        );

    \I__4804\ : Odrv4
    port map (
            O => \N__20571\,
            I => \c0.data_in_6_Z0Z_6\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__20564\,
            I => \N__20561\
        );

    \I__4802\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__20558\,
            I => \c0.data_in_frame_6_Z0Z_6\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20552\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__4798\ : Span4Mux_v
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__4797\ : Span4Mux_h
    port map (
            O => \N__20546\,
            I => \N__20542\
        );

    \I__4796\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20539\
        );

    \I__4795\ : Odrv4
    port map (
            O => \N__20542\,
            I => \c0.data_in_4_Z0Z_6\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__20539\,
            I => \c0.data_in_4_Z0Z_6\
        );

    \I__4793\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20529\
        );

    \I__4792\ : InMux
    port map (
            O => \N__20533\,
            I => \N__20525\
        );

    \I__4791\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20522\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__20529\,
            I => \N__20519\
        );

    \I__4789\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20516\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__20525\,
            I => \N__20508\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__20522\,
            I => \N__20508\
        );

    \I__4786\ : Span4Mux_h
    port map (
            O => \N__20519\,
            I => \N__20508\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__20516\,
            I => \N__20501\
        );

    \I__4784\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20498\
        );

    \I__4783\ : Span4Mux_v
    port map (
            O => \N__20508\,
            I => \N__20495\
        );

    \I__4782\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20486\
        );

    \I__4781\ : InMux
    port map (
            O => \N__20506\,
            I => \N__20486\
        );

    \I__4780\ : InMux
    port map (
            O => \N__20505\,
            I => \N__20486\
        );

    \I__4779\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20486\
        );

    \I__4778\ : Span4Mux_v
    port map (
            O => \N__20501\,
            I => \N__20483\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__20498\,
            I => \c0.d_4_38\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__20495\,
            I => \c0.d_4_38\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__20486\,
            I => \c0.d_4_38\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__20483\,
            I => \c0.d_4_38\
        );

    \I__4773\ : InMux
    port map (
            O => \N__20474\,
            I => \N__20471\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__20471\,
            I => \N__20465\
        );

    \I__4771\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20462\
        );

    \I__4770\ : InMux
    port map (
            O => \N__20469\,
            I => \N__20457\
        );

    \I__4769\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20457\
        );

    \I__4768\ : Odrv4
    port map (
            O => \N__20465\,
            I => \c0.d_4_5\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__20462\,
            I => \c0.d_4_5\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__20457\,
            I => \c0.d_4_5\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__20450\,
            I => \N__20447\
        );

    \I__4764\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__20444\,
            I => \N__20439\
        );

    \I__4762\ : InMux
    port map (
            O => \N__20443\,
            I => \N__20434\
        );

    \I__4761\ : InMux
    port map (
            O => \N__20442\,
            I => \N__20434\
        );

    \I__4760\ : Span4Mux_v
    port map (
            O => \N__20439\,
            I => \N__20431\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__20434\,
            I => \N__20427\
        );

    \I__4758\ : Span4Mux_h
    port map (
            O => \N__20431\,
            I => \N__20424\
        );

    \I__4757\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20421\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__20427\,
            I => \N__20418\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__20424\,
            I => \c0.d_4_21\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__20421\,
            I => \c0.d_4_21\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__20418\,
            I => \c0.d_4_21\
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__20411\,
            I => \N__20404\
        );

    \I__4751\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20399\
        );

    \I__4750\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20399\
        );

    \I__4749\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20392\
        );

    \I__4748\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20392\
        );

    \I__4747\ : InMux
    port map (
            O => \N__20404\,
            I => \N__20392\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__20399\,
            I => \N__20385\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__20392\,
            I => \N__20382\
        );

    \I__4744\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20375\
        );

    \I__4743\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20375\
        );

    \I__4742\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20375\
        );

    \I__4741\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20372\
        );

    \I__4740\ : Span4Mux_h
    port map (
            O => \N__20385\,
            I => \N__20365\
        );

    \I__4739\ : Span4Mux_h
    port map (
            O => \N__20382\,
            I => \N__20365\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__20375\,
            I => \N__20365\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__20372\,
            I => \c0.N_203\
        );

    \I__4736\ : Odrv4
    port map (
            O => \N__20365\,
            I => \c0.N_203\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__20360\,
            I => \c0.tx2_data_1_iv_5_1_5_cascade_\
        );

    \I__4734\ : InMux
    port map (
            O => \N__20357\,
            I => \N__20349\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20356\,
            I => \N__20349\
        );

    \I__4732\ : InMux
    port map (
            O => \N__20355\,
            I => \N__20346\
        );

    \I__4731\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20335\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__20349\,
            I => \N__20329\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__20346\,
            I => \N__20321\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20312\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20312\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20312\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20312\
        );

    \I__4724\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20309\
        );

    \I__4723\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20306\
        );

    \I__4722\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20301\
        );

    \I__4721\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20301\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__20335\,
            I => \N__20298\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20295\
        );

    \I__4718\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20290\
        );

    \I__4717\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20290\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__20329\,
            I => \N__20286\
        );

    \I__4715\ : InMux
    port map (
            O => \N__20328\,
            I => \N__20283\
        );

    \I__4714\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20280\
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__20326\,
            I => \N__20271\
        );

    \I__4712\ : CascadeMux
    port map (
            O => \N__20325\,
            I => \N__20267\
        );

    \I__4711\ : CascadeMux
    port map (
            O => \N__20324\,
            I => \N__20264\
        );

    \I__4710\ : Span4Mux_v
    port map (
            O => \N__20321\,
            I => \N__20255\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__20312\,
            I => \N__20255\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__20309\,
            I => \N__20255\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__20306\,
            I => \N__20255\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__20301\,
            I => \N__20252\
        );

    \I__4705\ : Span4Mux_v
    port map (
            O => \N__20298\,
            I => \N__20245\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__20295\,
            I => \N__20245\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__20290\,
            I => \N__20245\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20242\
        );

    \I__4701\ : Span4Mux_h
    port map (
            O => \N__20286\,
            I => \N__20237\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__20283\,
            I => \N__20237\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20280\,
            I => \N__20234\
        );

    \I__4698\ : InMux
    port map (
            O => \N__20279\,
            I => \N__20229\
        );

    \I__4697\ : InMux
    port map (
            O => \N__20278\,
            I => \N__20229\
        );

    \I__4696\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20216\
        );

    \I__4695\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20216\
        );

    \I__4694\ : InMux
    port map (
            O => \N__20275\,
            I => \N__20216\
        );

    \I__4693\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20216\
        );

    \I__4692\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20216\
        );

    \I__4691\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20216\
        );

    \I__4690\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20211\
        );

    \I__4689\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20211\
        );

    \I__4688\ : Span4Mux_v
    port map (
            O => \N__20255\,
            I => \N__20204\
        );

    \I__4687\ : Span4Mux_v
    port map (
            O => \N__20252\,
            I => \N__20204\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__20245\,
            I => \N__20204\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__20242\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__20237\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__20234\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__20229\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__20216\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__20211\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__20204\,
            I => \c0.byte_transmit_counter2Z0Z_2\
        );

    \I__4678\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__20180\,
            I => \c0.tx2_data_1_iv_5_5\
        );

    \I__4674\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__20174\,
            I => \N__20171\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__20171\,
            I => \c0.data_in_frame_6_Z0Z_5\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20165\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__20165\,
            I => \N__20162\
        );

    \I__4669\ : Span4Mux_v
    port map (
            O => \N__20162\,
            I => \N__20153\
        );

    \I__4668\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20150\
        );

    \I__4667\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20145\
        );

    \I__4666\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20145\
        );

    \I__4665\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20142\
        );

    \I__4664\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20137\
        );

    \I__4663\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20137\
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__20153\,
            I => \c0.d_4_37\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__20150\,
            I => \c0.d_4_37\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20145\,
            I => \c0.d_4_37\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__20142\,
            I => \c0.d_4_37\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__20137\,
            I => \c0.d_4_37\
        );

    \I__4657\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__20123\,
            I => \c0.tx2_data_1_iv_5_1_0_5\
        );

    \I__4655\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__4653\ : Span4Mux_h
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__20111\,
            I => \c0.rx.r_Rx_Bytece_1_6\
        );

    \I__4651\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20104\
        );

    \I__4650\ : CascadeMux
    port map (
            O => \N__20107\,
            I => \N__20101\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20098\
        );

    \I__4648\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20095\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__20098\,
            I => \c0.rx_data_6\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__20095\,
            I => \c0.rx_data_6\
        );

    \I__4645\ : CascadeMux
    port map (
            O => \N__20090\,
            I => \c0.un1_byte_transmit_counter2_1_ac0_3_out_cascade_\
        );

    \I__4644\ : CascadeMux
    port map (
            O => \N__20087\,
            I => \N__20079\
        );

    \I__4643\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20069\
        );

    \I__4642\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20069\
        );

    \I__4641\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20069\
        );

    \I__4640\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20069\
        );

    \I__4639\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20066\
        );

    \I__4638\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20061\
        );

    \I__4637\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20061\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__20069\,
            I => \c0.wait_for_transmission_RNI9PP5BZ0Z1\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__20066\,
            I => \c0.wait_for_transmission_RNI9PP5BZ0Z1\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__20061\,
            I => \c0.wait_for_transmission_RNI9PP5BZ0Z1\
        );

    \I__4633\ : SRMux
    port map (
            O => \N__20054\,
            I => \N__20050\
        );

    \I__4632\ : SRMux
    port map (
            O => \N__20053\,
            I => \N__20047\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__20050\,
            I => \N__20042\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__20047\,
            I => \N__20039\
        );

    \I__4629\ : SRMux
    port map (
            O => \N__20046\,
            I => \N__20036\
        );

    \I__4628\ : SRMux
    port map (
            O => \N__20045\,
            I => \N__20033\
        );

    \I__4627\ : Span4Mux_h
    port map (
            O => \N__20042\,
            I => \N__20028\
        );

    \I__4626\ : Span4Mux_v
    port map (
            O => \N__20039\,
            I => \N__20028\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__20036\,
            I => \N__20025\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__20033\,
            I => \N__20022\
        );

    \I__4623\ : Sp12to4
    port map (
            O => \N__20028\,
            I => \N__20019\
        );

    \I__4622\ : Span12Mux_v
    port map (
            O => \N__20025\,
            I => \N__20016\
        );

    \I__4621\ : Odrv4
    port map (
            O => \N__20022\,
            I => \c0.tx2_transmit_0_sqmuxa\
        );

    \I__4620\ : Odrv12
    port map (
            O => \N__20019\,
            I => \c0.tx2_transmit_0_sqmuxa\
        );

    \I__4619\ : Odrv12
    port map (
            O => \N__20016\,
            I => \c0.tx2_transmit_0_sqmuxa\
        );

    \I__4618\ : InMux
    port map (
            O => \N__20009\,
            I => \N__20006\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__20006\,
            I => \N__20003\
        );

    \I__4616\ : Span4Mux_v
    port map (
            O => \N__20003\,
            I => \N__19999\
        );

    \I__4615\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19996\
        );

    \I__4614\ : Span4Mux_h
    port map (
            O => \N__19999\,
            I => \N__19993\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__19996\,
            I => \N__19990\
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__19993\,
            I => \c0.data_in_4_Z0Z_5\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__19990\,
            I => \c0.data_in_4_Z0Z_5\
        );

    \I__4610\ : InMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__19982\,
            I => \N__19979\
        );

    \I__4608\ : Span12Mux_h
    port map (
            O => \N__19979\,
            I => \N__19975\
        );

    \I__4607\ : InMux
    port map (
            O => \N__19978\,
            I => \N__19972\
        );

    \I__4606\ : Odrv12
    port map (
            O => \N__19975\,
            I => \c0.data_in_5_Z0Z_5\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__19972\,
            I => \c0.data_in_5_Z0Z_5\
        );

    \I__4604\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__19964\,
            I => \N__19958\
        );

    \I__4602\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19955\
        );

    \I__4601\ : CascadeMux
    port map (
            O => \N__19962\,
            I => \N__19951\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__19961\,
            I => \N__19948\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__19958\,
            I => \N__19945\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__19955\,
            I => \N__19942\
        );

    \I__4597\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19935\
        );

    \I__4596\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19935\
        );

    \I__4595\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19935\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__19945\,
            I => \c0.data_in_7_Z0Z_5\
        );

    \I__4593\ : Odrv12
    port map (
            O => \N__19942\,
            I => \c0.data_in_7_Z0Z_5\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__19935\,
            I => \c0.data_in_7_Z0Z_5\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__19928\,
            I => \N__19924\
        );

    \I__4590\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19921\
        );

    \I__4589\ : InMux
    port map (
            O => \N__19924\,
            I => \N__19918\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__19921\,
            I => \N__19915\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__19918\,
            I => \N__19911\
        );

    \I__4586\ : Span4Mux_v
    port map (
            O => \N__19915\,
            I => \N__19908\
        );

    \I__4585\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19905\
        );

    \I__4584\ : Span4Mux_h
    port map (
            O => \N__19911\,
            I => \N__19902\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__19908\,
            I => \c0.data_in_6_Z0Z_5\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__19905\,
            I => \c0.data_in_6_Z0Z_5\
        );

    \I__4581\ : Odrv4
    port map (
            O => \N__19902\,
            I => \c0.data_in_6_Z0Z_5\
        );

    \I__4580\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__4578\ : Span4Mux_v
    port map (
            O => \N__19889\,
            I => \N__19885\
        );

    \I__4577\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19882\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__19885\,
            I => \c0.data_in_5_Z0Z_6\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__19882\,
            I => \c0.data_in_5_Z0Z_6\
        );

    \I__4574\ : CascadeMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__4573\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__19871\,
            I => \N__19866\
        );

    \I__4571\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19863\
        );

    \I__4570\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19860\
        );

    \I__4569\ : Span4Mux_h
    port map (
            O => \N__19866\,
            I => \N__19857\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__19863\,
            I => \c0.data_in_7_Z0Z_6\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__19860\,
            I => \c0.data_in_7_Z0Z_6\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__19857\,
            I => \c0.data_in_7_Z0Z_6\
        );

    \I__4565\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19846\
        );

    \I__4564\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19843\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__19846\,
            I => \N__19840\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__19843\,
            I => \N__19837\
        );

    \I__4561\ : Span12Mux_v
    port map (
            O => \N__19840\,
            I => \N__19834\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__19837\,
            I => \N__19831\
        );

    \I__4559\ : Odrv12
    port map (
            O => \N__19834\,
            I => \c0.d_4_RNII9QU3Z0Z_14\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__19831\,
            I => \c0.d_4_RNII9QU3Z0Z_14\
        );

    \I__4557\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19822\
        );

    \I__4556\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19819\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__19822\,
            I => \N__19814\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__19819\,
            I => \N__19814\
        );

    \I__4553\ : Odrv12
    port map (
            O => \N__19814\,
            I => \c0.wait_for_transmission_RNI94LSZ0Z6\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__4551\ : InMux
    port map (
            O => \N__19808\,
            I => \N__19804\
        );

    \I__4550\ : InMux
    port map (
            O => \N__19807\,
            I => \N__19800\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__19804\,
            I => \N__19797\
        );

    \I__4548\ : InMux
    port map (
            O => \N__19803\,
            I => \N__19794\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__19800\,
            I => \N__19789\
        );

    \I__4546\ : Sp12to4
    port map (
            O => \N__19797\,
            I => \N__19784\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__19794\,
            I => \N__19784\
        );

    \I__4544\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19781\
        );

    \I__4543\ : InMux
    port map (
            O => \N__19792\,
            I => \N__19778\
        );

    \I__4542\ : Odrv4
    port map (
            O => \N__19789\,
            I => \c0.wait_for_transmissionZ0\
        );

    \I__4541\ : Odrv12
    port map (
            O => \N__19784\,
            I => \c0.wait_for_transmissionZ0\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__19781\,
            I => \c0.wait_for_transmissionZ0\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__19778\,
            I => \c0.wait_for_transmissionZ0\
        );

    \I__4538\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__19766\,
            I => \c0.d_4_RNI9LFUVZ0Z_43\
        );

    \I__4536\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__19760\,
            I => \N__19755\
        );

    \I__4534\ : InMux
    port map (
            O => \N__19759\,
            I => \N__19750\
        );

    \I__4533\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19750\
        );

    \I__4532\ : Span12Mux_h
    port map (
            O => \N__19755\,
            I => \N__19747\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__19750\,
            I => \N__19744\
        );

    \I__4530\ : Odrv12
    port map (
            O => \N__19747\,
            I => \c0.tx2_transmitZ0\
        );

    \I__4529\ : Odrv12
    port map (
            O => \N__19744\,
            I => \c0.tx2_transmitZ0\
        );

    \I__4528\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19735\
        );

    \I__4527\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19732\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__19735\,
            I => \c0.m2_e_0_2\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__19732\,
            I => \c0.m2_e_0_2\
        );

    \I__4524\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19723\
        );

    \I__4523\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19720\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__19723\,
            I => \N__19717\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__19720\,
            I => \N__19714\
        );

    \I__4520\ : Span4Mux_v
    port map (
            O => \N__19717\,
            I => \N__19707\
        );

    \I__4519\ : Span4Mux_v
    port map (
            O => \N__19714\,
            I => \N__19707\
        );

    \I__4518\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19702\
        );

    \I__4517\ : InMux
    port map (
            O => \N__19712\,
            I => \N__19702\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__19707\,
            I => \c0.d_4_20\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__19702\,
            I => \c0.d_4_20\
        );

    \I__4514\ : CascadeMux
    port map (
            O => \N__19697\,
            I => \c0.N_203_cascade_\
        );

    \I__4513\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19691\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__19688\,
            I => \N__19684\
        );

    \I__4510\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19681\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__19684\,
            I => \c0.d_4_4\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19681\,
            I => \c0.d_4_4\
        );

    \I__4507\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19673\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__19673\,
            I => \c0.tx2_data_1_iv_5_1_4\
        );

    \I__4505\ : CascadeMux
    port map (
            O => \N__19670\,
            I => \c0.un1_m4_0_a2_2_cascade_\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19663\
        );

    \I__4503\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19660\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__19663\,
            I => \c0.byte_transmit_counter2Z0Z_7\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19660\,
            I => \c0.byte_transmit_counter2Z0Z_7\
        );

    \I__4500\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__19652\,
            I => \c0.un1_m4_0_a2_1_0\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__19649\,
            I => \N__19644\
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__19648\,
            I => \N__19641\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__19647\,
            I => \N__19638\
        );

    \I__4495\ : InMux
    port map (
            O => \N__19644\,
            I => \N__19634\
        );

    \I__4494\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19631\
        );

    \I__4493\ : InMux
    port map (
            O => \N__19638\,
            I => \N__19625\
        );

    \I__4492\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19625\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N__19622\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__19631\,
            I => \N__19619\
        );

    \I__4489\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19616\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__19625\,
            I => \c0.byte_transmit_counter2Z0Z_6\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__19622\,
            I => \c0.byte_transmit_counter2Z0Z_6\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__19619\,
            I => \c0.byte_transmit_counter2Z0Z_6\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__19616\,
            I => \c0.byte_transmit_counter2Z0Z_6\
        );

    \I__4484\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19601\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19606\,
            I => \N__19596\
        );

    \I__4482\ : InMux
    port map (
            O => \N__19605\,
            I => \N__19591\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19591\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__19601\,
            I => \N__19588\
        );

    \I__4479\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19583\
        );

    \I__4478\ : InMux
    port map (
            O => \N__19599\,
            I => \N__19583\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__19596\,
            I => \c0.byte_transmit_counter2Z0Z_5\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__19591\,
            I => \c0.byte_transmit_counter2Z0Z_5\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__19588\,
            I => \c0.byte_transmit_counter2Z0Z_5\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__19583\,
            I => \c0.byte_transmit_counter2Z0Z_5\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__19574\,
            I => \N__19569\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__19573\,
            I => \N__19565\
        );

    \I__4471\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19560\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19553\
        );

    \I__4469\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19553\
        );

    \I__4468\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19553\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__19564\,
            I => \N__19550\
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__19563\,
            I => \N__19547\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__19560\,
            I => \N__19542\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19542\
        );

    \I__4463\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19536\
        );

    \I__4462\ : InMux
    port map (
            O => \N__19547\,
            I => \N__19533\
        );

    \I__4461\ : Span4Mux_h
    port map (
            O => \N__19542\,
            I => \N__19530\
        );

    \I__4460\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19527\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__19540\,
            I => \N__19524\
        );

    \I__4458\ : CascadeMux
    port map (
            O => \N__19539\,
            I => \N__19520\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__19536\,
            I => \N__19515\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__19533\,
            I => \N__19515\
        );

    \I__4455\ : Span4Mux_h
    port map (
            O => \N__19530\,
            I => \N__19510\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__19527\,
            I => \N__19510\
        );

    \I__4453\ : InMux
    port map (
            O => \N__19524\,
            I => \N__19503\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19503\
        );

    \I__4451\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19503\
        );

    \I__4450\ : Span4Mux_v
    port map (
            O => \N__19515\,
            I => \N__19497\
        );

    \I__4449\ : Span4Mux_v
    port map (
            O => \N__19510\,
            I => \N__19497\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__19503\,
            I => \N__19494\
        );

    \I__4447\ : CascadeMux
    port map (
            O => \N__19502\,
            I => \N__19489\
        );

    \I__4446\ : Span4Mux_h
    port map (
            O => \N__19497\,
            I => \N__19475\
        );

    \I__4445\ : Span4Mux_v
    port map (
            O => \N__19494\,
            I => \N__19475\
        );

    \I__4444\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19466\
        );

    \I__4443\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19466\
        );

    \I__4442\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19466\
        );

    \I__4441\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19466\
        );

    \I__4440\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19459\
        );

    \I__4439\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19459\
        );

    \I__4438\ : InMux
    port map (
            O => \N__19485\,
            I => \N__19459\
        );

    \I__4437\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19454\
        );

    \I__4436\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19454\
        );

    \I__4435\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19449\
        );

    \I__4434\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19449\
        );

    \I__4433\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19446\
        );

    \I__4432\ : Sp12to4
    port map (
            O => \N__19475\,
            I => \N__19441\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__19466\,
            I => \N__19441\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__19459\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__19454\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__19449\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19446\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4426\ : Odrv12
    port map (
            O => \N__19441\,
            I => \c0.byte_transmit_counter2Z0Z_0\
        );

    \I__4425\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__4423\ : Span4Mux_h
    port map (
            O => \N__19424\,
            I => \N__19420\
        );

    \I__4422\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19417\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__19420\,
            I => \c0.N_201\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__19417\,
            I => \c0.N_201\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19407\
        );

    \I__4418\ : InMux
    port map (
            O => \N__19411\,
            I => \N__19404\
        );

    \I__4417\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19393\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__19407\,
            I => \N__19388\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__19404\,
            I => \N__19388\
        );

    \I__4414\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19381\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19381\
        );

    \I__4412\ : InMux
    port map (
            O => \N__19401\,
            I => \N__19381\
        );

    \I__4411\ : InMux
    port map (
            O => \N__19400\,
            I => \N__19376\
        );

    \I__4410\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19376\
        );

    \I__4409\ : InMux
    port map (
            O => \N__19398\,
            I => \N__19367\
        );

    \I__4408\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19364\
        );

    \I__4407\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19358\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__19393\,
            I => \N__19351\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__19388\,
            I => \N__19351\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__19381\,
            I => \N__19351\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19376\,
            I => \N__19348\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19375\,
            I => \N__19337\
        );

    \I__4401\ : InMux
    port map (
            O => \N__19374\,
            I => \N__19337\
        );

    \I__4400\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19337\
        );

    \I__4399\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19337\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19337\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19334\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__19367\,
            I => \N__19331\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__19364\,
            I => \N__19328\
        );

    \I__4394\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19323\
        );

    \I__4393\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19323\
        );

    \I__4392\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19315\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__19358\,
            I => \N__19302\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__19351\,
            I => \N__19302\
        );

    \I__4389\ : Span4Mux_v
    port map (
            O => \N__19348\,
            I => \N__19302\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__19337\,
            I => \N__19302\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__19334\,
            I => \N__19293\
        );

    \I__4386\ : Span4Mux_v
    port map (
            O => \N__19331\,
            I => \N__19293\
        );

    \I__4385\ : Span4Mux_v
    port map (
            O => \N__19328\,
            I => \N__19293\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__19323\,
            I => \N__19293\
        );

    \I__4383\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19288\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19321\,
            I => \N__19288\
        );

    \I__4381\ : InMux
    port map (
            O => \N__19320\,
            I => \N__19283\
        );

    \I__4380\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19278\
        );

    \I__4379\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19278\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__19315\,
            I => \N__19275\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19266\
        );

    \I__4376\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19266\
        );

    \I__4375\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19266\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19266\
        );

    \I__4373\ : Span4Mux_h
    port map (
            O => \N__19302\,
            I => \N__19263\
        );

    \I__4372\ : Span4Mux_h
    port map (
            O => \N__19293\,
            I => \N__19258\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__19288\,
            I => \N__19258\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19253\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19253\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__19283\,
            I => \c0.N_129_mux\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__19278\,
            I => \c0.N_129_mux\
        );

    \I__4366\ : Odrv12
    port map (
            O => \N__19275\,
            I => \c0.N_129_mux\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__19266\,
            I => \c0.N_129_mux\
        );

    \I__4364\ : Odrv4
    port map (
            O => \N__19263\,
            I => \c0.N_129_mux\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__19258\,
            I => \c0.N_129_mux\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__19253\,
            I => \c0.N_129_mux\
        );

    \I__4361\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19229\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__19237\,
            I => \N__19226\
        );

    \I__4359\ : CascadeMux
    port map (
            O => \N__19236\,
            I => \N__19223\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__19235\,
            I => \N__19219\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__19234\,
            I => \N__19215\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__19233\,
            I => \N__19210\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__19232\,
            I => \N__19206\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__19229\,
            I => \N__19197\
        );

    \I__4353\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19186\
        );

    \I__4352\ : InMux
    port map (
            O => \N__19223\,
            I => \N__19186\
        );

    \I__4351\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19186\
        );

    \I__4350\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19186\
        );

    \I__4349\ : InMux
    port map (
            O => \N__19218\,
            I => \N__19186\
        );

    \I__4348\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19182\
        );

    \I__4347\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19179\
        );

    \I__4346\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19174\
        );

    \I__4345\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19174\
        );

    \I__4344\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19163\
        );

    \I__4343\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19163\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19159\
        );

    \I__4341\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19153\
        );

    \I__4340\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19153\
        );

    \I__4339\ : InMux
    port map (
            O => \N__19202\,
            I => \N__19146\
        );

    \I__4338\ : InMux
    port map (
            O => \N__19201\,
            I => \N__19146\
        );

    \I__4337\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19146\
        );

    \I__4336\ : Span4Mux_h
    port map (
            O => \N__19197\,
            I => \N__19143\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__19186\,
            I => \N__19140\
        );

    \I__4334\ : InMux
    port map (
            O => \N__19185\,
            I => \N__19137\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__19182\,
            I => \N__19134\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__19179\,
            I => \N__19129\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__19174\,
            I => \N__19129\
        );

    \I__4330\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19120\
        );

    \I__4329\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19120\
        );

    \I__4328\ : InMux
    port map (
            O => \N__19171\,
            I => \N__19120\
        );

    \I__4327\ : InMux
    port map (
            O => \N__19170\,
            I => \N__19120\
        );

    \I__4326\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19115\
        );

    \I__4325\ : InMux
    port map (
            O => \N__19168\,
            I => \N__19115\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__19163\,
            I => \N__19110\
        );

    \I__4323\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19107\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__19159\,
            I => \N__19104\
        );

    \I__4321\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19101\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__19153\,
            I => \N__19096\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19146\,
            I => \N__19096\
        );

    \I__4318\ : Span4Mux_h
    port map (
            O => \N__19143\,
            I => \N__19081\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__19140\,
            I => \N__19081\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__19137\,
            I => \N__19081\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__19134\,
            I => \N__19081\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__19129\,
            I => \N__19081\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__19120\,
            I => \N__19081\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__19115\,
            I => \N__19081\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__19114\,
            I => \N__19078\
        );

    \I__4310\ : InMux
    port map (
            O => \N__19113\,
            I => \N__19073\
        );

    \I__4309\ : Span12Mux_h
    port map (
            O => \N__19110\,
            I => \N__19070\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__19107\,
            I => \N__19061\
        );

    \I__4307\ : Span12Mux_s8_h
    port map (
            O => \N__19104\,
            I => \N__19061\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__19101\,
            I => \N__19061\
        );

    \I__4305\ : Span12Mux_s9_v
    port map (
            O => \N__19096\,
            I => \N__19061\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__19081\,
            I => \N__19058\
        );

    \I__4303\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19051\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19077\,
            I => \N__19051\
        );

    \I__4301\ : InMux
    port map (
            O => \N__19076\,
            I => \N__19051\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__19073\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__4299\ : Odrv12
    port map (
            O => \N__19070\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__4298\ : Odrv12
    port map (
            O => \N__19061\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__4297\ : Odrv4
    port map (
            O => \N__19058\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__19051\,
            I => \c0.byte_transmit_counterZ0Z_2\
        );

    \I__4295\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__19037\,
            I => \c0.byte_transmit_counterZ0Z_7\
        );

    \I__4293\ : CEMux
    port map (
            O => \N__19034\,
            I => \N__19031\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__19031\,
            I => \N__19026\
        );

    \I__4291\ : CEMux
    port map (
            O => \N__19030\,
            I => \N__19023\
        );

    \I__4290\ : CEMux
    port map (
            O => \N__19029\,
            I => \N__19020\
        );

    \I__4289\ : Span4Mux_h
    port map (
            O => \N__19026\,
            I => \N__19016\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__19023\,
            I => \N__19013\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__19020\,
            I => \N__19010\
        );

    \I__4286\ : InMux
    port map (
            O => \N__19019\,
            I => \N__19007\
        );

    \I__4285\ : Odrv4
    port map (
            O => \N__19016\,
            I => \c0.byte_transmit_counter15\
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__19013\,
            I => \c0.byte_transmit_counter15\
        );

    \I__4283\ : Odrv12
    port map (
            O => \N__19010\,
            I => \c0.byte_transmit_counter15\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__19007\,
            I => \c0.byte_transmit_counter15\
        );

    \I__4281\ : CascadeMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__4280\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__18992\,
            I => \N__18989\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__18989\,
            I => \c0.tx2_data_1_iv_5_1_0_4\
        );

    \I__4277\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18982\
        );

    \I__4276\ : InMux
    port map (
            O => \N__18985\,
            I => \N__18979\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__18982\,
            I => \N__18976\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__18979\,
            I => \c0.N_207\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__18976\,
            I => \c0.N_207\
        );

    \I__4272\ : CascadeMux
    port map (
            O => \N__18971\,
            I => \c0.N_207_cascade_\
        );

    \I__4271\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18964\
        );

    \I__4270\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18961\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__18964\,
            I => \N__18958\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18953\
        );

    \I__4267\ : Span12Mux_h
    port map (
            O => \N__18958\,
            I => \N__18950\
        );

    \I__4266\ : InMux
    port map (
            O => \N__18957\,
            I => \N__18947\
        );

    \I__4265\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18944\
        );

    \I__4264\ : Span4Mux_h
    port map (
            O => \N__18953\,
            I => \N__18941\
        );

    \I__4263\ : Odrv12
    port map (
            O => \N__18950\,
            I => \c0.d_4_28\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__18947\,
            I => \c0.d_4_28\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__18944\,
            I => \c0.d_4_28\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__18941\,
            I => \c0.d_4_28\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__18932\,
            I => \c0.m2_e_0_2_cascade_\
        );

    \I__4258\ : InMux
    port map (
            O => \N__18929\,
            I => \N__18912\
        );

    \I__4257\ : InMux
    port map (
            O => \N__18928\,
            I => \N__18912\
        );

    \I__4256\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18912\
        );

    \I__4255\ : InMux
    port map (
            O => \N__18926\,
            I => \N__18912\
        );

    \I__4254\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18907\
        );

    \I__4253\ : InMux
    port map (
            O => \N__18924\,
            I => \N__18898\
        );

    \I__4252\ : InMux
    port map (
            O => \N__18923\,
            I => \N__18898\
        );

    \I__4251\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18898\
        );

    \I__4250\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18898\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__18912\,
            I => \N__18892\
        );

    \I__4248\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18889\
        );

    \I__4247\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18886\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__18907\,
            I => \N__18881\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__18898\,
            I => \N__18881\
        );

    \I__4244\ : InMux
    port map (
            O => \N__18897\,
            I => \N__18874\
        );

    \I__4243\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18874\
        );

    \I__4242\ : InMux
    port map (
            O => \N__18895\,
            I => \N__18874\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__18892\,
            I => \N__18868\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__18889\,
            I => \N__18868\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__18886\,
            I => \N__18861\
        );

    \I__4238\ : Span4Mux_v
    port map (
            O => \N__18881\,
            I => \N__18861\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__18874\,
            I => \N__18861\
        );

    \I__4236\ : InMux
    port map (
            O => \N__18873\,
            I => \N__18858\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__18868\,
            I => \N__18853\
        );

    \I__4234\ : Span4Mux_h
    port map (
            O => \N__18861\,
            I => \N__18853\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__18858\,
            I => \c0.N_71_mux\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__18853\,
            I => \c0.N_71_mux\
        );

    \I__4231\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18845\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__18842\,
            I => \N__18838\
        );

    \I__4228\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18835\
        );

    \I__4227\ : Span4Mux_h
    port map (
            O => \N__18838\,
            I => \N__18830\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__18835\,
            I => \N__18830\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__18830\,
            I => \c0.data_in_4_Z0Z_7\
        );

    \I__4224\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18823\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__18826\,
            I => \N__18820\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__18823\,
            I => \N__18817\
        );

    \I__4221\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18814\
        );

    \I__4220\ : Odrv12
    port map (
            O => \N__18817\,
            I => \c0.rx_data_7\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__18814\,
            I => \c0.rx_data_7\
        );

    \I__4218\ : InMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__18806\,
            I => \N__18802\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18798\
        );

    \I__4215\ : Span4Mux_h
    port map (
            O => \N__18802\,
            I => \N__18795\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18792\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__18798\,
            I => \N__18789\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__18795\,
            I => \c0.data_in_6_Z0Z_1\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__18792\,
            I => \c0.data_in_6_Z0Z_1\
        );

    \I__4210\ : Odrv4
    port map (
            O => \N__18789\,
            I => \c0.data_in_6_Z0Z_1\
        );

    \I__4209\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18778\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__18781\,
            I => \N__18775\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__18778\,
            I => \N__18772\
        );

    \I__4206\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18769\
        );

    \I__4205\ : Span4Mux_h
    port map (
            O => \N__18772\,
            I => \N__18766\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__18769\,
            I => \N__18762\
        );

    \I__4203\ : Span4Mux_h
    port map (
            O => \N__18766\,
            I => \N__18759\
        );

    \I__4202\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18756\
        );

    \I__4201\ : Span4Mux_h
    port map (
            O => \N__18762\,
            I => \N__18753\
        );

    \I__4200\ : Odrv4
    port map (
            O => \N__18759\,
            I => \c0.data_in_6_Z0Z_0\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__18756\,
            I => \c0.data_in_6_Z0Z_0\
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__18753\,
            I => \c0.data_in_6_Z0Z_0\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__4196\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18739\
        );

    \I__4195\ : InMux
    port map (
            O => \N__18742\,
            I => \N__18735\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__18739\,
            I => \N__18732\
        );

    \I__4193\ : InMux
    port map (
            O => \N__18738\,
            I => \N__18729\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__18735\,
            I => \N__18724\
        );

    \I__4191\ : Span4Mux_v
    port map (
            O => \N__18732\,
            I => \N__18724\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__18729\,
            I => \c0.data_in_7_Z0Z_0\
        );

    \I__4189\ : Odrv4
    port map (
            O => \N__18724\,
            I => \c0.data_in_7_Z0Z_0\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18715\
        );

    \I__4187\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18712\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__18715\,
            I => \N__18709\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__18712\,
            I => \N__18706\
        );

    \I__4184\ : Span12Mux_h
    port map (
            O => \N__18709\,
            I => \N__18703\
        );

    \I__4183\ : Span4Mux_h
    port map (
            O => \N__18706\,
            I => \N__18700\
        );

    \I__4182\ : Odrv12
    port map (
            O => \N__18703\,
            I => \c0.data_in_5_Z0Z_4\
        );

    \I__4181\ : Odrv4
    port map (
            O => \N__18700\,
            I => \c0.data_in_5_Z0Z_4\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__18692\,
            I => \c0.byte_transmit_counterZ0Z_5\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18689\,
            I => \N__18686\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__18686\,
            I => \c0.d_4_RNIU6U8Z0Z_22\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__18683\,
            I => \c0.d_4_RNIU6U8_0Z0Z_22_cascade_\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18677\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__18677\,
            I => \c0.d_4_RNIMI4KZ0Z_37\
        );

    \I__4173\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18670\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18667\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__18670\,
            I => \N__18663\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__18667\,
            I => \N__18660\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18657\
        );

    \I__4168\ : Odrv4
    port map (
            O => \N__18663\,
            I => \c0.data_in_3_Z0Z_0\
        );

    \I__4167\ : Odrv12
    port map (
            O => \N__18660\,
            I => \c0.data_in_3_Z0Z_0\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__18657\,
            I => \c0.data_in_3_Z0Z_0\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__18650\,
            I => \N__18645\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18641\
        );

    \I__4163\ : InMux
    port map (
            O => \N__18648\,
            I => \N__18637\
        );

    \I__4162\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18634\
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__18644\,
            I => \N__18631\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__18641\,
            I => \N__18628\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__18640\,
            I => \N__18623\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__18637\,
            I => \N__18620\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__18634\,
            I => \N__18617\
        );

    \I__4156\ : InMux
    port map (
            O => \N__18631\,
            I => \N__18614\
        );

    \I__4155\ : Span4Mux_h
    port map (
            O => \N__18628\,
            I => \N__18611\
        );

    \I__4154\ : InMux
    port map (
            O => \N__18627\,
            I => \N__18604\
        );

    \I__4153\ : InMux
    port map (
            O => \N__18626\,
            I => \N__18604\
        );

    \I__4152\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18604\
        );

    \I__4151\ : Span4Mux_h
    port map (
            O => \N__18620\,
            I => \N__18599\
        );

    \I__4150\ : Span4Mux_h
    port map (
            O => \N__18617\,
            I => \N__18599\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__18614\,
            I => \c0.d_4_24\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__18611\,
            I => \c0.d_4_24\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__18604\,
            I => \c0.d_4_24\
        );

    \I__4146\ : Odrv4
    port map (
            O => \N__18599\,
            I => \c0.d_4_24\
        );

    \I__4145\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18586\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__18589\,
            I => \N__18583\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__18586\,
            I => \N__18579\
        );

    \I__4142\ : InMux
    port map (
            O => \N__18583\,
            I => \N__18576\
        );

    \I__4141\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18573\
        );

    \I__4140\ : Span4Mux_v
    port map (
            O => \N__18579\,
            I => \N__18569\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__18576\,
            I => \N__18564\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18564\
        );

    \I__4137\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18561\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__18569\,
            I => \c0.N_126\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__18564\,
            I => \c0.N_126\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__18561\,
            I => \c0.N_126\
        );

    \I__4133\ : InMux
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__18551\,
            I => \N__18546\
        );

    \I__4131\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18541\
        );

    \I__4130\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18541\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__18546\,
            I => \c0.un1_data_in_6__1_0_a2_4_a2_1\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__18541\,
            I => \c0.un1_data_in_6__1_0_a2_4_a2_1\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__4124\ : Span12Mux_v
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__4123\ : Odrv12
    port map (
            O => \N__18524\,
            I => \c0.un1_data_in_6__1_0\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__4120\ : Span4Mux_v
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__4119\ : Span4Mux_h
    port map (
            O => \N__18512\,
            I => \N__18508\
        );

    \I__4118\ : InMux
    port map (
            O => \N__18511\,
            I => \N__18505\
        );

    \I__4117\ : Odrv4
    port map (
            O => \N__18508\,
            I => \c0.data_in_4_Z0Z_4\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__18505\,
            I => \c0.data_in_4_Z0Z_4\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__4114\ : InMux
    port map (
            O => \N__18497\,
            I => \N__18487\
        );

    \I__4113\ : InMux
    port map (
            O => \N__18496\,
            I => \N__18487\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__18495\,
            I => \N__18483\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18494\,
            I => \N__18477\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18493\,
            I => \N__18477\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18492\,
            I => \N__18474\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__18487\,
            I => \N__18471\
        );

    \I__4107\ : InMux
    port map (
            O => \N__18486\,
            I => \N__18464\
        );

    \I__4106\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18464\
        );

    \I__4105\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18464\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__18477\,
            I => \c0.d_4_36\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__18474\,
            I => \c0.d_4_36\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__18471\,
            I => \c0.d_4_36\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__18464\,
            I => \c0.d_4_36\
        );

    \I__4100\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18452\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__18452\,
            I => \c0.data_in_frame_6_Z0Z_4\
        );

    \I__4098\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__18440\,
            I => \c0.tx2_data_1_iv_4_1_0_6\
        );

    \I__4094\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__18434\,
            I => \c0.data_in_frame_7_Z0Z_6\
        );

    \I__4092\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18424\
        );

    \I__4091\ : InMux
    port map (
            O => \N__18430\,
            I => \N__18424\
        );

    \I__4090\ : InMux
    port map (
            O => \N__18429\,
            I => \N__18420\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18424\,
            I => \N__18416\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__18423\,
            I => \N__18413\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18420\,
            I => \N__18408\
        );

    \I__4086\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18405\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__18416\,
            I => \N__18402\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18397\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18412\,
            I => \N__18397\
        );

    \I__4082\ : InMux
    port map (
            O => \N__18411\,
            I => \N__18394\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__18408\,
            I => \N__18391\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__18405\,
            I => \N__18388\
        );

    \I__4079\ : Span4Mux_h
    port map (
            O => \N__18402\,
            I => \N__18385\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__18397\,
            I => \N__18382\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__18394\,
            I => \c0.d_4_42\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__18391\,
            I => \c0.d_4_42\
        );

    \I__4075\ : Odrv12
    port map (
            O => \N__18388\,
            I => \c0.d_4_42\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__18385\,
            I => \c0.d_4_42\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__18382\,
            I => \c0.d_4_42\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__18371\,
            I => \N__18365\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__18370\,
            I => \N__18362\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18357\
        );

    \I__4069\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18357\
        );

    \I__4068\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18352\
        );

    \I__4067\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18352\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__18357\,
            I => \c0.d_4_46\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__18352\,
            I => \c0.d_4_46\
        );

    \I__4064\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__4062\ : Span4Mux_v
    port map (
            O => \N__18341\,
            I => \N__18338\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__18338\,
            I => \c0.un1_data_in_7__2_0_a2_0_a2_4\
        );

    \I__4060\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18331\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18328\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__18331\,
            I => \N__18323\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__18328\,
            I => \N__18323\
        );

    \I__4056\ : Span4Mux_v
    port map (
            O => \N__18323\,
            I => \N__18318\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18322\,
            I => \N__18313\
        );

    \I__4054\ : InMux
    port map (
            O => \N__18321\,
            I => \N__18313\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__18318\,
            I => \c0.d_4_7\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__18313\,
            I => \c0.d_4_7\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__4049\ : Span4Mux_v
    port map (
            O => \N__18302\,
            I => \N__18298\
        );

    \I__4048\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18294\
        );

    \I__4047\ : Span4Mux_h
    port map (
            O => \N__18298\,
            I => \N__18291\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18297\,
            I => \N__18288\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__18294\,
            I => \c0.data_in_1_Z0Z_0\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__18291\,
            I => \c0.data_in_1_Z0Z_0\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__18288\,
            I => \c0.data_in_1_Z0Z_0\
        );

    \I__4042\ : InMux
    port map (
            O => \N__18281\,
            I => \N__18277\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__18280\,
            I => \N__18274\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__18277\,
            I => \N__18269\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18262\
        );

    \I__4038\ : InMux
    port map (
            O => \N__18273\,
            I => \N__18262\
        );

    \I__4037\ : InMux
    port map (
            O => \N__18272\,
            I => \N__18262\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__18269\,
            I => \c0.d_4_8\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__18262\,
            I => \c0.d_4_8\
        );

    \I__4034\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__18254\,
            I => \N__18249\
        );

    \I__4032\ : InMux
    port map (
            O => \N__18253\,
            I => \N__18245\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18252\,
            I => \N__18242\
        );

    \I__4030\ : Span4Mux_v
    port map (
            O => \N__18249\,
            I => \N__18238\
        );

    \I__4029\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18235\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__18245\,
            I => \N__18230\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__18242\,
            I => \N__18230\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18241\,
            I => \N__18227\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__18238\,
            I => \c0.d_4_9\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__18235\,
            I => \c0.d_4_9\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__18230\,
            I => \c0.d_4_9\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__18227\,
            I => \c0.d_4_9\
        );

    \I__4021\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18215\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__18215\,
            I => \N__18212\
        );

    \I__4019\ : Span4Mux_v
    port map (
            O => \N__18212\,
            I => \N__18206\
        );

    \I__4018\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18203\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18210\,
            I => \N__18200\
        );

    \I__4016\ : InMux
    port map (
            O => \N__18209\,
            I => \N__18197\
        );

    \I__4015\ : Odrv4
    port map (
            O => \N__18206\,
            I => \c0.d_4_39\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__18203\,
            I => \c0.d_4_39\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__18200\,
            I => \c0.d_4_39\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__18197\,
            I => \c0.d_4_39\
        );

    \I__4011\ : InMux
    port map (
            O => \N__18188\,
            I => \N__18185\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__18185\,
            I => \c0.un1_data_in_6__2_0\
        );

    \I__4009\ : InMux
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__18179\,
            I => \N__18174\
        );

    \I__4007\ : InMux
    port map (
            O => \N__18178\,
            I => \N__18171\
        );

    \I__4006\ : InMux
    port map (
            O => \N__18177\,
            I => \N__18168\
        );

    \I__4005\ : Span4Mux_h
    port map (
            O => \N__18174\,
            I => \N__18165\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__18171\,
            I => \N__18162\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__18168\,
            I => \c0.N_107\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__18165\,
            I => \c0.N_107\
        );

    \I__4001\ : Odrv4
    port map (
            O => \N__18162\,
            I => \c0.N_107\
        );

    \I__4000\ : InMux
    port map (
            O => \N__18155\,
            I => \N__18149\
        );

    \I__3999\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18149\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__18149\,
            I => \c0.un1_data_in_6__2_0_a2_6_a2_2\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__18146\,
            I => \c0.N_107_cascade_\
        );

    \I__3996\ : InMux
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__18140\,
            I => \N__18136\
        );

    \I__3994\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18133\
        );

    \I__3993\ : Span4Mux_h
    port map (
            O => \N__18136\,
            I => \N__18130\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__18133\,
            I => \N__18127\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__18130\,
            I => \c0.un1_data_in_6__2\
        );

    \I__3990\ : Odrv4
    port map (
            O => \N__18127\,
            I => \c0.un1_data_in_6__2\
        );

    \I__3989\ : InMux
    port map (
            O => \N__18122\,
            I => \N__18118\
        );

    \I__3988\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18115\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__18118\,
            I => \N__18111\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__18115\,
            I => \N__18108\
        );

    \I__3985\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18105\
        );

    \I__3984\ : Span4Mux_h
    port map (
            O => \N__18111\,
            I => \N__18102\
        );

    \I__3983\ : Span4Mux_h
    port map (
            O => \N__18108\,
            I => \N__18099\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__18105\,
            I => \c0.data_in_2_Z0Z_6\
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__18102\,
            I => \c0.data_in_2_Z0Z_6\
        );

    \I__3980\ : Odrv4
    port map (
            O => \N__18099\,
            I => \c0.data_in_2_Z0Z_6\
        );

    \I__3979\ : InMux
    port map (
            O => \N__18092\,
            I => \N__18089\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__18086\,
            I => \N__18080\
        );

    \I__3976\ : InMux
    port map (
            O => \N__18085\,
            I => \N__18073\
        );

    \I__3975\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18073\
        );

    \I__3974\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18073\
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__18080\,
            I => \c0.d_4_22\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__18073\,
            I => \c0.d_4_22\
        );

    \I__3971\ : CascadeMux
    port map (
            O => \N__18068\,
            I => \c0.d_4_RNI9LFUVZ0Z_43_cascade_\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__18065\,
            I => \c0.wait_for_transmission_RNI9PP5BZ0Z1_cascade_\
        );

    \I__3969\ : InMux
    port map (
            O => \N__18062\,
            I => \N__18059\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__18059\,
            I => \N__18056\
        );

    \I__3967\ : Span4Mux_v
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__3966\ : Odrv4
    port map (
            O => \N__18053\,
            I => \c0.un1_data_in_6__1_1\
        );

    \I__3965\ : InMux
    port map (
            O => \N__18050\,
            I => \N__18047\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__18047\,
            I => \c0.g0_2_3\
        );

    \I__3963\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18041\,
            I => \N__18037\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__18040\,
            I => \N__18032\
        );

    \I__3960\ : Span4Mux_v
    port map (
            O => \N__18037\,
            I => \N__18029\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18036\,
            I => \N__18026\
        );

    \I__3958\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18021\
        );

    \I__3957\ : InMux
    port map (
            O => \N__18032\,
            I => \N__18021\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__18029\,
            I => \c0.d_4_23\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__18026\,
            I => \c0.d_4_23\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__18021\,
            I => \c0.d_4_23\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__18014\,
            I => \c0.N_126_cascade_\
        );

    \I__3952\ : InMux
    port map (
            O => \N__18011\,
            I => \N__18008\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__18008\,
            I => \c0.un1_data_in_6__1\
        );

    \I__3950\ : InMux
    port map (
            O => \N__18005\,
            I => \N__18000\
        );

    \I__3949\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17996\
        );

    \I__3948\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17992\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__18000\,
            I => \N__17988\
        );

    \I__3946\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17985\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__17996\,
            I => \N__17982\
        );

    \I__3944\ : InMux
    port map (
            O => \N__17995\,
            I => \N__17979\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__17992\,
            I => \N__17976\
        );

    \I__3942\ : InMux
    port map (
            O => \N__17991\,
            I => \N__17973\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__17988\,
            I => \c0.d_4_35\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__17985\,
            I => \c0.d_4_35\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__17982\,
            I => \c0.d_4_35\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__17979\,
            I => \c0.d_4_35\
        );

    \I__3937\ : Odrv4
    port map (
            O => \N__17976\,
            I => \c0.d_4_35\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__17973\,
            I => \c0.d_4_35\
        );

    \I__3935\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17957\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__17957\,
            I => \N__17953\
        );

    \I__3933\ : InMux
    port map (
            O => \N__17956\,
            I => \N__17950\
        );

    \I__3932\ : Odrv12
    port map (
            O => \N__17953\,
            I => \c0.data_in_0_Z0Z_7\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__17950\,
            I => \c0.data_in_0_Z0Z_7\
        );

    \I__3930\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17942\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17942\,
            I => \N__17938\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__17941\,
            I => \N__17934\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__17938\,
            I => \N__17931\
        );

    \I__3926\ : InMux
    port map (
            O => \N__17937\,
            I => \N__17926\
        );

    \I__3925\ : InMux
    port map (
            O => \N__17934\,
            I => \N__17926\
        );

    \I__3924\ : Odrv4
    port map (
            O => \N__17931\,
            I => \c0.d_4_15\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__17926\,
            I => \c0.d_4_15\
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__17921\,
            I => \c0.data_in_frame_1__m_7_cascade_\
        );

    \I__3921\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17914\
        );

    \I__3920\ : InMux
    port map (
            O => \N__17917\,
            I => \N__17911\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__17914\,
            I => \N__17906\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__17911\,
            I => \N__17906\
        );

    \I__3917\ : Span4Mux_h
    port map (
            O => \N__17906\,
            I => \N__17897\
        );

    \I__3916\ : InMux
    port map (
            O => \N__17905\,
            I => \N__17890\
        );

    \I__3915\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17890\
        );

    \I__3914\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17890\
        );

    \I__3913\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17883\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17883\
        );

    \I__3911\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17883\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__17897\,
            I => \c0.d_4_31\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__17890\,
            I => \c0.d_4_31\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__17883\,
            I => \c0.d_4_31\
        );

    \I__3907\ : InMux
    port map (
            O => \N__17876\,
            I => \N__17873\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__17873\,
            I => \c0.tx2_data_1_iv_1_7\
        );

    \I__3905\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17866\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__17869\,
            I => \N__17862\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__17866\,
            I => \N__17859\
        );

    \I__3902\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17851\
        );

    \I__3901\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17851\
        );

    \I__3900\ : Span4Mux_h
    port map (
            O => \N__17859\,
            I => \N__17847\
        );

    \I__3899\ : CascadeMux
    port map (
            O => \N__17858\,
            I => \N__17844\
        );

    \I__3898\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17839\
        );

    \I__3897\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17839\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__17851\,
            I => \N__17836\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__17850\,
            I => \N__17832\
        );

    \I__3894\ : Span4Mux_h
    port map (
            O => \N__17847\,
            I => \N__17829\
        );

    \I__3893\ : InMux
    port map (
            O => \N__17844\,
            I => \N__17826\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__17839\,
            I => \N__17821\
        );

    \I__3891\ : Span12Mux_v
    port map (
            O => \N__17836\,
            I => \N__17821\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17816\
        );

    \I__3889\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17816\
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__17829\,
            I => \c0.N_205\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__17826\,
            I => \c0.N_205\
        );

    \I__3886\ : Odrv12
    port map (
            O => \N__17821\,
            I => \c0.N_205\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__17816\,
            I => \c0.N_205\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17804\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__17804\,
            I => \N__17801\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__17801\,
            I => \N__17795\
        );

    \I__3881\ : InMux
    port map (
            O => \N__17800\,
            I => \N__17790\
        );

    \I__3880\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17790\
        );

    \I__3879\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17787\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__17795\,
            I => \c0.d_4_27\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__17790\,
            I => \c0.d_4_27\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__17787\,
            I => \c0.d_4_27\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__17780\,
            I => \c0.N_205_cascade_\
        );

    \I__3874\ : InMux
    port map (
            O => \N__17777\,
            I => \N__17774\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__17774\,
            I => \N__17771\
        );

    \I__3872\ : Span4Mux_h
    port map (
            O => \N__17771\,
            I => \N__17767\
        );

    \I__3871\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17764\
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__17767\,
            I => \c0.d_4_11\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__17764\,
            I => \c0.d_4_11\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17759\,
            I => \N__17756\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__17753\,
            I => \N__17750\
        );

    \I__3865\ : Span4Mux_h
    port map (
            O => \N__17750\,
            I => \N__17747\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__17747\,
            I => \c0.tx2_data_1_iv_4_1_3\
        );

    \I__3863\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17740\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__17743\,
            I => \N__17737\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__17740\,
            I => \N__17734\
        );

    \I__3860\ : InMux
    port map (
            O => \N__17737\,
            I => \N__17731\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__17734\,
            I => \c0.un1_data_in_6__5\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__17731\,
            I => \c0.un1_data_in_6__5\
        );

    \I__3857\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17721\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17718\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17715\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__17721\,
            I => \N__17712\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__17718\,
            I => \c0.i12_THRU_CO\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__17715\,
            I => \c0.i12_THRU_CO\
        );

    \I__3851\ : Odrv12
    port map (
            O => \N__17712\,
            I => \c0.i12_THRU_CO\
        );

    \I__3850\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17701\
        );

    \I__3849\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17698\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__17701\,
            I => \c0.N_136\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__17698\,
            I => \c0.N_136\
        );

    \I__3846\ : InMux
    port map (
            O => \N__17693\,
            I => \N__17688\
        );

    \I__3845\ : InMux
    port map (
            O => \N__17692\,
            I => \N__17685\
        );

    \I__3844\ : InMux
    port map (
            O => \N__17691\,
            I => \N__17682\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17688\,
            I => \N__17679\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17685\,
            I => \N__17676\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__17682\,
            I => \N__17673\
        );

    \I__3840\ : Span4Mux_v
    port map (
            O => \N__17679\,
            I => \N__17670\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__17676\,
            I => \c0.wait_for_transmission4_13_1\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__17673\,
            I => \c0.wait_for_transmission4_13_1\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__17670\,
            I => \c0.wait_for_transmission4_13_1\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__17663\,
            I => \c0.g1_3_cascade_\
        );

    \I__3835\ : InMux
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__17657\,
            I => \N__17654\
        );

    \I__3833\ : Span4Mux_v
    port map (
            O => \N__17654\,
            I => \N__17650\
        );

    \I__3832\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17647\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__17650\,
            I => \N__17642\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__17647\,
            I => \N__17642\
        );

    \I__3829\ : Sp12to4
    port map (
            O => \N__17642\,
            I => \N__17639\
        );

    \I__3828\ : Odrv12
    port map (
            O => \N__17639\,
            I => \c0.un1_data_in_7__0_0_a2_1_a2_5_0\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__17636\,
            I => \c0.i12_7_c_RNIP740G_cascade_\
        );

    \I__3826\ : InMux
    port map (
            O => \N__17633\,
            I => \N__17630\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__17630\,
            I => \c0.g1_2\
        );

    \I__3824\ : InMux
    port map (
            O => \N__17627\,
            I => \N__17624\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__17624\,
            I => \N__17621\
        );

    \I__3822\ : Span4Mux_v
    port map (
            O => \N__17621\,
            I => \N__17617\
        );

    \I__3821\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17614\
        );

    \I__3820\ : Odrv4
    port map (
            O => \N__17617\,
            I => \c0.wait_for_transmission4_12_5\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__17614\,
            I => \c0.wait_for_transmission4_12_5\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17609\,
            I => \N__17606\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__17606\,
            I => \N__17602\
        );

    \I__3816\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17599\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__17602\,
            I => \N__17596\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__17599\,
            I => \c0.un1_data_in_7__3_i\
        );

    \I__3813\ : Odrv4
    port map (
            O => \N__17596\,
            I => \c0.un1_data_in_7__3_i\
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__17591\,
            I => \c0.g1_5_cascade_\
        );

    \I__3811\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17584\
        );

    \I__3810\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17581\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__17584\,
            I => \N__17578\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__17581\,
            I => \c0.wait_for_transmission4_12_4\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__17578\,
            I => \c0.wait_for_transmission4_12_4\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17570\,
            I => \c0.byte_transmit_counterZ0Z_4\
        );

    \I__3804\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17558\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17555\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17550\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17547\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17544\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17541\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17561\,
            I => \N__17537\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__17558\,
            I => \N__17534\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__17555\,
            I => \N__17531\
        );

    \I__3795\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17528\
        );

    \I__3794\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17525\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__17550\,
            I => \N__17522\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__17547\,
            I => \N__17517\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__17544\,
            I => \N__17512\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__17541\,
            I => \N__17512\
        );

    \I__3789\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17509\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17506\
        );

    \I__3787\ : Span4Mux_v
    port map (
            O => \N__17534\,
            I => \N__17492\
        );

    \I__3786\ : Span4Mux_v
    port map (
            O => \N__17531\,
            I => \N__17492\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17528\,
            I => \N__17492\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__17525\,
            I => \N__17492\
        );

    \I__3783\ : Span4Mux_v
    port map (
            O => \N__17522\,
            I => \N__17492\
        );

    \I__3782\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17489\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17486\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__17517\,
            I => \N__17483\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__17512\,
            I => \N__17476\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__17509\,
            I => \N__17476\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__17506\,
            I => \N__17476\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17505\,
            I => \N__17470\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17470\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17467\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__17492\,
            I => \N__17462\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17489\,
            I => \N__17462\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17486\,
            I => \N__17455\
        );

    \I__3770\ : Span4Mux_h
    port map (
            O => \N__17483\,
            I => \N__17455\
        );

    \I__3769\ : Span4Mux_h
    port map (
            O => \N__17476\,
            I => \N__17455\
        );

    \I__3768\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17452\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__17470\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__17467\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__17462\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__17455\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__17452\,
            I => \c0.byte_transmit_counterZ0Z_0\
        );

    \I__3762\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17438\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__17438\,
            I => \c0.un144_newcrc_3\
        );

    \I__3760\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17430\
        );

    \I__3759\ : InMux
    port map (
            O => \N__17434\,
            I => \N__17427\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17433\,
            I => \N__17424\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__17430\,
            I => \N__17419\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__17427\,
            I => \N__17419\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__17424\,
            I => \N__17415\
        );

    \I__3754\ : Span4Mux_h
    port map (
            O => \N__17419\,
            I => \N__17412\
        );

    \I__3753\ : InMux
    port map (
            O => \N__17418\,
            I => \N__17409\
        );

    \I__3752\ : Odrv12
    port map (
            O => \N__17415\,
            I => \c0.d_2_34\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__17412\,
            I => \c0.d_2_34\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__17409\,
            I => \c0.d_2_34\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__17396\,
            I => \c0.un144_newcrc_4\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17393\,
            I => \N__17389\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__17392\,
            I => \N__17386\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__17389\,
            I => \N__17383\
        );

    \I__3743\ : InMux
    port map (
            O => \N__17386\,
            I => \N__17380\
        );

    \I__3742\ : Span4Mux_v
    port map (
            O => \N__17383\,
            I => \N__17373\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__17380\,
            I => \N__17373\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17379\,
            I => \N__17370\
        );

    \I__3739\ : InMux
    port map (
            O => \N__17378\,
            I => \N__17367\
        );

    \I__3738\ : Span4Mux_h
    port map (
            O => \N__17373\,
            I => \N__17362\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__17370\,
            I => \N__17362\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__17367\,
            I => \c0.d_2_33\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__17362\,
            I => \c0.d_2_33\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17357\,
            I => \N__17354\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__17354\,
            I => \N__17351\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__17351\,
            I => \c0.data_out_7_Z0Z_6\
        );

    \I__3731\ : SRMux
    port map (
            O => \N__17348\,
            I => \N__17334\
        );

    \I__3730\ : SRMux
    port map (
            O => \N__17347\,
            I => \N__17331\
        );

    \I__3729\ : SRMux
    port map (
            O => \N__17346\,
            I => \N__17328\
        );

    \I__3728\ : SRMux
    port map (
            O => \N__17345\,
            I => \N__17325\
        );

    \I__3727\ : SRMux
    port map (
            O => \N__17344\,
            I => \N__17322\
        );

    \I__3726\ : SRMux
    port map (
            O => \N__17343\,
            I => \N__17319\
        );

    \I__3725\ : SRMux
    port map (
            O => \N__17342\,
            I => \N__17316\
        );

    \I__3724\ : SRMux
    port map (
            O => \N__17341\,
            I => \N__17313\
        );

    \I__3723\ : SRMux
    port map (
            O => \N__17340\,
            I => \N__17310\
        );

    \I__3722\ : SRMux
    port map (
            O => \N__17339\,
            I => \N__17307\
        );

    \I__3721\ : SRMux
    port map (
            O => \N__17338\,
            I => \N__17304\
        );

    \I__3720\ : SRMux
    port map (
            O => \N__17337\,
            I => \N__17301\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17334\,
            I => \N__17284\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__17331\,
            I => \N__17281\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__17328\,
            I => \N__17278\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__17325\,
            I => \N__17275\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__17322\,
            I => \N__17272\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17269\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__17316\,
            I => \N__17266\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__17313\,
            I => \N__17263\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__17310\,
            I => \N__17260\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__17307\,
            I => \N__17257\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__17304\,
            I => \N__17254\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__17301\,
            I => \N__17251\
        );

    \I__3707\ : CEMux
    port map (
            O => \N__17300\,
            I => \N__17198\
        );

    \I__3706\ : CEMux
    port map (
            O => \N__17299\,
            I => \N__17198\
        );

    \I__3705\ : CEMux
    port map (
            O => \N__17298\,
            I => \N__17198\
        );

    \I__3704\ : CEMux
    port map (
            O => \N__17297\,
            I => \N__17198\
        );

    \I__3703\ : CEMux
    port map (
            O => \N__17296\,
            I => \N__17198\
        );

    \I__3702\ : CEMux
    port map (
            O => \N__17295\,
            I => \N__17198\
        );

    \I__3701\ : CEMux
    port map (
            O => \N__17294\,
            I => \N__17198\
        );

    \I__3700\ : CEMux
    port map (
            O => \N__17293\,
            I => \N__17198\
        );

    \I__3699\ : CEMux
    port map (
            O => \N__17292\,
            I => \N__17198\
        );

    \I__3698\ : CEMux
    port map (
            O => \N__17291\,
            I => \N__17198\
        );

    \I__3697\ : CEMux
    port map (
            O => \N__17290\,
            I => \N__17198\
        );

    \I__3696\ : CEMux
    port map (
            O => \N__17289\,
            I => \N__17198\
        );

    \I__3695\ : CEMux
    port map (
            O => \N__17288\,
            I => \N__17198\
        );

    \I__3694\ : CEMux
    port map (
            O => \N__17287\,
            I => \N__17198\
        );

    \I__3693\ : Glb2LocalMux
    port map (
            O => \N__17284\,
            I => \N__17198\
        );

    \I__3692\ : Glb2LocalMux
    port map (
            O => \N__17281\,
            I => \N__17198\
        );

    \I__3691\ : Glb2LocalMux
    port map (
            O => \N__17278\,
            I => \N__17198\
        );

    \I__3690\ : Glb2LocalMux
    port map (
            O => \N__17275\,
            I => \N__17198\
        );

    \I__3689\ : Glb2LocalMux
    port map (
            O => \N__17272\,
            I => \N__17198\
        );

    \I__3688\ : Glb2LocalMux
    port map (
            O => \N__17269\,
            I => \N__17198\
        );

    \I__3687\ : Glb2LocalMux
    port map (
            O => \N__17266\,
            I => \N__17198\
        );

    \I__3686\ : Glb2LocalMux
    port map (
            O => \N__17263\,
            I => \N__17198\
        );

    \I__3685\ : Glb2LocalMux
    port map (
            O => \N__17260\,
            I => \N__17198\
        );

    \I__3684\ : Glb2LocalMux
    port map (
            O => \N__17257\,
            I => \N__17198\
        );

    \I__3683\ : Glb2LocalMux
    port map (
            O => \N__17254\,
            I => \N__17198\
        );

    \I__3682\ : Glb2LocalMux
    port map (
            O => \N__17251\,
            I => \N__17198\
        );

    \I__3681\ : GlobalMux
    port map (
            O => \N__17198\,
            I => \N__17195\
        );

    \I__3680\ : gio2CtrlBuf
    port map (
            O => \N__17195\,
            I => \c0.data_out_0__1_sqmuxa_g\
        );

    \I__3679\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__17189\,
            I => \N__17185\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17188\,
            I => \N__17181\
        );

    \I__3676\ : Span4Mux_v
    port map (
            O => \N__17185\,
            I => \N__17175\
        );

    \I__3675\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17172\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__17181\,
            I => \N__17168\
        );

    \I__3673\ : InMux
    port map (
            O => \N__17180\,
            I => \N__17161\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17161\
        );

    \I__3671\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17161\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__17175\,
            I => \N__17158\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__17172\,
            I => \N__17155\
        );

    \I__3668\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17152\
        );

    \I__3667\ : Span4Mux_h
    port map (
            O => \N__17168\,
            I => \N__17147\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__17161\,
            I => \N__17147\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__17158\,
            I => \c0.d_4_12\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__17155\,
            I => \c0.d_4_12\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17152\,
            I => \c0.d_4_12\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__17147\,
            I => \c0.d_4_12\
        );

    \I__3661\ : InMux
    port map (
            O => \N__17138\,
            I => \N__17135\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__17135\,
            I => \N__17132\
        );

    \I__3659\ : Span4Mux_h
    port map (
            O => \N__17132\,
            I => \N__17129\
        );

    \I__3658\ : Span4Mux_v
    port map (
            O => \N__17129\,
            I => \N__17122\
        );

    \I__3657\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17119\
        );

    \I__3656\ : InMux
    port map (
            O => \N__17127\,
            I => \N__17116\
        );

    \I__3655\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17111\
        );

    \I__3654\ : InMux
    port map (
            O => \N__17125\,
            I => \N__17111\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__17122\,
            I => \c0.d_4_44\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__17119\,
            I => \c0.d_4_44\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__17116\,
            I => \c0.d_4_44\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__17111\,
            I => \c0.d_4_44\
        );

    \I__3649\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17099\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__17099\,
            I => \N__17096\
        );

    \I__3647\ : Odrv12
    port map (
            O => \N__17096\,
            I => \c0.tx2_data_1_iv_5_7\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__17093\,
            I => \N__17090\
        );

    \I__3645\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17087\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__17087\,
            I => \N__17084\
        );

    \I__3643\ : Odrv12
    port map (
            O => \N__17084\,
            I => \c0.tx2_data_1_0_i_1_7\
        );

    \I__3642\ : InMux
    port map (
            O => \N__17081\,
            I => \N__17078\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__17078\,
            I => \N__17075\
        );

    \I__3640\ : Span4Mux_h
    port map (
            O => \N__17075\,
            I => \N__17072\
        );

    \I__3639\ : Span4Mux_v
    port map (
            O => \N__17072\,
            I => \N__17069\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__17069\,
            I => \c0.tx2.r_Tx_DataZ0Z_7\
        );

    \I__3637\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17063\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__17063\,
            I => \N__17059\
        );

    \I__3635\ : InMux
    port map (
            O => \N__17062\,
            I => \N__17056\
        );

    \I__3634\ : Span4Mux_h
    port map (
            O => \N__17059\,
            I => \N__17050\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__17056\,
            I => \N__17050\
        );

    \I__3632\ : InMux
    port map (
            O => \N__17055\,
            I => \N__17047\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__17050\,
            I => \c0.d_4_13\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__17047\,
            I => \c0.d_4_13\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__17039\,
            I => \N__17036\
        );

    \I__3627\ : Span4Mux_h
    port map (
            O => \N__17036\,
            I => \N__17032\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17029\
        );

    \I__3625\ : Span4Mux_h
    port map (
            O => \N__17032\,
            I => \N__17024\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__17029\,
            I => \N__17024\
        );

    \I__3623\ : Span4Mux_v
    port map (
            O => \N__17024\,
            I => \N__17019\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__17023\,
            I => \N__17016\
        );

    \I__3621\ : InMux
    port map (
            O => \N__17022\,
            I => \N__17012\
        );

    \I__3620\ : Span4Mux_h
    port map (
            O => \N__17019\,
            I => \N__17009\
        );

    \I__3619\ : InMux
    port map (
            O => \N__17016\,
            I => \N__17004\
        );

    \I__3618\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17004\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__17012\,
            I => \c0.d_4_29\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__17009\,
            I => \c0.d_4_29\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__17004\,
            I => \c0.d_4_29\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__16997\,
            I => \c0.data_in_frame_1__m_5_cascade_\
        );

    \I__3613\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__16988\,
            I => \c0.tx2_data_1_0_i_1_5\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__16985\,
            I => \c0.tx2_data_1_iv_1_5_cascade_\
        );

    \I__3609\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__16979\,
            I => \N__16976\
        );

    \I__3607\ : Span4Mux_v
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__3606\ : Span4Mux_v
    port map (
            O => \N__16973\,
            I => \N__16970\
        );

    \I__3605\ : Odrv4
    port map (
            O => \N__16970\,
            I => \c0.tx2.r_Tx_DataZ0Z_5\
        );

    \I__3604\ : InMux
    port map (
            O => \N__16967\,
            I => \N__16964\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__16964\,
            I => \c0.data_out_6_Z0Z_6\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__16961\,
            I => \c0.N_4_0_cascade_\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__16955\,
            I => \N__16952\
        );

    \I__3599\ : Odrv12
    port map (
            O => \N__16952\,
            I => \c0.N_197\
        );

    \I__3598\ : IoInMux
    port map (
            O => \N__16949\,
            I => \N__16946\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__16946\,
            I => \N__16943\
        );

    \I__3596\ : IoSpan4Mux
    port map (
            O => \N__16943\,
            I => \N__16940\
        );

    \I__3595\ : Span4Mux_s1_v
    port map (
            O => \N__16940\,
            I => \N__16937\
        );

    \I__3594\ : Span4Mux_v
    port map (
            O => \N__16937\,
            I => \N__16934\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__16934\,
            I => \c0.data_out_0__1_sqmuxa\
        );

    \I__3592\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__16928\,
            I => \c0.byte_transmit_counterZ0Z_6\
        );

    \I__3590\ : InMux
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__16922\,
            I => \c0.byte_transmit_counterZ0Z_3\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__16919\,
            I => \c0.m2_e_1_cascade_\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__16916\,
            I => \c0.N_129_mux_cascade_\
        );

    \I__3586\ : InMux
    port map (
            O => \N__16913\,
            I => \N__16910\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__16910\,
            I => \N__16905\
        );

    \I__3584\ : InMux
    port map (
            O => \N__16909\,
            I => \N__16902\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16899\
        );

    \I__3582\ : Span4Mux_h
    port map (
            O => \N__16905\,
            I => \N__16894\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16902\,
            I => \N__16894\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__16899\,
            I => \N__16891\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__16894\,
            I => \N__16888\
        );

    \I__3578\ : Odrv12
    port map (
            O => \N__16891\,
            I => \c0.N_86\
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__16888\,
            I => \c0.N_86\
        );

    \I__3576\ : InMux
    port map (
            O => \N__16883\,
            I => \N__16878\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__16882\,
            I => \N__16872\
        );

    \I__3574\ : InMux
    port map (
            O => \N__16881\,
            I => \N__16864\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__16878\,
            I => \N__16861\
        );

    \I__3572\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16856\
        );

    \I__3571\ : InMux
    port map (
            O => \N__16876\,
            I => \N__16856\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16875\,
            I => \N__16851\
        );

    \I__3569\ : InMux
    port map (
            O => \N__16872\,
            I => \N__16851\
        );

    \I__3568\ : InMux
    port map (
            O => \N__16871\,
            I => \N__16844\
        );

    \I__3567\ : InMux
    port map (
            O => \N__16870\,
            I => \N__16844\
        );

    \I__3566\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16844\
        );

    \I__3565\ : InMux
    port map (
            O => \N__16868\,
            I => \N__16839\
        );

    \I__3564\ : InMux
    port map (
            O => \N__16867\,
            I => \N__16836\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__16864\,
            I => \N__16833\
        );

    \I__3562\ : Span4Mux_v
    port map (
            O => \N__16861\,
            I => \N__16828\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__16856\,
            I => \N__16828\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__16851\,
            I => \N__16825\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__16844\,
            I => \N__16822\
        );

    \I__3558\ : InMux
    port map (
            O => \N__16843\,
            I => \N__16819\
        );

    \I__3557\ : InMux
    port map (
            O => \N__16842\,
            I => \N__16816\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__16839\,
            I => \N__16813\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__16836\,
            I => \N__16810\
        );

    \I__3554\ : Span4Mux_v
    port map (
            O => \N__16833\,
            I => \N__16800\
        );

    \I__3553\ : Span4Mux_v
    port map (
            O => \N__16828\,
            I => \N__16800\
        );

    \I__3552\ : Span4Mux_v
    port map (
            O => \N__16825\,
            I => \N__16800\
        );

    \I__3551\ : Sp12to4
    port map (
            O => \N__16822\,
            I => \N__16795\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__16819\,
            I => \N__16795\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__16816\,
            I => \N__16788\
        );

    \I__3548\ : Span4Mux_h
    port map (
            O => \N__16813\,
            I => \N__16788\
        );

    \I__3547\ : Span4Mux_v
    port map (
            O => \N__16810\,
            I => \N__16788\
        );

    \I__3546\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16783\
        );

    \I__3545\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16783\
        );

    \I__3544\ : InMux
    port map (
            O => \N__16807\,
            I => \N__16778\
        );

    \I__3543\ : Span4Mux_h
    port map (
            O => \N__16800\,
            I => \N__16775\
        );

    \I__3542\ : Span12Mux_s7_v
    port map (
            O => \N__16795\,
            I => \N__16768\
        );

    \I__3541\ : Sp12to4
    port map (
            O => \N__16788\,
            I => \N__16768\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__16783\,
            I => \N__16768\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16763\
        );

    \I__3538\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16763\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__16778\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3536\ : Odrv4
    port map (
            O => \N__16775\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3535\ : Odrv12
    port map (
            O => \N__16768\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__16763\,
            I => \c0.byte_transmit_counterZ0Z_1\
        );

    \I__3533\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16751\,
            I => \N__16748\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__16748\,
            I => \c0.data_in_frame_6_Z0Z_0\
        );

    \I__3530\ : InMux
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__16742\,
            I => \N__16738\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__16741\,
            I => \N__16734\
        );

    \I__3527\ : Span4Mux_v
    port map (
            O => \N__16738\,
            I => \N__16731\
        );

    \I__3526\ : InMux
    port map (
            O => \N__16737\,
            I => \N__16726\
        );

    \I__3525\ : InMux
    port map (
            O => \N__16734\,
            I => \N__16726\
        );

    \I__3524\ : Odrv4
    port map (
            O => \N__16731\,
            I => \c0.data_in_3_Z0Z_2\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__16726\,
            I => \c0.data_in_3_Z0Z_2\
        );

    \I__3522\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16718\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__16718\,
            I => \N__16712\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16709\
        );

    \I__3519\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16703\
        );

    \I__3518\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16703\
        );

    \I__3517\ : Span4Mux_v
    port map (
            O => \N__16712\,
            I => \N__16698\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__16709\,
            I => \N__16698\
        );

    \I__3515\ : InMux
    port map (
            O => \N__16708\,
            I => \N__16695\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__16703\,
            I => \N__16692\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__16698\,
            I => \N__16688\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__16695\,
            I => \N__16685\
        );

    \I__3511\ : Span4Mux_h
    port map (
            O => \N__16692\,
            I => \N__16682\
        );

    \I__3510\ : InMux
    port map (
            O => \N__16691\,
            I => \N__16679\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__16688\,
            I => \c0.d_4_26\
        );

    \I__3508\ : Odrv12
    port map (
            O => \N__16685\,
            I => \c0.d_4_26\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__16682\,
            I => \c0.d_4_26\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__16679\,
            I => \c0.d_4_26\
        );

    \I__3505\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__3503\ : Span4Mux_h
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__3502\ : Span4Mux_h
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__16658\,
            I => \c0.data_in_frame_6_Z0Z_1\
        );

    \I__3500\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3498\ : Span4Mux_h
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3497\ : Span4Mux_h
    port map (
            O => \N__16646\,
            I => \N__16641\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16638\
        );

    \I__3495\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16635\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__16641\,
            I => \c0.data_in_1_Z0Z_2\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__16638\,
            I => \c0.data_in_1_Z0Z_2\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__16635\,
            I => \c0.data_in_1_Z0Z_2\
        );

    \I__3491\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16624\
        );

    \I__3490\ : CascadeMux
    port map (
            O => \N__16627\,
            I => \N__16621\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__16624\,
            I => \N__16616\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16621\,
            I => \N__16612\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16620\,
            I => \N__16607\
        );

    \I__3486\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16607\
        );

    \I__3485\ : Span4Mux_v
    port map (
            O => \N__16616\,
            I => \N__16604\
        );

    \I__3484\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16601\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16612\,
            I => \N__16598\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__16607\,
            I => \N__16595\
        );

    \I__3481\ : Span4Mux_h
    port map (
            O => \N__16604\,
            I => \N__16588\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__16601\,
            I => \N__16588\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__16598\,
            I => \N__16588\
        );

    \I__3478\ : Odrv12
    port map (
            O => \N__16595\,
            I => \c0.d_4_10\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__16588\,
            I => \c0.d_4_10\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__3475\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__16577\,
            I => \N__16574\
        );

    \I__3473\ : Span4Mux_h
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__16571\,
            I => \c0.data_in_frame_7_Z0Z_0\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16563\
        );

    \I__3470\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16560\
        );

    \I__3469\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16557\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__16563\,
            I => \N__16554\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__16560\,
            I => \N__16551\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__16557\,
            I => \N__16548\
        );

    \I__3465\ : Span4Mux_v
    port map (
            O => \N__16554\,
            I => \N__16545\
        );

    \I__3464\ : Sp12to4
    port map (
            O => \N__16551\,
            I => \N__16542\
        );

    \I__3463\ : Span4Mux_h
    port map (
            O => \N__16548\,
            I => \N__16538\
        );

    \I__3462\ : Sp12to4
    port map (
            O => \N__16545\,
            I => \N__16533\
        );

    \I__3461\ : Span12Mux_v
    port map (
            O => \N__16542\,
            I => \N__16533\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16541\,
            I => \N__16530\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__16538\,
            I => \c0.d_2_36\
        );

    \I__3458\ : Odrv12
    port map (
            O => \N__16533\,
            I => \c0.d_2_36\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__16530\,
            I => \c0.d_2_36\
        );

    \I__3456\ : InMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__3454\ : Span4Mux_v
    port map (
            O => \N__16517\,
            I => \N__16512\
        );

    \I__3453\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16509\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16506\
        );

    \I__3451\ : Span4Mux_h
    port map (
            O => \N__16512\,
            I => \N__16501\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__16509\,
            I => \N__16501\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__16506\,
            I => \N__16498\
        );

    \I__3448\ : Span4Mux_h
    port map (
            O => \N__16501\,
            I => \N__16495\
        );

    \I__3447\ : Span4Mux_h
    port map (
            O => \N__16498\,
            I => \N__16491\
        );

    \I__3446\ : Span4Mux_v
    port map (
            O => \N__16495\,
            I => \N__16488\
        );

    \I__3445\ : InMux
    port map (
            O => \N__16494\,
            I => \N__16485\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__16491\,
            I => \c0.d_2_35\
        );

    \I__3443\ : Odrv4
    port map (
            O => \N__16488\,
            I => \c0.d_2_35\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__16485\,
            I => \c0.d_2_35\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__3440\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16472\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__16472\,
            I => \N__16469\
        );

    \I__3438\ : Span4Mux_h
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__16466\,
            I => \c0.N_71\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__16463\,
            I => \N__16458\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16462\,
            I => \N__16454\
        );

    \I__3434\ : InMux
    port map (
            O => \N__16461\,
            I => \N__16451\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16446\
        );

    \I__3432\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16446\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__16454\,
            I => \c0.tx2.r_Bit_IndexZ0Z_0\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__16451\,
            I => \c0.tx2.r_Bit_IndexZ0Z_0\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__16446\,
            I => \c0.tx2.r_Bit_IndexZ0Z_0\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16439\,
            I => \N__16429\
        );

    \I__3427\ : InMux
    port map (
            O => \N__16438\,
            I => \N__16424\
        );

    \I__3426\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16424\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16415\
        );

    \I__3424\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16415\
        );

    \I__3423\ : InMux
    port map (
            O => \N__16434\,
            I => \N__16408\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16408\
        );

    \I__3421\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16408\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__16429\,
            I => \N__16403\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__16424\,
            I => \N__16403\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16423\,
            I => \N__16400\
        );

    \I__3417\ : InMux
    port map (
            O => \N__16422\,
            I => \N__16393\
        );

    \I__3416\ : InMux
    port map (
            O => \N__16421\,
            I => \N__16393\
        );

    \I__3415\ : InMux
    port map (
            O => \N__16420\,
            I => \N__16393\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__16415\,
            I => \c0.tx2.r_Clock_Count12_THRU_CO\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__16408\,
            I => \c0.tx2.r_Clock_Count12_THRU_CO\
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__16403\,
            I => \c0.tx2.r_Clock_Count12_THRU_CO\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__16400\,
            I => \c0.tx2.r_Clock_Count12_THRU_CO\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__16393\,
            I => \c0.tx2.r_Clock_Count12_THRU_CO\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16382\,
            I => \N__16378\
        );

    \I__3408\ : InMux
    port map (
            O => \N__16381\,
            I => \N__16375\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__16378\,
            I => \c0.tx2.N_257\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__16375\,
            I => \c0.tx2.N_257\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__16370\,
            I => \c0.tx2.N_258_cascade_\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16362\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16359\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16356\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__16362\,
            I => \N__16353\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__16359\,
            I => \N__16341\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__16356\,
            I => \N__16341\
        );

    \I__3398\ : Span4Mux_h
    port map (
            O => \N__16353\,
            I => \N__16338\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16352\,
            I => \N__16331\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16351\,
            I => \N__16331\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16350\,
            I => \N__16331\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16349\,
            I => \N__16326\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16348\,
            I => \N__16326\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16321\
        );

    \I__3391\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16321\
        );

    \I__3390\ : Span4Mux_h
    port map (
            O => \N__16341\,
            I => \N__16318\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__16338\,
            I => \c0.tx2.r_SM_MainZ0Z_1\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__16331\,
            I => \c0.tx2.r_SM_MainZ0Z_1\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__16326\,
            I => \c0.tx2.r_SM_MainZ0Z_1\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__16321\,
            I => \c0.tx2.r_SM_MainZ0Z_1\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__16318\,
            I => \c0.tx2.r_SM_MainZ0Z_1\
        );

    \I__3384\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16293\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16293\
        );

    \I__3382\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16293\
        );

    \I__3381\ : InMux
    port map (
            O => \N__16304\,
            I => \N__16293\
        );

    \I__3380\ : InMux
    port map (
            O => \N__16303\,
            I => \N__16290\
        );

    \I__3379\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16287\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__16293\,
            I => \N__16284\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__16290\,
            I => \c0.tx2.r_Bit_IndexZ0Z_1\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16287\,
            I => \c0.tx2.r_Bit_IndexZ0Z_1\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__16284\,
            I => \c0.tx2.r_Bit_IndexZ0Z_1\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__16277\,
            I => \N__16274\
        );

    \I__3373\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16271\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__16271\,
            I => \c0.un1_data_in_7__7_0_a2_0_a2_2\
        );

    \I__3371\ : InMux
    port map (
            O => \N__16268\,
            I => \N__16265\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__16265\,
            I => \N__16262\
        );

    \I__3369\ : Span4Mux_h
    port map (
            O => \N__16262\,
            I => \N__16259\
        );

    \I__3368\ : Span4Mux_h
    port map (
            O => \N__16259\,
            I => \N__16255\
        );

    \I__3367\ : InMux
    port map (
            O => \N__16258\,
            I => \N__16252\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__16255\,
            I => \c0.data_in_0_Z0Z_5\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__16252\,
            I => \c0.data_in_0_Z0Z_5\
        );

    \I__3364\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__16244\,
            I => \N__16241\
        );

    \I__3362\ : Span4Mux_h
    port map (
            O => \N__16241\,
            I => \N__16238\
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__16238\,
            I => \c0.wait_for_transmission_RNOZ0Z_9\
        );

    \I__3360\ : InMux
    port map (
            O => \N__16235\,
            I => \N__16232\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__16232\,
            I => \N__16228\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__16231\,
            I => \N__16224\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__16228\,
            I => \N__16221\
        );

    \I__3356\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16218\
        );

    \I__3355\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16215\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__16221\,
            I => \c0.data_in_2_Z0Z_2\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16218\,
            I => \c0.data_in_2_Z0Z_2\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__16215\,
            I => \c0.data_in_2_Z0Z_2\
        );

    \I__3351\ : InMux
    port map (
            O => \N__16208\,
            I => \N__16205\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__16205\,
            I => \N__16202\
        );

    \I__3349\ : Span4Mux_h
    port map (
            O => \N__16202\,
            I => \N__16198\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__16201\,
            I => \N__16194\
        );

    \I__3347\ : Span4Mux_v
    port map (
            O => \N__16198\,
            I => \N__16191\
        );

    \I__3346\ : InMux
    port map (
            O => \N__16197\,
            I => \N__16186\
        );

    \I__3345\ : InMux
    port map (
            O => \N__16194\,
            I => \N__16186\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__16191\,
            I => \c0.data_in_2_Z0Z_4\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__16186\,
            I => \c0.data_in_2_Z0Z_4\
        );

    \I__3342\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16177\
        );

    \I__3341\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16174\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__16177\,
            I => \N__16171\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__16174\,
            I => \N__16168\
        );

    \I__3338\ : Span4Mux_h
    port map (
            O => \N__16171\,
            I => \N__16161\
        );

    \I__3337\ : Span4Mux_v
    port map (
            O => \N__16168\,
            I => \N__16161\
        );

    \I__3336\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16156\
        );

    \I__3335\ : InMux
    port map (
            O => \N__16166\,
            I => \N__16156\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__16161\,
            I => \c0.d_4_18\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__16156\,
            I => \c0.d_4_18\
        );

    \I__3332\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16147\
        );

    \I__3331\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16144\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__16147\,
            I => \N__16139\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__16144\,
            I => \N__16139\
        );

    \I__3328\ : Odrv12
    port map (
            O => \N__16139\,
            I => \c0.N_124\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__16136\,
            I => \c0.N_124_cascade_\
        );

    \I__3326\ : InMux
    port map (
            O => \N__16133\,
            I => \N__16129\
        );

    \I__3325\ : InMux
    port map (
            O => \N__16132\,
            I => \N__16126\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__16129\,
            I => \N__16121\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__16126\,
            I => \N__16118\
        );

    \I__3322\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16115\
        );

    \I__3321\ : InMux
    port map (
            O => \N__16124\,
            I => \N__16112\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__16121\,
            I => \c0.d_4_RNI21N6Z0Z_11\
        );

    \I__3319\ : Odrv4
    port map (
            O => \N__16118\,
            I => \c0.d_4_RNI21N6Z0Z_11\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__16115\,
            I => \c0.d_4_RNI21N6Z0Z_11\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__16112\,
            I => \c0.d_4_RNI21N6Z0Z_11\
        );

    \I__3316\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16100\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__16100\,
            I => \N__16096\
        );

    \I__3314\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16093\
        );

    \I__3313\ : Span4Mux_h
    port map (
            O => \N__16096\,
            I => \N__16090\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__16093\,
            I => \c0.d_4_RNIPF9J2Z0Z_37\
        );

    \I__3311\ : Odrv4
    port map (
            O => \N__16090\,
            I => \c0.d_4_RNIPF9J2Z0Z_37\
        );

    \I__3310\ : InMux
    port map (
            O => \N__16085\,
            I => \N__16082\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__16082\,
            I => \N__16079\
        );

    \I__3308\ : Span4Mux_v
    port map (
            O => \N__16079\,
            I => \N__16075\
        );

    \I__3307\ : InMux
    port map (
            O => \N__16078\,
            I => \N__16072\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__16075\,
            I => \c0.data_in_4_Z0Z_1\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__16072\,
            I => \c0.data_in_4_Z0Z_1\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__16067\,
            I => \N__16064\
        );

    \I__3303\ : InMux
    port map (
            O => \N__16064\,
            I => \N__16060\
        );

    \I__3302\ : InMux
    port map (
            O => \N__16063\,
            I => \N__16057\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__16060\,
            I => \N__16054\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__16057\,
            I => \N__16051\
        );

    \I__3299\ : Span4Mux_h
    port map (
            O => \N__16054\,
            I => \N__16044\
        );

    \I__3298\ : Span4Mux_h
    port map (
            O => \N__16051\,
            I => \N__16044\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16039\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16039\
        );

    \I__3295\ : Odrv4
    port map (
            O => \N__16044\,
            I => \c0.d_4_33\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__16039\,
            I => \c0.d_4_33\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__16034\,
            I => \c0.un1_data_in_6__3_0_a2_5_a2_2_cascade_\
        );

    \I__3292\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16026\
        );

    \I__3291\ : InMux
    port map (
            O => \N__16030\,
            I => \N__16022\
        );

    \I__3290\ : InMux
    port map (
            O => \N__16029\,
            I => \N__16019\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__16026\,
            I => \N__16015\
        );

    \I__3288\ : InMux
    port map (
            O => \N__16025\,
            I => \N__16012\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__16022\,
            I => \N__16007\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__16019\,
            I => \N__16007\
        );

    \I__3285\ : InMux
    port map (
            O => \N__16018\,
            I => \N__16004\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__16015\,
            I => \c0.d_4_25\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__16012\,
            I => \c0.d_4_25\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__16007\,
            I => \c0.d_4_25\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__16004\,
            I => \c0.d_4_25\
        );

    \I__3280\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15992\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__15992\,
            I => \N__15989\
        );

    \I__3278\ : Span4Mux_v
    port map (
            O => \N__15989\,
            I => \N__15986\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__15986\,
            I => \c0.un1_data_in_6__3\
        );

    \I__3276\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15980\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__15980\,
            I => \c0.un1_data_in_6__3_0_a2_5_a2_1\
        );

    \I__3274\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15973\
        );

    \I__3273\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15970\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__15973\,
            I => \N__15967\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__15970\,
            I => \N__15964\
        );

    \I__3270\ : Span4Mux_h
    port map (
            O => \N__15967\,
            I => \N__15961\
        );

    \I__3269\ : Span4Mux_h
    port map (
            O => \N__15964\,
            I => \N__15955\
        );

    \I__3268\ : Span4Mux_h
    port map (
            O => \N__15961\,
            I => \N__15955\
        );

    \I__3267\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15952\
        );

    \I__3266\ : Odrv4
    port map (
            O => \N__15955\,
            I => \c0.data_in_1_Z0Z_1\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__15952\,
            I => \c0.data_in_1_Z0Z_1\
        );

    \I__3264\ : InMux
    port map (
            O => \N__15947\,
            I => \N__15943\
        );

    \I__3263\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15940\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__15943\,
            I => \N__15936\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__15940\,
            I => \N__15933\
        );

    \I__3260\ : InMux
    port map (
            O => \N__15939\,
            I => \N__15930\
        );

    \I__3259\ : Span12Mux_v
    port map (
            O => \N__15936\,
            I => \N__15927\
        );

    \I__3258\ : Span4Mux_h
    port map (
            O => \N__15933\,
            I => \N__15922\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__15930\,
            I => \N__15922\
        );

    \I__3256\ : Odrv12
    port map (
            O => \N__15927\,
            I => \c0.data_in_2_Z0Z_7\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__15922\,
            I => \c0.data_in_2_Z0Z_7\
        );

    \I__3254\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15914\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__15914\,
            I => \N__15910\
        );

    \I__3252\ : InMux
    port map (
            O => \N__15913\,
            I => \N__15907\
        );

    \I__3251\ : Odrv12
    port map (
            O => \N__15910\,
            I => \c0.data_in_5_Z0Z_0\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__15907\,
            I => \c0.data_in_5_Z0Z_0\
        );

    \I__3249\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15899\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__15899\,
            I => \N__15895\
        );

    \I__3247\ : CascadeMux
    port map (
            O => \N__15898\,
            I => \N__15892\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__15895\,
            I => \N__15887\
        );

    \I__3245\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15884\
        );

    \I__3244\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15881\
        );

    \I__3243\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15878\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__15887\,
            I => \c0.d_4_40\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__15884\,
            I => \c0.d_4_40\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__15881\,
            I => \c0.d_4_40\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__15878\,
            I => \c0.d_4_40\
        );

    \I__3238\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15866\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15863\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__15863\,
            I => \N__15859\
        );

    \I__3235\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15856\
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__15859\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_4_1_0\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__15856\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_4_1_0\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15848\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__15848\,
            I => \N__15845\
        );

    \I__3230\ : Span4Mux_h
    port map (
            O => \N__15845\,
            I => \N__15841\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15838\
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__15841\,
            I => \c0.data_in_4_Z0Z_3\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__15838\,
            I => \c0.data_in_4_Z0Z_3\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__15833\,
            I => \c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_\
        );

    \I__3225\ : InMux
    port map (
            O => \N__15830\,
            I => \N__15827\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__15827\,
            I => \N__15824\
        );

    \I__3223\ : Odrv12
    port map (
            O => \N__15824\,
            I => \c0.g3_2\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__15821\,
            I => \c0.un1_data_in_6__6_0_a2_0_a2_3_cascade_\
        );

    \I__3221\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15815\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__15815\,
            I => \N__15812\
        );

    \I__3219\ : Span4Mux_h
    port map (
            O => \N__15812\,
            I => \N__15804\
        );

    \I__3218\ : InMux
    port map (
            O => \N__15811\,
            I => \N__15801\
        );

    \I__3217\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15798\
        );

    \I__3216\ : InMux
    port map (
            O => \N__15809\,
            I => \N__15791\
        );

    \I__3215\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15791\
        );

    \I__3214\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15791\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__15804\,
            I => \c0.N_128\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__15801\,
            I => \c0.N_128\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__15798\,
            I => \c0.N_128\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__15791\,
            I => \c0.N_128\
        );

    \I__3209\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15777\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15781\,
            I => \N__15774\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__15780\,
            I => \N__15771\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__15777\,
            I => \N__15768\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__15774\,
            I => \N__15765\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15762\
        );

    \I__3203\ : Span4Mux_h
    port map (
            O => \N__15768\,
            I => \N__15757\
        );

    \I__3202\ : Span4Mux_h
    port map (
            O => \N__15765\,
            I => \N__15752\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__15762\,
            I => \N__15752\
        );

    \I__3200\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15749\
        );

    \I__3199\ : InMux
    port map (
            O => \N__15760\,
            I => \N__15746\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__15757\,
            I => \c0.d_4_41\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__15752\,
            I => \c0.d_4_41\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__15749\,
            I => \c0.d_4_41\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__15746\,
            I => \c0.d_4_41\
        );

    \I__3194\ : CascadeMux
    port map (
            O => \N__15737\,
            I => \c0.un1_data_in_6__5_0_a2_5_a2_2_cascade_\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15734\,
            I => \N__15729\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15733\,
            I => \N__15724\
        );

    \I__3191\ : InMux
    port map (
            O => \N__15732\,
            I => \N__15724\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__15729\,
            I => \N__15720\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__15724\,
            I => \N__15717\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__15723\,
            I => \N__15714\
        );

    \I__3187\ : Span4Mux_v
    port map (
            O => \N__15720\,
            I => \N__15711\
        );

    \I__3186\ : Span4Mux_v
    port map (
            O => \N__15717\,
            I => \N__15708\
        );

    \I__3185\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15705\
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__15711\,
            I => \c0.N_132\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__15708\,
            I => \c0.N_132\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__15705\,
            I => \c0.N_132\
        );

    \I__3181\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15695\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__15695\,
            I => \N__15691\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15694\,
            I => \N__15688\
        );

    \I__3178\ : Odrv12
    port map (
            O => \N__15691\,
            I => \c0.un1_data_in_6__6_0_a2_0_a2_3\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__15688\,
            I => \c0.un1_data_in_6__6_0_a2_0_a2_3\
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__15683\,
            I => \c0.un1_data_in_6__5_cascade_\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15677\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__15677\,
            I => \N__15674\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__15674\,
            I => \c0.g0_2_0\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15671\,
            I => \N__15666\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15670\,
            I => \N__15661\
        );

    \I__3170\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15661\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__15666\,
            I => \N__15655\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__15661\,
            I => \N__15655\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15660\,
            I => \N__15652\
        );

    \I__3166\ : Span4Mux_h
    port map (
            O => \N__15655\,
            I => \N__15649\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__15652\,
            I => \c0.d_4_43\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__15649\,
            I => \c0.d_4_43\
        );

    \I__3163\ : InMux
    port map (
            O => \N__15644\,
            I => \N__15641\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__15641\,
            I => \c0.un1_data_in_7__0_0_a2_1_a2_2\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15635\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__15635\,
            I => \c0.un1_data_in_6__4\
        );

    \I__3159\ : CascadeMux
    port map (
            O => \N__15632\,
            I => \c0.wait_for_transmission4_12_5_1_cascade_\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15629\,
            I => \N__15625\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15622\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__15625\,
            I => \N__15619\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__15622\,
            I => \N__15613\
        );

    \I__3154\ : Span4Mux_h
    port map (
            O => \N__15619\,
            I => \N__15613\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15610\
        );

    \I__3152\ : Odrv4
    port map (
            O => \N__15613\,
            I => \c0.N_108\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__15610\,
            I => \c0.N_108\
        );

    \I__3150\ : InMux
    port map (
            O => \N__15605\,
            I => \N__15602\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__15602\,
            I => \N__15598\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15601\,
            I => \N__15590\
        );

    \I__3147\ : Span4Mux_h
    port map (
            O => \N__15598\,
            I => \N__15587\
        );

    \I__3146\ : InMux
    port map (
            O => \N__15597\,
            I => \N__15580\
        );

    \I__3145\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15580\
        );

    \I__3144\ : InMux
    port map (
            O => \N__15595\,
            I => \N__15580\
        );

    \I__3143\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15577\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15574\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__15590\,
            I => \c0.d_4_32\
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__15587\,
            I => \c0.d_4_32\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__15580\,
            I => \c0.d_4_32\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15577\,
            I => \c0.d_4_32\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__15574\,
            I => \c0.d_4_32\
        );

    \I__3136\ : InMux
    port map (
            O => \N__15563\,
            I => \N__15560\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__15560\,
            I => \c0.un1_data_in_7__6_0_a2_5_a2_2\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15554\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__15554\,
            I => \c0.wait_for_transmission_RNOZ0Z_11\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15551\,
            I => \N__15547\
        );

    \I__3131\ : InMux
    port map (
            O => \N__15550\,
            I => \N__15544\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__15547\,
            I => \N__15541\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__15544\,
            I => \N__15538\
        );

    \I__3128\ : Span4Mux_v
    port map (
            O => \N__15541\,
            I => \N__15533\
        );

    \I__3127\ : Span4Mux_h
    port map (
            O => \N__15538\,
            I => \N__15533\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__15533\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_4_1\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__15530\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_4_1_cascade_\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__15527\,
            I => \N__15521\
        );

    \I__3123\ : InMux
    port map (
            O => \N__15526\,
            I => \N__15518\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__15525\,
            I => \N__15515\
        );

    \I__3121\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15510\
        );

    \I__3120\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15510\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__15518\,
            I => \N__15507\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15515\,
            I => \N__15504\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__15510\,
            I => \c0.d_4_47\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__15507\,
            I => \c0.d_4_47\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__15504\,
            I => \c0.d_4_47\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__15494\,
            I => \N__15491\
        );

    \I__3112\ : Span4Mux_h
    port map (
            O => \N__15491\,
            I => \N__15487\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15484\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__15487\,
            I => \c0.N_125\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15484\,
            I => \c0.N_125\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__15476\,
            I => \N__15473\
        );

    \I__3106\ : Span4Mux_h
    port map (
            O => \N__15473\,
            I => \N__15469\
        );

    \I__3105\ : InMux
    port map (
            O => \N__15472\,
            I => \N__15466\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__15469\,
            I => \c0.data_in_0_Z0Z_6\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__15466\,
            I => \c0.data_in_0_Z0Z_6\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15461\,
            I => \N__15457\
        );

    \I__3101\ : InMux
    port map (
            O => \N__15460\,
            I => \N__15453\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__15457\,
            I => \N__15449\
        );

    \I__3099\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15446\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__15453\,
            I => \N__15443\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15440\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__15449\,
            I => \c0.d_4_6\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15446\,
            I => \c0.d_4_6\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__15443\,
            I => \c0.d_4_6\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__15440\,
            I => \c0.d_4_6\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15428\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__3090\ : Span4Mux_h
    port map (
            O => \N__15425\,
            I => \N__15420\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15424\,
            I => \N__15417\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15423\,
            I => \N__15414\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__15420\,
            I => \c0.data_in_2_Z0Z_3\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__15417\,
            I => \c0.data_in_2_Z0Z_3\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__15414\,
            I => \c0.data_in_2_Z0Z_3\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__15407\,
            I => \N__15403\
        );

    \I__3083\ : InMux
    port map (
            O => \N__15406\,
            I => \N__15398\
        );

    \I__3082\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15391\
        );

    \I__3081\ : InMux
    port map (
            O => \N__15402\,
            I => \N__15391\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15401\,
            I => \N__15391\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__15398\,
            I => \N__15387\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__15391\,
            I => \N__15384\
        );

    \I__3077\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15380\
        );

    \I__3076\ : Span4Mux_h
    port map (
            O => \N__15387\,
            I => \N__15375\
        );

    \I__3075\ : Span4Mux_v
    port map (
            O => \N__15384\,
            I => \N__15375\
        );

    \I__3074\ : InMux
    port map (
            O => \N__15383\,
            I => \N__15372\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__15380\,
            I => \c0.d_4_19\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__15375\,
            I => \c0.d_4_19\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__15372\,
            I => \c0.d_4_19\
        );

    \I__3070\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15362\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__15362\,
            I => \N__15357\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15354\
        );

    \I__3067\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15351\
        );

    \I__3066\ : Span4Mux_v
    port map (
            O => \N__15357\,
            I => \N__15345\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__15354\,
            I => \N__15345\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__15351\,
            I => \N__15342\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15339\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__15345\,
            I => \c0.d_2_31\
        );

    \I__3061\ : Odrv4
    port map (
            O => \N__15342\,
            I => \c0.d_2_31\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__15339\,
            I => \c0.d_2_31\
        );

    \I__3059\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15327\
        );

    \I__3058\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15324\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__15330\,
            I => \N__15321\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__15327\,
            I => \N__15318\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__15324\,
            I => \N__15315\
        );

    \I__3054\ : InMux
    port map (
            O => \N__15321\,
            I => \N__15312\
        );

    \I__3053\ : Span4Mux_v
    port map (
            O => \N__15318\,
            I => \N__15309\
        );

    \I__3052\ : Span4Mux_v
    port map (
            O => \N__15315\,
            I => \N__15303\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__15312\,
            I => \N__15303\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__15309\,
            I => \N__15300\
        );

    \I__3049\ : InMux
    port map (
            O => \N__15308\,
            I => \N__15297\
        );

    \I__3048\ : Span4Mux_h
    port map (
            O => \N__15303\,
            I => \N__15294\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__15300\,
            I => \c0.d_2_43\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__15297\,
            I => \c0.d_2_43\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__15294\,
            I => \c0.d_2_43\
        );

    \I__3044\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15283\
        );

    \I__3043\ : InMux
    port map (
            O => \N__15286\,
            I => \N__15279\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__15283\,
            I => \N__15276\
        );

    \I__3041\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15273\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15279\,
            I => \N__15270\
        );

    \I__3039\ : Span4Mux_h
    port map (
            O => \N__15276\,
            I => \N__15265\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__15273\,
            I => \N__15265\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__15270\,
            I => \N__15260\
        );

    \I__3036\ : Span4Mux_h
    port map (
            O => \N__15265\,
            I => \N__15260\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__15260\,
            I => \c0.d_2_15\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__15257\,
            I => \N__15254\
        );

    \I__3033\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15251\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__15251\,
            I => \N__15248\
        );

    \I__3031\ : Span4Mux_v
    port map (
            O => \N__15248\,
            I => \N__15243\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15247\,
            I => \N__15240\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__15246\,
            I => \N__15236\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__15243\,
            I => \N__15231\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__15240\,
            I => \N__15231\
        );

    \I__3026\ : InMux
    port map (
            O => \N__15239\,
            I => \N__15228\
        );

    \I__3025\ : InMux
    port map (
            O => \N__15236\,
            I => \N__15225\
        );

    \I__3024\ : Span4Mux_h
    port map (
            O => \N__15231\,
            I => \N__15222\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__15228\,
            I => \N__15217\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__15225\,
            I => \N__15217\
        );

    \I__3021\ : Span4Mux_h
    port map (
            O => \N__15222\,
            I => \N__15214\
        );

    \I__3020\ : Odrv12
    port map (
            O => \N__15217\,
            I => \c0.d_2_2\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__15214\,
            I => \c0.d_2_2\
        );

    \I__3018\ : InMux
    port map (
            O => \N__15209\,
            I => \N__15205\
        );

    \I__3017\ : CascadeMux
    port map (
            O => \N__15208\,
            I => \N__15202\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__15205\,
            I => \N__15199\
        );

    \I__3015\ : InMux
    port map (
            O => \N__15202\,
            I => \N__15196\
        );

    \I__3014\ : Span4Mux_v
    port map (
            O => \N__15199\,
            I => \N__15192\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__15196\,
            I => \N__15189\
        );

    \I__3012\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15186\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__15192\,
            I => \c0.d_2_47\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__15189\,
            I => \c0.d_2_47\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__15186\,
            I => \c0.d_2_47\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__15179\,
            I => \c0.un105_newcrc_0_a2_3_cascade_\
        );

    \I__3007\ : InMux
    port map (
            O => \N__15176\,
            I => \N__15173\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__15173\,
            I => \c0.un105_newcrc_0_a2_4\
        );

    \I__3005\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__15167\,
            I => \N__15163\
        );

    \I__3003\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15160\
        );

    \I__3002\ : Span4Mux_v
    port map (
            O => \N__15163\,
            I => \N__15154\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__15160\,
            I => \N__15154\
        );

    \I__3000\ : InMux
    port map (
            O => \N__15159\,
            I => \N__15151\
        );

    \I__2999\ : Span4Mux_h
    port map (
            O => \N__15154\,
            I => \N__15148\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__15151\,
            I => \c0.d_2_5\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__15148\,
            I => \c0.d_2_5\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15143\,
            I => \N__15139\
        );

    \I__2995\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15136\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__15139\,
            I => \N__15130\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__15136\,
            I => \N__15130\
        );

    \I__2992\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15127\
        );

    \I__2991\ : Span4Mux_v
    port map (
            O => \N__15130\,
            I => \N__15123\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__15127\,
            I => \N__15120\
        );

    \I__2989\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15117\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__15123\,
            I => \c0.d_2_32\
        );

    \I__2987\ : Odrv12
    port map (
            O => \N__15120\,
            I => \c0.d_2_32\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__15117\,
            I => \c0.d_2_32\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__15110\,
            I => \N__15107\
        );

    \I__2984\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15102\
        );

    \I__2983\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15099\
        );

    \I__2982\ : InMux
    port map (
            O => \N__15105\,
            I => \N__15095\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__15102\,
            I => \N__15092\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__15099\,
            I => \N__15089\
        );

    \I__2979\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15086\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__15095\,
            I => \N__15083\
        );

    \I__2977\ : Span4Mux_v
    port map (
            O => \N__15092\,
            I => \N__15080\
        );

    \I__2976\ : Span4Mux_v
    port map (
            O => \N__15089\,
            I => \N__15073\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__15086\,
            I => \N__15073\
        );

    \I__2974\ : Span4Mux_v
    port map (
            O => \N__15083\,
            I => \N__15073\
        );

    \I__2973\ : Span4Mux_h
    port map (
            O => \N__15080\,
            I => \N__15070\
        );

    \I__2972\ : Span4Mux_h
    port map (
            O => \N__15073\,
            I => \N__15067\
        );

    \I__2971\ : Odrv4
    port map (
            O => \N__15070\,
            I => \c0.d_2_18\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__15067\,
            I => \c0.d_2_18\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__15062\,
            I => \N__15057\
        );

    \I__2968\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15052\
        );

    \I__2967\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15049\
        );

    \I__2966\ : InMux
    port map (
            O => \N__15057\,
            I => \N__15046\
        );

    \I__2965\ : InMux
    port map (
            O => \N__15056\,
            I => \N__15041\
        );

    \I__2964\ : InMux
    port map (
            O => \N__15055\,
            I => \N__15041\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__15052\,
            I => \N__15038\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__15049\,
            I => \N__15035\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__15046\,
            I => \N__15032\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__15041\,
            I => \c0.d_2_46\
        );

    \I__2959\ : Odrv12
    port map (
            O => \N__15038\,
            I => \c0.d_2_46\
        );

    \I__2958\ : Odrv12
    port map (
            O => \N__15035\,
            I => \c0.d_2_46\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__15032\,
            I => \c0.d_2_46\
        );

    \I__2956\ : InMux
    port map (
            O => \N__15023\,
            I => \N__15018\
        );

    \I__2955\ : InMux
    port map (
            O => \N__15022\,
            I => \N__15014\
        );

    \I__2954\ : InMux
    port map (
            O => \N__15021\,
            I => \N__15011\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__15018\,
            I => \N__15008\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__15017\,
            I => \N__15005\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__15014\,
            I => \N__15002\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__15011\,
            I => \N__14999\
        );

    \I__2949\ : Span4Mux_v
    port map (
            O => \N__15008\,
            I => \N__14996\
        );

    \I__2948\ : InMux
    port map (
            O => \N__15005\,
            I => \N__14993\
        );

    \I__2947\ : Span4Mux_v
    port map (
            O => \N__15002\,
            I => \N__14990\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__14999\,
            I => \N__14987\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__14996\,
            I => \c0.d_2_20\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__14993\,
            I => \c0.d_2_20\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__14990\,
            I => \c0.d_2_20\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__14987\,
            I => \c0.d_2_20\
        );

    \I__2941\ : InMux
    port map (
            O => \N__14978\,
            I => \N__14975\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__14975\,
            I => \N__14971\
        );

    \I__2939\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14968\
        );

    \I__2938\ : Span4Mux_v
    port map (
            O => \N__14971\,
            I => \N__14965\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__14968\,
            I => \c0.nextCRC16_3_3_1\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__14965\,
            I => \c0.nextCRC16_3_3_1\
        );

    \I__2935\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14956\
        );

    \I__2934\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14953\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__14956\,
            I => \N__14950\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__14953\,
            I => \N__14947\
        );

    \I__2931\ : Span4Mux_h
    port map (
            O => \N__14950\,
            I => \N__14944\
        );

    \I__2930\ : Span4Mux_v
    port map (
            O => \N__14947\,
            I => \N__14941\
        );

    \I__2929\ : Span4Mux_v
    port map (
            O => \N__14944\,
            I => \N__14934\
        );

    \I__2928\ : Span4Mux_h
    port map (
            O => \N__14941\,
            I => \N__14934\
        );

    \I__2927\ : InMux
    port map (
            O => \N__14940\,
            I => \N__14931\
        );

    \I__2926\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14928\
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__14934\,
            I => \c0.d_2_17\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__14931\,
            I => \c0.d_2_17\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__14928\,
            I => \c0.d_2_17\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__14921\,
            I => \N__14917\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__14920\,
            I => \N__14913\
        );

    \I__2920\ : InMux
    port map (
            O => \N__14917\,
            I => \N__14909\
        );

    \I__2919\ : InMux
    port map (
            O => \N__14916\,
            I => \N__14906\
        );

    \I__2918\ : InMux
    port map (
            O => \N__14913\,
            I => \N__14903\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__14912\,
            I => \N__14900\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__14909\,
            I => \N__14896\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__14906\,
            I => \N__14893\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__14903\,
            I => \N__14890\
        );

    \I__2913\ : InMux
    port map (
            O => \N__14900\,
            I => \N__14886\
        );

    \I__2912\ : InMux
    port map (
            O => \N__14899\,
            I => \N__14883\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__14896\,
            I => \N__14880\
        );

    \I__2910\ : Span4Mux_v
    port map (
            O => \N__14893\,
            I => \N__14875\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__14890\,
            I => \N__14875\
        );

    \I__2908\ : InMux
    port map (
            O => \N__14889\,
            I => \N__14872\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14886\,
            I => \c0.d_2_1\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__14883\,
            I => \c0.d_2_1\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__14880\,
            I => \c0.d_2_1\
        );

    \I__2904\ : Odrv4
    port map (
            O => \N__14875\,
            I => \c0.d_2_1\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__14872\,
            I => \c0.d_2_1\
        );

    \I__2902\ : InMux
    port map (
            O => \N__14861\,
            I => \N__14857\
        );

    \I__2901\ : InMux
    port map (
            O => \N__14860\,
            I => \N__14853\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__14857\,
            I => \N__14850\
        );

    \I__2899\ : InMux
    port map (
            O => \N__14856\,
            I => \N__14847\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__14853\,
            I => \N__14844\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__14850\,
            I => \N__14838\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__14847\,
            I => \N__14838\
        );

    \I__2895\ : Span4Mux_h
    port map (
            O => \N__14844\,
            I => \N__14835\
        );

    \I__2894\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14832\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__14838\,
            I => \c0.d_2_4\
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__14835\,
            I => \c0.d_2_4\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__14832\,
            I => \c0.d_2_4\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__14825\,
            I => \N__14822\
        );

    \I__2889\ : InMux
    port map (
            O => \N__14822\,
            I => \N__14819\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__14819\,
            I => \c0.nextCRC16_3_0_a2_1_1\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__14816\,
            I => \N__14813\
        );

    \I__2886\ : InMux
    port map (
            O => \N__14813\,
            I => \N__14810\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__14810\,
            I => \c0.un1_data_in_6__4_0_a2_5_a2_1\
        );

    \I__2884\ : InMux
    port map (
            O => \N__14807\,
            I => \N__14804\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__14804\,
            I => \N__14800\
        );

    \I__2882\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14795\
        );

    \I__2881\ : Span4Mux_v
    port map (
            O => \N__14800\,
            I => \N__14792\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14787\
        );

    \I__2879\ : InMux
    port map (
            O => \N__14798\,
            I => \N__14787\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__14795\,
            I => \c0.N_133\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__14792\,
            I => \c0.N_133\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__14787\,
            I => \c0.N_133\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__14780\,
            I => \N__14777\
        );

    \I__2874\ : InMux
    port map (
            O => \N__14777\,
            I => \N__14774\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__14774\,
            I => \N__14771\
        );

    \I__2872\ : Span4Mux_h
    port map (
            O => \N__14771\,
            I => \N__14768\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__14768\,
            I => \c0.un1_data_in_7__2_0_a2_0_a2_5\
        );

    \I__2870\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14762\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__14759\,
            I => \c0.tx2_data_1_iv_4_6\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__2866\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14750\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__14750\,
            I => \N__14747\
        );

    \I__2864\ : Odrv4
    port map (
            O => \N__14747\,
            I => \c0.tx2_data_1_iv_3_6\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__14744\,
            I => \N__14741\
        );

    \I__2862\ : InMux
    port map (
            O => \N__14741\,
            I => \N__14738\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__14738\,
            I => \c0.tx2.r_Tx_DataZ0Z_6\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__2859\ : InMux
    port map (
            O => \N__14732\,
            I => \N__14728\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__14731\,
            I => \N__14725\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__14728\,
            I => \N__14722\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14725\,
            I => \N__14719\
        );

    \I__2855\ : Span4Mux_v
    port map (
            O => \N__14722\,
            I => \N__14714\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__14719\,
            I => \N__14714\
        );

    \I__2853\ : Span4Mux_h
    port map (
            O => \N__14714\,
            I => \N__14711\
        );

    \I__2852\ : Span4Mux_h
    port map (
            O => \N__14711\,
            I => \N__14708\
        );

    \I__2851\ : Odrv4
    port map (
            O => \N__14708\,
            I => \c0.d_2_27\
        );

    \I__2850\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14702\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__14702\,
            I => \N__14699\
        );

    \I__2848\ : Span4Mux_h
    port map (
            O => \N__14699\,
            I => \N__14696\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__14696\,
            I => \c0.tx_data_RNO_1Z0Z_3\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__14693\,
            I => \N__14690\
        );

    \I__2845\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14687\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__2843\ : Odrv12
    port map (
            O => \N__14684\,
            I => \c0.data_out_7_Z0Z_7\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__14681\,
            I => \N__14678\
        );

    \I__2841\ : InMux
    port map (
            O => \N__14678\,
            I => \N__14675\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__14675\,
            I => \N__14672\
        );

    \I__2839\ : Odrv12
    port map (
            O => \N__14672\,
            I => \c0.tx_data_RNO_1Z0Z_7\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__14669\,
            I => \c0.tx_data_RNO_3Z0Z_2_cascade_\
        );

    \I__2837\ : InMux
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__14660\,
            I => \c0.tx_data_1_0_i_ns_1_2\
        );

    \I__2834\ : InMux
    port map (
            O => \N__14657\,
            I => \N__14654\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14654\,
            I => \N__14650\
        );

    \I__2832\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14647\
        );

    \I__2831\ : Span4Mux_h
    port map (
            O => \N__14650\,
            I => \N__14642\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__14647\,
            I => \N__14642\
        );

    \I__2829\ : Span4Mux_h
    port map (
            O => \N__14642\,
            I => \N__14638\
        );

    \I__2828\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14635\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__14638\,
            I => \c0.d_2_10\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__14635\,
            I => \c0.d_2_10\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__14630\,
            I => \N__14625\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__14629\,
            I => \N__14622\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__14628\,
            I => \N__14619\
        );

    \I__2822\ : InMux
    port map (
            O => \N__14625\,
            I => \N__14615\
        );

    \I__2821\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14610\
        );

    \I__2820\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14610\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14607\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__14615\,
            I => \N__14604\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__14610\,
            I => \N__14600\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__14607\,
            I => \N__14595\
        );

    \I__2815\ : Span4Mux_v
    port map (
            O => \N__14604\,
            I => \N__14595\
        );

    \I__2814\ : InMux
    port map (
            O => \N__14603\,
            I => \N__14592\
        );

    \I__2813\ : Span4Mux_h
    port map (
            O => \N__14600\,
            I => \N__14589\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__14595\,
            I => \c0.d_2_42\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__14592\,
            I => \c0.d_2_42\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__14589\,
            I => \c0.d_2_42\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14579\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__14579\,
            I => \c0.tx_data_RNO_4Z0Z_2\
        );

    \I__2807\ : InMux
    port map (
            O => \N__14576\,
            I => \N__14573\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__14573\,
            I => \N__14570\
        );

    \I__2805\ : Span4Mux_h
    port map (
            O => \N__14570\,
            I => \N__14566\
        );

    \I__2804\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14563\
        );

    \I__2803\ : Odrv4
    port map (
            O => \N__14566\,
            I => \c0.N_81\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__14563\,
            I => \c0.N_81\
        );

    \I__2801\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14554\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14551\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__14554\,
            I => \N__14547\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__14551\,
            I => \N__14543\
        );

    \I__2797\ : InMux
    port map (
            O => \N__14550\,
            I => \N__14540\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__14547\,
            I => \N__14537\
        );

    \I__2795\ : InMux
    port map (
            O => \N__14546\,
            I => \N__14534\
        );

    \I__2794\ : Span4Mux_h
    port map (
            O => \N__14543\,
            I => \N__14529\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__14540\,
            I => \N__14529\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__14537\,
            I => \N__14526\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14534\,
            I => \c0.d_2_29\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__14529\,
            I => \c0.d_2_29\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__14526\,
            I => \c0.d_2_29\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__14519\,
            I => \N__14515\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__14518\,
            I => \N__14512\
        );

    \I__2786\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14506\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14506\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14511\,
            I => \N__14502\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14506\,
            I => \N__14497\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__14505\,
            I => \N__14494\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__14502\,
            I => \N__14491\
        );

    \I__2780\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14488\
        );

    \I__2779\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14485\
        );

    \I__2778\ : Span4Mux_h
    port map (
            O => \N__14497\,
            I => \N__14482\
        );

    \I__2777\ : InMux
    port map (
            O => \N__14494\,
            I => \N__14479\
        );

    \I__2776\ : Span4Mux_h
    port map (
            O => \N__14491\,
            I => \N__14474\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14474\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__14485\,
            I => \c0.d_2_30\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__14482\,
            I => \c0.d_2_30\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__14479\,
            I => \c0.d_2_30\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__14474\,
            I => \c0.d_2_30\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__14462\,
            I => \N__14459\
        );

    \I__2768\ : Odrv12
    port map (
            O => \N__14459\,
            I => \c0.data_out_7_Z0Z_3\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__14456\,
            I => \c0.tx2_data_1_iv_4_1_6_cascade_\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14450\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__14450\,
            I => \N__14447\
        );

    \I__2764\ : Span4Mux_h
    port map (
            O => \N__14447\,
            I => \N__14443\
        );

    \I__2763\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14440\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__14443\,
            I => \c0.data_in_5_Z0Z_3\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__14440\,
            I => \c0.data_in_5_Z0Z_3\
        );

    \I__2760\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14422\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14434\,
            I => \N__14422\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14422\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__14432\,
            I => \N__14416\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__14431\,
            I => \N__14413\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__14430\,
            I => \N__14410\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__14429\,
            I => \N__14405\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__14422\,
            I => \N__14402\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__14421\,
            I => \N__14399\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14420\,
            I => \N__14391\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14391\
        );

    \I__2749\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14391\
        );

    \I__2748\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14384\
        );

    \I__2747\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14384\
        );

    \I__2746\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14384\
        );

    \I__2745\ : InMux
    port map (
            O => \N__14408\,
            I => \N__14379\
        );

    \I__2744\ : InMux
    port map (
            O => \N__14405\,
            I => \N__14379\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__14402\,
            I => \N__14376\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14373\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14370\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__14391\,
            I => \N__14367\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__14384\,
            I => \c0.tx2.r_SM_MainZ0Z_2\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__14379\,
            I => \c0.tx2.r_SM_MainZ0Z_2\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__14376\,
            I => \c0.tx2.r_SM_MainZ0Z_2\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14373\,
            I => \c0.tx2.r_SM_MainZ0Z_2\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__14370\,
            I => \c0.tx2.r_SM_MainZ0Z_2\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__14367\,
            I => \c0.tx2.r_SM_MainZ0Z_2\
        );

    \I__2733\ : InMux
    port map (
            O => \N__14354\,
            I => \N__14351\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__14351\,
            I => \N__14344\
        );

    \I__2731\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14337\
        );

    \I__2730\ : InMux
    port map (
            O => \N__14349\,
            I => \N__14330\
        );

    \I__2729\ : InMux
    port map (
            O => \N__14348\,
            I => \N__14330\
        );

    \I__2728\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14330\
        );

    \I__2727\ : Span4Mux_h
    port map (
            O => \N__14344\,
            I => \N__14327\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14343\,
            I => \N__14322\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14342\,
            I => \N__14322\
        );

    \I__2724\ : InMux
    port map (
            O => \N__14341\,
            I => \N__14317\
        );

    \I__2723\ : InMux
    port map (
            O => \N__14340\,
            I => \N__14317\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14337\,
            I => \N__14314\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__14330\,
            I => \c0.tx2.r_SM_MainZ0Z_0\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__14327\,
            I => \c0.tx2.r_SM_MainZ0Z_0\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__14322\,
            I => \c0.tx2.r_SM_MainZ0Z_0\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__14317\,
            I => \c0.tx2.r_SM_MainZ0Z_0\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__14314\,
            I => \c0.tx2.r_SM_MainZ0Z_0\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__14303\,
            I => \c0.tx2.N_257_cascade_\
        );

    \I__2715\ : InMux
    port map (
            O => \N__14300\,
            I => \N__14297\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__14297\,
            I => \c0.tx2.N_261\
        );

    \I__2713\ : InMux
    port map (
            O => \N__14294\,
            I => \N__14288\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__14293\,
            I => \N__14284\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__14292\,
            I => \N__14281\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__14291\,
            I => \N__14278\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__14288\,
            I => \N__14275\
        );

    \I__2708\ : SRMux
    port map (
            O => \N__14287\,
            I => \N__14272\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14269\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14266\
        );

    \I__2705\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14263\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__14275\,
            I => \N__14260\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__14272\,
            I => \N__14257\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__14269\,
            I => \N__14246\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__14266\,
            I => \N__14246\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14246\
        );

    \I__2699\ : Span4Mux_h
    port map (
            O => \N__14260\,
            I => \N__14246\
        );

    \I__2698\ : Span4Mux_v
    port map (
            O => \N__14257\,
            I => \N__14246\
        );

    \I__2697\ : Span4Mux_h
    port map (
            O => \N__14246\,
            I => \N__14243\
        );

    \I__2696\ : Sp12to4
    port map (
            O => \N__14243\,
            I => \N__14240\
        );

    \I__2695\ : Odrv12
    port map (
            O => \N__14240\,
            I => \c0.tx2.o_Tx_Serial12\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__14237\,
            I => \c0.tx2.N_261_cascade_\
        );

    \I__2693\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14229\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__14233\,
            I => \N__14226\
        );

    \I__2691\ : InMux
    port map (
            O => \N__14232\,
            I => \N__14222\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__14229\,
            I => \N__14219\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14226\,
            I => \N__14214\
        );

    \I__2688\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14214\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__14222\,
            I => \c0.tx2.r_Bit_IndexZ0Z_2\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__14219\,
            I => \c0.tx2.r_Bit_IndexZ0Z_2\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__14214\,
            I => \c0.tx2.r_Bit_IndexZ0Z_2\
        );

    \I__2684\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14204\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__14204\,
            I => \N__14201\
        );

    \I__2682\ : Span4Mux_h
    port map (
            O => \N__14201\,
            I => \N__14196\
        );

    \I__2681\ : InMux
    port map (
            O => \N__14200\,
            I => \N__14191\
        );

    \I__2680\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14191\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__14196\,
            I => \c0.tx_transmitZ0\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__14191\,
            I => \c0.tx_transmitZ0\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14179\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14179\
        );

    \I__2675\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14176\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__14179\,
            I => \N__14173\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__14176\,
            I => \N__14168\
        );

    \I__2672\ : Span4Mux_h
    port map (
            O => \N__14173\,
            I => \N__14168\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__14168\,
            I => \c0.tx_active\
        );

    \I__2670\ : InMux
    port map (
            O => \N__14165\,
            I => \N__14162\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__14162\,
            I => \N__14159\
        );

    \I__2668\ : Span4Mux_h
    port map (
            O => \N__14159\,
            I => \N__14155\
        );

    \I__2667\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14152\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__14155\,
            I => \N__14147\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__14152\,
            I => \N__14144\
        );

    \I__2664\ : InMux
    port map (
            O => \N__14151\,
            I => \N__14139\
        );

    \I__2663\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14139\
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__14147\,
            I => \c0.d_4_34\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__14144\,
            I => \c0.d_4_34\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__14139\,
            I => \c0.d_4_34\
        );

    \I__2659\ : InMux
    port map (
            O => \N__14132\,
            I => \N__14129\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__14129\,
            I => \N__14126\
        );

    \I__2657\ : Span4Mux_h
    port map (
            O => \N__14126\,
            I => \N__14123\
        );

    \I__2656\ : Odrv4
    port map (
            O => \N__14123\,
            I => \c0.un1_data_in_7__7_i\
        );

    \I__2655\ : InMux
    port map (
            O => \N__14120\,
            I => \N__14117\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__14117\,
            I => \N__14114\
        );

    \I__2653\ : Odrv12
    port map (
            O => \N__14114\,
            I => \c0.tx2_data_1_0_i_1_3\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__14111\,
            I => \N__14108\
        );

    \I__2651\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14105\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__14105\,
            I => \N__14102\
        );

    \I__2649\ : Span4Mux_h
    port map (
            O => \N__14102\,
            I => \N__14099\
        );

    \I__2648\ : Span4Mux_h
    port map (
            O => \N__14099\,
            I => \N__14096\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__14096\,
            I => \c0.tx2_data_1_iv_4_1_0_3\
        );

    \I__2646\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14090\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__14090\,
            I => \N__14087\
        );

    \I__2644\ : Span4Mux_v
    port map (
            O => \N__14087\,
            I => \N__14083\
        );

    \I__2643\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14079\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__14083\,
            I => \N__14076\
        );

    \I__2641\ : InMux
    port map (
            O => \N__14082\,
            I => \N__14073\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__14079\,
            I => \c0.data_in_1_Z0Z_4\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__14076\,
            I => \c0.data_in_1_Z0Z_4\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__14073\,
            I => \c0.data_in_1_Z0Z_4\
        );

    \I__2637\ : InMux
    port map (
            O => \N__14066\,
            I => \N__14061\
        );

    \I__2636\ : InMux
    port map (
            O => \N__14065\,
            I => \N__14058\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__14064\,
            I => \N__14055\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__14061\,
            I => \N__14052\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__14058\,
            I => \N__14049\
        );

    \I__2632\ : InMux
    port map (
            O => \N__14055\,
            I => \N__14046\
        );

    \I__2631\ : Span4Mux_h
    port map (
            O => \N__14052\,
            I => \N__14043\
        );

    \I__2630\ : Span4Mux_v
    port map (
            O => \N__14049\,
            I => \N__14040\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__14046\,
            I => \N__14037\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__14043\,
            I => \c0.data_in_7_Z0Z_3\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__14040\,
            I => \c0.data_in_7_Z0Z_3\
        );

    \I__2626\ : Odrv12
    port map (
            O => \N__14037\,
            I => \c0.data_in_7_Z0Z_3\
        );

    \I__2625\ : InMux
    port map (
            O => \N__14030\,
            I => \N__14027\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__14027\,
            I => \c0.data_in_frame_7_Z0Z_3\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__14024\,
            I => \N__14019\
        );

    \I__2622\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14016\
        );

    \I__2621\ : InMux
    port map (
            O => \N__14022\,
            I => \N__14013\
        );

    \I__2620\ : InMux
    port map (
            O => \N__14019\,
            I => \N__14010\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__14016\,
            I => \N__14005\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__14013\,
            I => \N__14002\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__14010\,
            I => \N__13999\
        );

    \I__2616\ : InMux
    port map (
            O => \N__14009\,
            I => \N__13996\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__14008\,
            I => \N__13993\
        );

    \I__2614\ : Span4Mux_h
    port map (
            O => \N__14005\,
            I => \N__13990\
        );

    \I__2613\ : Span4Mux_h
    port map (
            O => \N__14002\,
            I => \N__13987\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__13999\,
            I => \N__13982\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__13996\,
            I => \N__13982\
        );

    \I__2610\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13979\
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__13990\,
            I => \c0.d_4_14\
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__13987\,
            I => \c0.d_4_14\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__13982\,
            I => \c0.d_4_14\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__13979\,
            I => \c0.d_4_14\
        );

    \I__2605\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13966\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__13969\,
            I => \N__13963\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__13966\,
            I => \N__13958\
        );

    \I__2602\ : InMux
    port map (
            O => \N__13963\,
            I => \N__13955\
        );

    \I__2601\ : InMux
    port map (
            O => \N__13962\,
            I => \N__13950\
        );

    \I__2600\ : InMux
    port map (
            O => \N__13961\,
            I => \N__13950\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__13958\,
            I => \c0.d_4_30\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__13955\,
            I => \c0.d_4_30\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__13950\,
            I => \c0.d_4_30\
        );

    \I__2596\ : InMux
    port map (
            O => \N__13943\,
            I => \N__13940\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__13940\,
            I => \N__13936\
        );

    \I__2594\ : InMux
    port map (
            O => \N__13939\,
            I => \N__13933\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__13936\,
            I => \c0.data_in_4_Z0Z_2\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__13933\,
            I => \c0.data_in_4_Z0Z_2\
        );

    \I__2591\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13924\
        );

    \I__2590\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13920\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__13924\,
            I => \N__13917\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__13923\,
            I => \N__13914\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__13920\,
            I => \N__13911\
        );

    \I__2586\ : Span4Mux_v
    port map (
            O => \N__13917\,
            I => \N__13908\
        );

    \I__2585\ : InMux
    port map (
            O => \N__13914\,
            I => \N__13905\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__13911\,
            I => \c0.data_in_1_Z0Z_3\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__13908\,
            I => \c0.data_in_1_Z0Z_3\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__13905\,
            I => \c0.data_in_1_Z0Z_3\
        );

    \I__2581\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__13892\,
            I => \N__13888\
        );

    \I__2578\ : InMux
    port map (
            O => \N__13891\,
            I => \N__13884\
        );

    \I__2577\ : Span4Mux_h
    port map (
            O => \N__13888\,
            I => \N__13881\
        );

    \I__2576\ : InMux
    port map (
            O => \N__13887\,
            I => \N__13878\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__13884\,
            I => \c0.data_in_1_Z0Z_5\
        );

    \I__2574\ : Odrv4
    port map (
            O => \N__13881\,
            I => \c0.data_in_1_Z0Z_5\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__13878\,
            I => \c0.data_in_1_Z0Z_5\
        );

    \I__2572\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__13868\,
            I => \N__13864\
        );

    \I__2570\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13860\
        );

    \I__2569\ : Span4Mux_h
    port map (
            O => \N__13864\,
            I => \N__13857\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13854\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__13860\,
            I => \c0.data_in_2_Z0Z_5\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__13857\,
            I => \c0.data_in_2_Z0Z_5\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__13854\,
            I => \c0.data_in_2_Z0Z_5\
        );

    \I__2564\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13843\
        );

    \I__2563\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13840\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__13843\,
            I => \N__13836\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__13840\,
            I => \N__13833\
        );

    \I__2560\ : InMux
    port map (
            O => \N__13839\,
            I => \N__13830\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__13836\,
            I => \c0.data_in_3_Z0Z_1\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__13833\,
            I => \c0.data_in_3_Z0Z_1\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__13830\,
            I => \c0.data_in_3_Z0Z_1\
        );

    \I__2556\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13820\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__13820\,
            I => \N__13816\
        );

    \I__2554\ : InMux
    port map (
            O => \N__13819\,
            I => \N__13813\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__13816\,
            I => \c0.data_in_5_Z0Z_1\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__13813\,
            I => \c0.data_in_5_Z0Z_1\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13808\,
            I => \N__13805\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__13805\,
            I => \N__13800\
        );

    \I__2549\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13795\
        );

    \I__2548\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13795\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__13800\,
            I => \c0.data_in_3_Z0Z_3\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__13795\,
            I => \c0.data_in_3_Z0Z_3\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__13790\,
            I => \c0.tx2_data_1_iv_3_1_6_cascade_\
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__13787\,
            I => \c0.un1_data_in_7__3_0_a2_0_a2_3_cascade_\
        );

    \I__2543\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13778\
        );

    \I__2542\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13775\
        );

    \I__2541\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13770\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13770\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__13778\,
            I => \c0.N_129\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__13775\,
            I => \c0.N_129\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__13770\,
            I => \c0.N_129\
        );

    \I__2536\ : InMux
    port map (
            O => \N__13763\,
            I => \N__13760\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__13760\,
            I => \N__13757\
        );

    \I__2534\ : Span4Mux_h
    port map (
            O => \N__13757\,
            I => \N__13752\
        );

    \I__2533\ : InMux
    port map (
            O => \N__13756\,
            I => \N__13749\
        );

    \I__2532\ : InMux
    port map (
            O => \N__13755\,
            I => \N__13746\
        );

    \I__2531\ : Odrv4
    port map (
            O => \N__13752\,
            I => \c0.data_in_2_Z0Z_1\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__13749\,
            I => \c0.data_in_2_Z0Z_1\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__13746\,
            I => \c0.data_in_2_Z0Z_1\
        );

    \I__2528\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13735\
        );

    \I__2527\ : InMux
    port map (
            O => \N__13738\,
            I => \N__13732\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13735\,
            I => \N__13726\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__13732\,
            I => \N__13726\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13731\,
            I => \N__13722\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__13726\,
            I => \N__13719\
        );

    \I__2522\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13716\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__13722\,
            I => \c0.d_4_17\
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__13719\,
            I => \c0.d_4_17\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__13716\,
            I => \c0.d_4_17\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__13706\,
            I => \N__13702\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__13705\,
            I => \N__13698\
        );

    \I__2515\ : Span4Mux_v
    port map (
            O => \N__13702\,
            I => \N__13695\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13701\,
            I => \N__13690\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13698\,
            I => \N__13690\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__13695\,
            I => \c0.data_in_3_Z0Z_6\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__13690\,
            I => \c0.data_in_3_Z0Z_6\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13682\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__13682\,
            I => \N__13679\
        );

    \I__2508\ : Span4Mux_h
    port map (
            O => \N__13679\,
            I => \N__13675\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13678\,
            I => \N__13672\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__13675\,
            I => \c0.data_in_0_Z0Z_0\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13672\,
            I => \c0.data_in_0_Z0Z_0\
        );

    \I__2504\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13664\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__13664\,
            I => \N__13661\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__13661\,
            I => \N__13656\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13660\,
            I => \N__13653\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13659\,
            I => \N__13650\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__13656\,
            I => \c0.data_in_2_Z0Z_0\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__13653\,
            I => \c0.data_in_2_Z0Z_0\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__13650\,
            I => \c0.data_in_2_Z0Z_0\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13639\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13636\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__13639\,
            I => \N__13630\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__13636\,
            I => \N__13630\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13626\
        );

    \I__2491\ : Span4Mux_v
    port map (
            O => \N__13630\,
            I => \N__13623\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13620\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__13626\,
            I => \c0.d_4_16\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__13623\,
            I => \c0.d_4_16\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__13620\,
            I => \c0.d_4_16\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__13613\,
            I => \N__13610\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13604\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13609\,
            I => \N__13604\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__13604\,
            I => \c0.d_4_0\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13601\,
            I => \N__13598\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__13598\,
            I => \N__13595\
        );

    \I__2480\ : Span4Mux_v
    port map (
            O => \N__13595\,
            I => \N__13592\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__13592\,
            I => \c0.tx2_data_RNO_3Z0Z_0\
        );

    \I__2478\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13586\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__13586\,
            I => \N__13582\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__13585\,
            I => \N__13579\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__13582\,
            I => \N__13576\
        );

    \I__2474\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13573\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__13576\,
            I => \c0.data_in_0_Z0Z_4\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__13573\,
            I => \c0.data_in_0_Z0Z_4\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__13568\,
            I => \c0.wait_for_transmission_RNOZ0Z_10_cascade_\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__13565\,
            I => \N__13562\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13559\,
            I => \N__13556\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__13556\,
            I => \N__13553\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__13553\,
            I => \c0.g0_5_4\
        );

    \I__2465\ : InMux
    port map (
            O => \N__13550\,
            I => \N__13547\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__13547\,
            I => \N__13541\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13546\,
            I => \N__13538\
        );

    \I__2462\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13535\
        );

    \I__2461\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13532\
        );

    \I__2460\ : Span4Mux_h
    port map (
            O => \N__13541\,
            I => \N__13529\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__13538\,
            I => \N__13526\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__13535\,
            I => \N__13521\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__13532\,
            I => \N__13521\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__13529\,
            I => \c0.d_4_3\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__13526\,
            I => \c0.d_4_3\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__13521\,
            I => \c0.d_4_3\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__13514\,
            I => \N__13511\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13511\,
            I => \N__13507\
        );

    \I__2451\ : InMux
    port map (
            O => \N__13510\,
            I => \N__13504\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__13507\,
            I => \N__13501\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13504\,
            I => \c0.d_4_45\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__13501\,
            I => \c0.d_4_45\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__13496\,
            I => \N__13493\
        );

    \I__2446\ : InMux
    port map (
            O => \N__13493\,
            I => \N__13490\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__13490\,
            I => \N__13487\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__13487\,
            I => \N__13484\
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__13484\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_2\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__13481\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_3_cascade_\
        );

    \I__2441\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__13475\,
            I => \c0.un1_data_in_6__7_0_a2_17_a2_5\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__13472\,
            I => \N__13469\
        );

    \I__2438\ : InMux
    port map (
            O => \N__13469\,
            I => \N__13466\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__2436\ : Span4Mux_h
    port map (
            O => \N__13463\,
            I => \N__13460\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__13460\,
            I => \N__13457\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__13457\,
            I => \c0.g3_2_1\
        );

    \I__2433\ : InMux
    port map (
            O => \N__13454\,
            I => \N__13451\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__13451\,
            I => \c0.g0_3_0\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__13448\,
            I => \c0.un1_data_in_7__0_0_a2_1_a2_3_cascade_\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__13445\,
            I => \c0.un1_data_in_7__0_0_a2_1_a2_5_0_cascade_\
        );

    \I__2429\ : InMux
    port map (
            O => \N__13442\,
            I => \N__13439\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__13439\,
            I => \c0.tx2_transmit_0_sqmuxa_1\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13433\,
            I => \N__13429\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__13432\,
            I => \N__13426\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__13429\,
            I => \N__13422\
        );

    \I__2423\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13419\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__13425\,
            I => \N__13415\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__13422\,
            I => \N__13410\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__13419\,
            I => \N__13410\
        );

    \I__2419\ : InMux
    port map (
            O => \N__13418\,
            I => \N__13405\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13415\,
            I => \N__13405\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__13410\,
            I => \N__13400\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13405\,
            I => \N__13400\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__13400\,
            I => \N__13397\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__13397\,
            I => \c0.d_2_24\
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__13394\,
            I => \N__13383\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13393\,
            I => \N__13370\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13392\,
            I => \N__13370\
        );

    \I__2410\ : InMux
    port map (
            O => \N__13391\,
            I => \N__13370\
        );

    \I__2409\ : InMux
    port map (
            O => \N__13390\,
            I => \N__13370\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13389\,
            I => \N__13370\
        );

    \I__2407\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13370\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__13387\,
            I => \N__13367\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__13386\,
            I => \N__13364\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13383\,
            I => \N__13345\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__13370\,
            I => \N__13342\
        );

    \I__2402\ : InMux
    port map (
            O => \N__13367\,
            I => \N__13331\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13364\,
            I => \N__13331\
        );

    \I__2400\ : InMux
    port map (
            O => \N__13363\,
            I => \N__13331\
        );

    \I__2399\ : InMux
    port map (
            O => \N__13362\,
            I => \N__13331\
        );

    \I__2398\ : InMux
    port map (
            O => \N__13361\,
            I => \N__13331\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13327\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13320\
        );

    \I__2395\ : InMux
    port map (
            O => \N__13358\,
            I => \N__13320\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13357\,
            I => \N__13320\
        );

    \I__2393\ : InMux
    port map (
            O => \N__13356\,
            I => \N__13315\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13315\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13354\,
            I => \N__13304\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13353\,
            I => \N__13304\
        );

    \I__2389\ : InMux
    port map (
            O => \N__13352\,
            I => \N__13304\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13351\,
            I => \N__13304\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13350\,
            I => \N__13304\
        );

    \I__2386\ : InMux
    port map (
            O => \N__13349\,
            I => \N__13295\
        );

    \I__2385\ : InMux
    port map (
            O => \N__13348\,
            I => \N__13292\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__13345\,
            I => \N__13289\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__13342\,
            I => \N__13284\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13331\,
            I => \N__13284\
        );

    \I__2381\ : InMux
    port map (
            O => \N__13330\,
            I => \N__13281\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13327\,
            I => \N__13278\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__13320\,
            I => \N__13271\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__13315\,
            I => \N__13271\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__13304\,
            I => \N__13271\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__13303\,
            I => \N__13268\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__13302\,
            I => \N__13265\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__13301\,
            I => \N__13262\
        );

    \I__2373\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13255\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13299\,
            I => \N__13255\
        );

    \I__2371\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13252\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__13295\,
            I => \N__13246\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__13292\,
            I => \N__13243\
        );

    \I__2368\ : Span4Mux_h
    port map (
            O => \N__13289\,
            I => \N__13236\
        );

    \I__2367\ : Span4Mux_h
    port map (
            O => \N__13284\,
            I => \N__13236\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__13281\,
            I => \N__13236\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__13278\,
            I => \N__13231\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__13271\,
            I => \N__13231\
        );

    \I__2363\ : InMux
    port map (
            O => \N__13268\,
            I => \N__13228\
        );

    \I__2362\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13219\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13219\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13219\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13219\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__13255\,
            I => \N__13214\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__13252\,
            I => \N__13214\
        );

    \I__2356\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13207\
        );

    \I__2355\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13207\
        );

    \I__2354\ : InMux
    port map (
            O => \N__13249\,
            I => \N__13207\
        );

    \I__2353\ : Odrv12
    port map (
            O => \N__13246\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__13243\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__13236\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__13231\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__13228\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__13219\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__13214\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__13207\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__13190\,
            I => \N__13187\
        );

    \I__2344\ : InMux
    port map (
            O => \N__13187\,
            I => \N__13183\
        );

    \I__2343\ : InMux
    port map (
            O => \N__13186\,
            I => \N__13180\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__13183\,
            I => \N__13176\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__13180\,
            I => \N__13173\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13170\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__13176\,
            I => \c0.N_105\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__13173\,
            I => \c0.N_105\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__13170\,
            I => \c0.N_105\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13163\,
            I => \N__13160\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__13160\,
            I => \N__13156\
        );

    \I__2334\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13153\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__13156\,
            I => \c0.nextCRC16_3_2_1\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__13153\,
            I => \c0.nextCRC16_3_2_1\
        );

    \I__2331\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13144\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13140\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13144\,
            I => \N__13137\
        );

    \I__2328\ : InMux
    port map (
            O => \N__13143\,
            I => \N__13134\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__13140\,
            I => \c0.N_106\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__13137\,
            I => \c0.N_106\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__13134\,
            I => \c0.N_106\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__13127\,
            I => \N__13124\
        );

    \I__2323\ : InMux
    port map (
            O => \N__13124\,
            I => \N__13121\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13121\,
            I => \N__13118\
        );

    \I__2321\ : Span4Mux_h
    port map (
            O => \N__13118\,
            I => \N__13115\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__13115\,
            I => \c0.data_out_7_Z0Z_1\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__13112\,
            I => \N__13109\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13106\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13106\,
            I => \c0.data_in_frame_7_Z0Z_5\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__13103\,
            I => \N__13100\
        );

    \I__2315\ : InMux
    port map (
            O => \N__13100\,
            I => \N__13097\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__13097\,
            I => \c0.data_in_frame_7_Z0Z_7\
        );

    \I__2313\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13087\
        );

    \I__2312\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13087\
        );

    \I__2311\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13084\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__13087\,
            I => \N__13081\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__13084\,
            I => \N__13078\
        );

    \I__2308\ : Span4Mux_v
    port map (
            O => \N__13081\,
            I => \N__13075\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__13078\,
            I => \c0.d_2_28\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__13075\,
            I => \c0.d_2_28\
        );

    \I__2305\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13067\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__13067\,
            I => \c0.nextCRC16_3_0_a2_1_2\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__13064\,
            I => \N__13061\
        );

    \I__2302\ : InMux
    port map (
            O => \N__13061\,
            I => \N__13056\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13060\,
            I => \N__13051\
        );

    \I__2300\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13051\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__13056\,
            I => \c0.d_2_0\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__13051\,
            I => \c0.d_2_0\
        );

    \I__2297\ : InMux
    port map (
            O => \N__13046\,
            I => \N__13043\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__13043\,
            I => \N__13040\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__13040\,
            I => \c0.nextCRC16_3_4_0\
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__13037\,
            I => \N__13034\
        );

    \I__2293\ : InMux
    port map (
            O => \N__13034\,
            I => \N__13031\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__13031\,
            I => \N__13026\
        );

    \I__2291\ : InMux
    port map (
            O => \N__13030\,
            I => \N__13021\
        );

    \I__2290\ : InMux
    port map (
            O => \N__13029\,
            I => \N__13021\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__13026\,
            I => \c0.d_2_13\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__13021\,
            I => \c0.d_2_13\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13016\,
            I => \N__13013\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__13013\,
            I => \N__13008\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13012\,
            I => \N__13005\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__13011\,
            I => \N__13000\
        );

    \I__2283\ : Span4Mux_v
    port map (
            O => \N__13008\,
            I => \N__12995\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__13005\,
            I => \N__12995\
        );

    \I__2281\ : InMux
    port map (
            O => \N__13004\,
            I => \N__12992\
        );

    \I__2280\ : InMux
    port map (
            O => \N__13003\,
            I => \N__12989\
        );

    \I__2279\ : InMux
    port map (
            O => \N__13000\,
            I => \N__12986\
        );

    \I__2278\ : Sp12to4
    port map (
            O => \N__12995\,
            I => \N__12981\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__12992\,
            I => \N__12981\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__12989\,
            I => \c0.d_2_26\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__12986\,
            I => \c0.d_2_26\
        );

    \I__2274\ : Odrv12
    port map (
            O => \N__12981\,
            I => \c0.d_2_26\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__12974\,
            I => \c0.nextCRC16_3_4_0_cascade_\
        );

    \I__2272\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12968\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__12968\,
            I => \N__12964\
        );

    \I__2270\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12961\
        );

    \I__2269\ : Span12Mux_s7_v
    port map (
            O => \N__12964\,
            I => \N__12957\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__12961\,
            I => \N__12954\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12960\,
            I => \N__12951\
        );

    \I__2266\ : Odrv12
    port map (
            O => \N__12957\,
            I => \c0.N_99\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__12954\,
            I => \c0.N_99\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__12951\,
            I => \c0.N_99\
        );

    \I__2263\ : InMux
    port map (
            O => \N__12944\,
            I => \N__12941\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__12941\,
            I => \c0.nextCRC16_3_0_a2_3_0\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__12938\,
            I => \N__12935\
        );

    \I__2260\ : InMux
    port map (
            O => \N__12935\,
            I => \N__12929\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12934\,
            I => \N__12926\
        );

    \I__2258\ : InMux
    port map (
            O => \N__12933\,
            I => \N__12923\
        );

    \I__2257\ : InMux
    port map (
            O => \N__12932\,
            I => \N__12920\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__12929\,
            I => \N__12916\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__12926\,
            I => \N__12913\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__12923\,
            I => \N__12910\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__12920\,
            I => \N__12907\
        );

    \I__2252\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12904\
        );

    \I__2251\ : Span4Mux_h
    port map (
            O => \N__12916\,
            I => \N__12901\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__12913\,
            I => \N__12896\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__12910\,
            I => \N__12896\
        );

    \I__2248\ : Odrv12
    port map (
            O => \N__12907\,
            I => \c0.d_2_39\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12904\,
            I => \c0.d_2_39\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__12901\,
            I => \c0.d_2_39\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__12896\,
            I => \c0.d_2_39\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__12887\,
            I => \N__12884\
        );

    \I__2243\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12881\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__12881\,
            I => \N__12878\
        );

    \I__2241\ : Span4Mux_h
    port map (
            O => \N__12878\,
            I => \N__12875\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__12875\,
            I => \c0.data_out_6_Z0Z_5\
        );

    \I__2239\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12869\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__12869\,
            I => \c0.nextCRC16_3_0_a2_4_15\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__12866\,
            I => \N__12863\
        );

    \I__2236\ : InMux
    port map (
            O => \N__12863\,
            I => \N__12860\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__12860\,
            I => \N__12857\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__12857\,
            I => \N__12854\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__12854\,
            I => \c0.nextCRC16_3_0_a2_3_15\
        );

    \I__2232\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12848\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__12848\,
            I => \N__12845\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__12845\,
            I => \N__12842\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__12842\,
            I => \c0.data_out_6_Z0Z_7\
        );

    \I__2228\ : InMux
    port map (
            O => \N__12839\,
            I => \N__12835\
        );

    \I__2227\ : InMux
    port map (
            O => \N__12838\,
            I => \N__12832\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__12835\,
            I => \N__12829\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__12832\,
            I => \N__12825\
        );

    \I__2224\ : Span4Mux_h
    port map (
            O => \N__12829\,
            I => \N__12822\
        );

    \I__2223\ : InMux
    port map (
            O => \N__12828\,
            I => \N__12817\
        );

    \I__2222\ : Span4Mux_v
    port map (
            O => \N__12825\,
            I => \N__12814\
        );

    \I__2221\ : Span4Mux_h
    port map (
            O => \N__12822\,
            I => \N__12811\
        );

    \I__2220\ : InMux
    port map (
            O => \N__12821\,
            I => \N__12806\
        );

    \I__2219\ : InMux
    port map (
            O => \N__12820\,
            I => \N__12806\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__12817\,
            I => \N__12803\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__12814\,
            I => \c0.d_2_16\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__12811\,
            I => \c0.d_2_16\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__12806\,
            I => \c0.d_2_16\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__12803\,
            I => \c0.d_2_16\
        );

    \I__2213\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12791\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__12791\,
            I => \N__12787\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12790\,
            I => \N__12783\
        );

    \I__2210\ : Span4Mux_h
    port map (
            O => \N__12787\,
            I => \N__12780\
        );

    \I__2209\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12777\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__12783\,
            I => \c0.d_2_9\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__12780\,
            I => \c0.d_2_9\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__12777\,
            I => \c0.d_2_9\
        );

    \I__2205\ : InMux
    port map (
            O => \N__12770\,
            I => \N__12766\
        );

    \I__2204\ : InMux
    port map (
            O => \N__12769\,
            I => \N__12763\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__12766\,
            I => \N__12760\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__12763\,
            I => \N__12757\
        );

    \I__2201\ : Span4Mux_h
    port map (
            O => \N__12760\,
            I => \N__12754\
        );

    \I__2200\ : Span4Mux_h
    port map (
            O => \N__12757\,
            I => \N__12751\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__12754\,
            I => \c0.N_94\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__12751\,
            I => \c0.N_94\
        );

    \I__2197\ : InMux
    port map (
            O => \N__12746\,
            I => \N__12743\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__12743\,
            I => \N__12740\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__12740\,
            I => \N__12737\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__12737\,
            I => \N__12734\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__12734\,
            I => \c0.tx_data_RNO_4Z0Z_5\
        );

    \I__2192\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12727\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12730\,
            I => \N__12724\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__12727\,
            I => \N__12721\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__12724\,
            I => \N__12718\
        );

    \I__2188\ : Span4Mux_h
    port map (
            O => \N__12721\,
            I => \N__12715\
        );

    \I__2187\ : Span4Mux_h
    port map (
            O => \N__12718\,
            I => \N__12712\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__12715\,
            I => \c0.d_2_45\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__12712\,
            I => \c0.d_2_45\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12707\,
            I => \N__12704\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__12704\,
            I => \c0.nextCRC16_3_0_a2_0_0\
        );

    \I__2182\ : InMux
    port map (
            O => \N__12701\,
            I => \N__12698\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__12698\,
            I => \c0.nextCRC16_3_0_a2_4_0\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12692\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__12692\,
            I => \N__12689\
        );

    \I__2178\ : Span4Mux_h
    port map (
            O => \N__12689\,
            I => \N__12686\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__12686\,
            I => \c0.tx2.r_Tx_DataZ0Z_3\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__12683\,
            I => \c0.tx2.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12680\,
            I => \N__12677\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__12677\,
            I => \c0.tx2.N_349\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__12674\,
            I => \c0.tx2.N_346_cascade_\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__12671\,
            I => \c0.tx2.N_279_cascade_\
        );

    \I__2171\ : IoInMux
    port map (
            O => \N__12668\,
            I => \N__12665\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12665\,
            I => \N__12661\
        );

    \I__2169\ : InMux
    port map (
            O => \N__12664\,
            I => \N__12658\
        );

    \I__2168\ : Span12Mux_s11_h
    port map (
            O => \N__12661\,
            I => \N__12655\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__12658\,
            I => \N__12652\
        );

    \I__2166\ : Odrv12
    port map (
            O => \N__12655\,
            I => \PIN_3_c\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__12652\,
            I => \PIN_3_c\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12647\,
            I => \N__12644\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__12644\,
            I => \N__12641\
        );

    \I__2162\ : Span12Mux_v
    port map (
            O => \N__12641\,
            I => \N__12638\
        );

    \I__2161\ : Odrv12
    port map (
            O => \N__12638\,
            I => \c0.tx2.r_Tx_Active_1_sqmuxa\
        );

    \I__2160\ : InMux
    port map (
            O => \N__12635\,
            I => \N__12632\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__12632\,
            I => \N__12629\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__12629\,
            I => \c0.tx_data_RNO_3Z0Z_1\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__12626\,
            I => \c0.tx2.m5_0_0_cascade_\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12623\,
            I => \N__12620\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__12620\,
            I => \N__12617\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__12617\,
            I => \N__12614\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__12614\,
            I => \c0.tx2_data_RNO_0Z0Z_0\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__12611\,
            I => \c0.tx2_data_1_0_i_ns_1_0_cascade_\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__12608\,
            I => \N__12605\
        );

    \I__2150\ : InMux
    port map (
            O => \N__12605\,
            I => \N__12602\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__12602\,
            I => \N__12595\
        );

    \I__2148\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12592\
        );

    \I__2147\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12587\
        );

    \I__2146\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12587\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12598\,
            I => \N__12584\
        );

    \I__2144\ : Odrv12
    port map (
            O => \N__12595\,
            I => \c0.d_4_1\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__12592\,
            I => \c0.d_4_1\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__12587\,
            I => \c0.d_4_1\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__12584\,
            I => \c0.d_4_1\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__12575\,
            I => \c0.tx2_data_RNO_3Z0Z_1_cascade_\
        );

    \I__2139\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12569\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__12569\,
            I => \N__12566\
        );

    \I__2137\ : Span4Mux_v
    port map (
            O => \N__12566\,
            I => \N__12563\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__12563\,
            I => \c0.tx2_data_RNO_1Z0Z_1\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__12560\,
            I => \c0.tx2_data_1_0_i_ns_1_1_cascade_\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12557\,
            I => \N__12554\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__12554\,
            I => \N__12551\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__12551\,
            I => \N__12548\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__12548\,
            I => \c0.tx2_data_RNO_0Z0Z_1\
        );

    \I__2130\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12542\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__12542\,
            I => \c0.tx2_data_RNO_4Z0Z_1\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12536\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__12536\,
            I => \c0.tx2_data_RNO_1Z0Z_0\
        );

    \I__2126\ : InMux
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__12530\,
            I => \N__12527\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__12527\,
            I => \N__12524\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__12524\,
            I => \c0.tx2.r_Tx_DataZ0Z_2\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12518\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__12518\,
            I => \c0.tx2.r_Tx_DataZ0Z_0\
        );

    \I__2120\ : InMux
    port map (
            O => \N__12515\,
            I => \N__12512\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__12512\,
            I => \c0.tx2.r_Tx_Data_pmux_3_i_m2_ns_1\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12506\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__12506\,
            I => \c0.tx2.r_Tx_DataZ0Z_1\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__12503\,
            I => \c0.un1_data_in_7__1_0_a2_24_a2_2_cascade_\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12497\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12497\,
            I => \N__12493\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__12496\,
            I => \N__12488\
        );

    \I__2112\ : Span4Mux_h
    port map (
            O => \N__12493\,
            I => \N__12484\
        );

    \I__2111\ : InMux
    port map (
            O => \N__12492\,
            I => \N__12481\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12491\,
            I => \N__12474\
        );

    \I__2109\ : InMux
    port map (
            O => \N__12488\,
            I => \N__12474\
        );

    \I__2108\ : InMux
    port map (
            O => \N__12487\,
            I => \N__12474\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__12484\,
            I => \c0.d_4_2\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__12481\,
            I => \c0.d_4_2\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__12474\,
            I => \c0.d_4_2\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12464\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__12464\,
            I => \N__12460\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12457\
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__12460\,
            I => \c0.N_103\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__12457\,
            I => \c0.N_103\
        );

    \I__2099\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12449\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__12449\,
            I => \c0.wait_for_transmission4_13_1_1\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__12446\,
            I => \c0.un1_data_in_7__1_0_a2_24_a2_6_cascade_\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__12443\,
            I => \c0.un1_data_in_7__1_0_a2_24_a2_1_cascade_\
        );

    \I__2095\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12437\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__12437\,
            I => \c0.un1_data_in_7__1_0_a2_24_a2_5\
        );

    \I__2093\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12431\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__12431\,
            I => \N__12428\
        );

    \I__2091\ : Odrv4
    port map (
            O => \N__12428\,
            I => \c0.d_4_RNITCRCZ0Z_29\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__12425\,
            I => \c0.tx2_data_RNO_4Z0Z_0_cascade_\
        );

    \I__2089\ : InMux
    port map (
            O => \N__12422\,
            I => \N__12419\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__12419\,
            I => \N__12416\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__12416\,
            I => \c0.un1_data_in_7__4_0_a2_0_a2_4\
        );

    \I__2086\ : InMux
    port map (
            O => \N__12413\,
            I => \N__12410\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__12410\,
            I => \N__12406\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__12409\,
            I => \N__12403\
        );

    \I__2083\ : Span4Mux_h
    port map (
            O => \N__12406\,
            I => \N__12400\
        );

    \I__2082\ : InMux
    port map (
            O => \N__12403\,
            I => \N__12397\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__12400\,
            I => \c0.data_in_0_Z0Z_2\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__12397\,
            I => \c0.data_in_0_Z0Z_2\
        );

    \I__2079\ : InMux
    port map (
            O => \N__12392\,
            I => \N__12389\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__12389\,
            I => \c0.d_4_RNID6K21_0Z0Z_15\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12386\,
            I => \N__12383\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__12383\,
            I => \c0.d_4_RNID6K21Z0Z_15\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12380\,
            I => \N__12377\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__12377\,
            I => \N__12374\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__12374\,
            I => \N__12370\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12373\,
            I => \N__12367\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__12370\,
            I => \c0.data_in_0_Z0Z_1\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__12367\,
            I => \c0.data_in_0_Z0Z_1\
        );

    \I__2069\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12357\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__12361\,
            I => \N__12354\
        );

    \I__2067\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12351\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__12357\,
            I => \N__12348\
        );

    \I__2065\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12345\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__12351\,
            I => \N__12340\
        );

    \I__2063\ : Span4Mux_h
    port map (
            O => \N__12348\,
            I => \N__12340\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__12345\,
            I => \N__12337\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__12340\,
            I => \c0.data_in_1_Z0Z_7\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__12337\,
            I => \c0.data_in_1_Z0Z_7\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12332\,
            I => \N__12328\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12325\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__12328\,
            I => \N__12321\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__12325\,
            I => \N__12318\
        );

    \I__2055\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12315\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__12321\,
            I => \c0.data_in_3_Z0Z_7\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__12318\,
            I => \c0.data_in_3_Z0Z_7\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__12315\,
            I => \c0.data_in_3_Z0Z_7\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__12308\,
            I => \c0.un1_data_in_6__0_0_a2_5_a2_2_cascade_\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__12305\,
            I => \c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__12302\,
            I => \c0.un1_data_in_7__4_i_cascade_\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12299\,
            I => \N__12296\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__12296\,
            I => \c0.un1_data_in_6__0\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__12293\,
            I => \c0.d_4_RNIF73E2Z0Z_14_cascade_\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__12290\,
            I => \c0.d_4_RNIMKFE3Z0Z_14_cascade_\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__12287\,
            I => \c0.un1_data_in_6__7_cascade_\
        );

    \I__2043\ : InMux
    port map (
            O => \N__12284\,
            I => \N__12281\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__12281\,
            I => \c0.wait_for_transmission4_12\
        );

    \I__2041\ : IoInMux
    port map (
            O => \N__12278\,
            I => \N__12275\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__12275\,
            I => \N__12272\
        );

    \I__2039\ : IoSpan4Mux
    port map (
            O => \N__12272\,
            I => \N__12269\
        );

    \I__2038\ : Span4Mux_s2_h
    port map (
            O => \N__12269\,
            I => \N__12266\
        );

    \I__2037\ : Sp12to4
    port map (
            O => \N__12266\,
            I => \N__12262\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12259\
        );

    \I__2035\ : Span12Mux_s10_h
    port map (
            O => \N__12262\,
            I => \N__12256\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__12259\,
            I => \c0.data_in_frame_0__0_sqmuxa\
        );

    \I__2033\ : Odrv12
    port map (
            O => \N__12256\,
            I => \c0.data_in_frame_0__0_sqmuxa\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__12251\,
            I => \c0.wait_for_transmission4_12_cascade_\
        );

    \I__2031\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12245\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__12245\,
            I => \N__12241\
        );

    \I__2029\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12238\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__12241\,
            I => \c0.dataZ0Z_15\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__12238\,
            I => \c0.dataZ0Z_15\
        );

    \I__2026\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12226\
        );

    \I__2025\ : InMux
    port map (
            O => \N__12232\,
            I => \N__12226\
        );

    \I__2024\ : InMux
    port map (
            O => \N__12231\,
            I => \N__12223\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12226\,
            I => \N__12220\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__12223\,
            I => \c0.tx2_active\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__12220\,
            I => \c0.tx2_active\
        );

    \I__2020\ : InMux
    port map (
            O => \N__12215\,
            I => \N__12212\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__12212\,
            I => \c0.tx2_data_1_iv_5_1_0_7\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__12209\,
            I => \c0.tx2_data_1_iv_5_1_7_cascade_\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12203\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__12203\,
            I => \c0.data_in_frame_6_Z0Z_7\
        );

    \I__2015\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12197\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__12197\,
            I => \N__12194\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__12194\,
            I => \N__12191\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__12191\,
            I => \c0.tx2_data_1_iv_3_1_3\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__12188\,
            I => \N__12185\
        );

    \I__2010\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12182\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__12182\,
            I => \N__12179\
        );

    \I__2008\ : Span4Mux_v
    port map (
            O => \N__12179\,
            I => \N__12176\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__12176\,
            I => \c0.tx2_data_1_iv_3_3\
        );

    \I__2006\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12170\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__12170\,
            I => \N__12167\
        );

    \I__2004\ : Span4Mux_h
    port map (
            O => \N__12167\,
            I => \N__12163\
        );

    \I__2003\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12160\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__12163\,
            I => \c0.data_in_0_Z0Z_3\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__12160\,
            I => \c0.data_in_0_Z0Z_3\
        );

    \I__2000\ : InMux
    port map (
            O => \N__12155\,
            I => \N__12152\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__12152\,
            I => \c0.N_247_0\
        );

    \I__1998\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12145\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__12148\,
            I => \N__12141\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__12145\,
            I => \N__12138\
        );

    \I__1995\ : InMux
    port map (
            O => \N__12144\,
            I => \N__12133\
        );

    \I__1994\ : InMux
    port map (
            O => \N__12141\,
            I => \N__12133\
        );

    \I__1993\ : Span4Mux_h
    port map (
            O => \N__12138\,
            I => \N__12130\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__12133\,
            I => \c0.d_2_41\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__12130\,
            I => \c0.d_2_41\
        );

    \I__1990\ : InMux
    port map (
            O => \N__12125\,
            I => \N__12118\
        );

    \I__1989\ : InMux
    port map (
            O => \N__12124\,
            I => \N__12118\
        );

    \I__1988\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12115\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__12118\,
            I => \c0.d_2_12\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__12115\,
            I => \c0.d_2_12\
        );

    \I__1985\ : InMux
    port map (
            O => \N__12110\,
            I => \N__12107\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__12107\,
            I => \N__12102\
        );

    \I__1983\ : InMux
    port map (
            O => \N__12106\,
            I => \N__12099\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__12105\,
            I => \N__12094\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__12102\,
            I => \N__12089\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__12099\,
            I => \N__12089\
        );

    \I__1979\ : InMux
    port map (
            O => \N__12098\,
            I => \N__12086\
        );

    \I__1978\ : InMux
    port map (
            O => \N__12097\,
            I => \N__12083\
        );

    \I__1977\ : InMux
    port map (
            O => \N__12094\,
            I => \N__12080\
        );

    \I__1976\ : Odrv4
    port map (
            O => \N__12089\,
            I => \c0.d_2_40\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__12086\,
            I => \c0.d_2_40\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__12083\,
            I => \c0.d_2_40\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__12080\,
            I => \c0.d_2_40\
        );

    \I__1972\ : InMux
    port map (
            O => \N__12071\,
            I => \N__12068\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__12068\,
            I => \c0.nextCRC16_3_0_a2_2_2\
        );

    \I__1970\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12061\
        );

    \I__1969\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12058\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__12061\,
            I => \N__12055\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__12058\,
            I => \N__12052\
        );

    \I__1966\ : Span4Mux_h
    port map (
            O => \N__12055\,
            I => \N__12049\
        );

    \I__1965\ : Span4Mux_v
    port map (
            O => \N__12052\,
            I => \N__12046\
        );

    \I__1964\ : Span4Mux_h
    port map (
            O => \N__12049\,
            I => \N__12043\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__12046\,
            I => \c0.d_2_3\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__12043\,
            I => \c0.d_2_3\
        );

    \I__1961\ : InMux
    port map (
            O => \N__12038\,
            I => \N__12035\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__12035\,
            I => \N__12031\
        );

    \I__1959\ : InMux
    port map (
            O => \N__12034\,
            I => \N__12028\
        );

    \I__1958\ : Odrv12
    port map (
            O => \N__12031\,
            I => \c0.N_75\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__12028\,
            I => \c0.N_75\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__12023\,
            I => \c0.N_75_cascade_\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__12020\,
            I => \N__12017\
        );

    \I__1954\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12014\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__12014\,
            I => \N__12010\
        );

    \I__1952\ : InMux
    port map (
            O => \N__12013\,
            I => \N__12007\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__12010\,
            I => \c0.d_2_44\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__12007\,
            I => \c0.d_2_44\
        );

    \I__1949\ : InMux
    port map (
            O => \N__12002\,
            I => \N__11999\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__11999\,
            I => \c0.N_95\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__11996\,
            I => \N__11992\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__11995\,
            I => \N__11988\
        );

    \I__1945\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11985\
        );

    \I__1944\ : InMux
    port map (
            O => \N__11991\,
            I => \N__11982\
        );

    \I__1943\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11979\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__11985\,
            I => \N__11974\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__11982\,
            I => \N__11974\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__11979\,
            I => \N__11971\
        );

    \I__1939\ : Span4Mux_h
    port map (
            O => \N__11974\,
            I => \N__11968\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__11971\,
            I => \N__11965\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__11968\,
            I => \c0.d_2_14\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__11965\,
            I => \c0.d_2_14\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__11960\,
            I => \c0.N_95_cascade_\
        );

    \I__1934\ : InMux
    port map (
            O => \N__11957\,
            I => \N__11951\
        );

    \I__1933\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11948\
        );

    \I__1932\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11945\
        );

    \I__1931\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11942\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__11951\,
            I => \N__11939\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__11948\,
            I => \N__11936\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__11945\,
            I => \N__11933\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__11942\,
            I => \N__11930\
        );

    \I__1926\ : Span4Mux_h
    port map (
            O => \N__11939\,
            I => \N__11927\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__11936\,
            I => \N__11924\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__11933\,
            I => \N__11919\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__11930\,
            I => \N__11919\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__11927\,
            I => \c0.d_2_25\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__11924\,
            I => \c0.d_2_25\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__11919\,
            I => \c0.d_2_25\
        );

    \I__1919\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11908\
        );

    \I__1918\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11904\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__11908\,
            I => \N__11900\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11907\,
            I => \N__11897\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__11904\,
            I => \N__11894\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__11903\,
            I => \N__11891\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__11900\,
            I => \N__11888\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__11897\,
            I => \N__11883\
        );

    \I__1911\ : Span12Mux_s6_v
    port map (
            O => \N__11894\,
            I => \N__11883\
        );

    \I__1910\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11880\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__11888\,
            I => \c0.d_2_11\
        );

    \I__1908\ : Odrv12
    port map (
            O => \N__11883\,
            I => \c0.d_2_11\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11880\,
            I => \c0.d_2_11\
        );

    \I__1906\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11870\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__11870\,
            I => \N__11866\
        );

    \I__1904\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11863\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__11866\,
            I => \c0.dataZ0Z_8\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__11863\,
            I => \c0.dataZ0Z_8\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__11858\,
            I => \N__11855\
        );

    \I__1900\ : InMux
    port map (
            O => \N__11855\,
            I => \N__11852\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__11852\,
            I => \c0.nextCRC16_3_0_a2_1_8\
        );

    \I__1898\ : InMux
    port map (
            O => \N__11849\,
            I => \N__11845\
        );

    \I__1897\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11842\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__11845\,
            I => \N__11837\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__11842\,
            I => \N__11837\
        );

    \I__1894\ : Span4Mux_h
    port map (
            O => \N__11837\,
            I => \N__11834\
        );

    \I__1893\ : Span4Mux_h
    port map (
            O => \N__11834\,
            I => \N__11830\
        );

    \I__1892\ : InMux
    port map (
            O => \N__11833\,
            I => \N__11827\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__11830\,
            I => \c0.N_77\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__11827\,
            I => \c0.N_77\
        );

    \I__1889\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11819\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__11819\,
            I => \c0.data_out_6_Z0Z_0\
        );

    \I__1887\ : InMux
    port map (
            O => \N__11816\,
            I => \N__11813\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__11813\,
            I => \N__11810\
        );

    \I__1885\ : Span4Mux_h
    port map (
            O => \N__11810\,
            I => \N__11806\
        );

    \I__1884\ : InMux
    port map (
            O => \N__11809\,
            I => \N__11803\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__11806\,
            I => \c0.dataZ0Z_0\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__11803\,
            I => \c0.dataZ0Z_0\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11798\,
            I => \N__11795\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__11795\,
            I => \c0.data_out_7_Z0Z_0\
        );

    \I__1879\ : InMux
    port map (
            O => \N__11792\,
            I => \N__11789\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__11789\,
            I => \N__11785\
        );

    \I__1877\ : InMux
    port map (
            O => \N__11788\,
            I => \N__11782\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__11785\,
            I => \c0.d_2_8\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__11782\,
            I => \c0.d_2_8\
        );

    \I__1874\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__11774\,
            I => \N__11771\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__11771\,
            I => \c0.tx_data_RNO_0Z0Z_0\
        );

    \I__1871\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11765\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__11765\,
            I => \c0.N_93\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__11762\,
            I => \N__11759\
        );

    \I__1868\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__11753\,
            I => \c0.nextCRC16_3_0_a2_0_10\
        );

    \I__1865\ : InMux
    port map (
            O => \N__11750\,
            I => \N__11743\
        );

    \I__1864\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11743\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__11748\,
            I => \N__11740\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__11743\,
            I => \N__11736\
        );

    \I__1861\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11731\
        );

    \I__1860\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11731\
        );

    \I__1859\ : Span4Mux_h
    port map (
            O => \N__11736\,
            I => \N__11728\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__11731\,
            I => \c0.d_2_22\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__11728\,
            I => \c0.d_2_22\
        );

    \I__1856\ : InMux
    port map (
            O => \N__11723\,
            I => \N__11720\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__11717\,
            I => \N__11713\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11710\
        );

    \I__1852\ : Span4Mux_h
    port map (
            O => \N__11713\,
            I => \N__11704\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__11710\,
            I => \N__11704\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11709\,
            I => \N__11700\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__11704\,
            I => \N__11697\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11694\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__11700\,
            I => \c0.d_2_6\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__11697\,
            I => \c0.d_2_6\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11694\,
            I => \c0.d_2_6\
        );

    \I__1844\ : InMux
    port map (
            O => \N__11687\,
            I => \N__11684\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__11684\,
            I => \N__11681\
        );

    \I__1842\ : Odrv12
    port map (
            O => \N__11681\,
            I => \c0.nextCRC16_3_9\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__11678\,
            I => \c0.nextCRC16_3_0_a2_6_0_15_cascade_\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11675\,
            I => \N__11672\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__11672\,
            I => \N__11668\
        );

    \I__1838\ : InMux
    port map (
            O => \N__11671\,
            I => \N__11665\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__11668\,
            I => \N__11660\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__11665\,
            I => \N__11660\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__11660\,
            I => \c0.N_92\
        );

    \I__1834\ : InMux
    port map (
            O => \N__11657\,
            I => \c0.tx2.r_Clock_Count12\
        );

    \I__1833\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11650\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__11653\,
            I => \N__11646\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__11650\,
            I => \N__11643\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11640\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11637\
        );

    \I__1828\ : Span4Mux_h
    port map (
            O => \N__11643\,
            I => \N__11634\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__11640\,
            I => \N__11631\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__11637\,
            I => \c0.N_76\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__11634\,
            I => \c0.N_76\
        );

    \I__1824\ : Odrv12
    port map (
            O => \N__11631\,
            I => \c0.N_76\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__11624\,
            I => \N__11621\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11618\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__11618\,
            I => \c0.data_out_6_Z0Z_2\
        );

    \I__1820\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11612\,
            I => \c0.tx_data_RNO_0Z0Z_2\
        );

    \I__1818\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__11606\,
            I => \N__11601\
        );

    \I__1816\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11598\
        );

    \I__1815\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11595\
        );

    \I__1814\ : Span4Mux_v
    port map (
            O => \N__11601\,
            I => \N__11588\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__11598\,
            I => \N__11588\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__11595\,
            I => \N__11588\
        );

    \I__1811\ : Span4Mux_h
    port map (
            O => \N__11588\,
            I => \N__11584\
        );

    \I__1810\ : InMux
    port map (
            O => \N__11587\,
            I => \N__11581\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__11584\,
            I => \c0.d_2_21\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__11581\,
            I => \c0.d_2_21\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__11576\,
            I => \c0.tx_data_1_iv_i_m2_0_ns_1_0_cascade_\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__11573\,
            I => \c0.N_304_cascade_\
        );

    \I__1805\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11567\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__11567\,
            I => \N__11564\
        );

    \I__1803\ : Span4Mux_h
    port map (
            O => \N__11564\,
            I => \N__11561\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__11561\,
            I => \c0.tx_data_1_iv_i_1_0\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11558\,
            I => \c0.tx2.un1_r_Clock_Count_cry_2\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11555\,
            I => \N__11552\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__11552\,
            I => \c0.tx2.r_Clock_Count_RNO_0_0_3\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__11549\,
            I => \N__11545\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11542\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11539\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__11542\,
            I => \c0.tx2.r_Clock_Count_0_sqmuxa\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__11539\,
            I => \c0.tx2.r_Clock_Count_0_sqmuxa\
        );

    \I__1793\ : InMux
    port map (
            O => \N__11534\,
            I => \N__11531\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__11531\,
            I => \c0.tx2.r_Clock_Count_RNO_0_0_0\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11524\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11527\,
            I => \N__11521\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__11524\,
            I => \c0.tx2.r_Clock_CountZ0Z_0\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__11521\,
            I => \c0.tx2.r_Clock_CountZ0Z_0\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11516\,
            I => \N__11513\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__11513\,
            I => \c0.tx2.r_Clock_Count_RNO_0_0_1\
        );

    \I__1785\ : InMux
    port map (
            O => \N__11510\,
            I => \N__11506\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11509\,
            I => \N__11503\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__11506\,
            I => \c0.tx2.r_Clock_Count_i_0\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11503\,
            I => \c0.tx2.r_Clock_Count_i_0\
        );

    \I__1781\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11494\
        );

    \I__1780\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11491\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__11494\,
            I => \c0.tx2.r_Clock_CountZ0Z_1\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__11491\,
            I => \c0.tx2.r_Clock_CountZ0Z_1\
        );

    \I__1777\ : InMux
    port map (
            O => \N__11486\,
            I => \N__11483\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__11483\,
            I => \c0.tx2.r_Clock_Count_i_1\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11476\
        );

    \I__1774\ : InMux
    port map (
            O => \N__11479\,
            I => \N__11473\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__11476\,
            I => \c0.tx2.r_Clock_CountZ0Z_2\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__11473\,
            I => \c0.tx2.r_Clock_CountZ0Z_2\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11465\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__11465\,
            I => \c0.tx2.r_Clock_Count_i_2\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11462\,
            I => \N__11458\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11461\,
            I => \N__11455\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11458\,
            I => \c0.tx2.r_Clock_CountZ0Z_3\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__11455\,
            I => \c0.tx2.r_Clock_CountZ0Z_3\
        );

    \I__1765\ : InMux
    port map (
            O => \N__11450\,
            I => \N__11447\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__11447\,
            I => \c0.tx2.r_Clock_Count_i_3\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11440\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11437\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__11440\,
            I => \N__11433\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__11437\,
            I => \N__11430\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11427\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__11433\,
            I => \c0.data_in_3_Z0Z_4\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__11430\,
            I => \c0.data_in_3_Z0Z_4\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__11427\,
            I => \c0.data_in_3_Z0Z_4\
        );

    \I__1755\ : InMux
    port map (
            O => \N__11420\,
            I => \N__11415\
        );

    \I__1754\ : InMux
    port map (
            O => \N__11419\,
            I => \N__11412\
        );

    \I__1753\ : InMux
    port map (
            O => \N__11418\,
            I => \N__11409\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__11415\,
            I => \N__11406\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__11412\,
            I => \N__11403\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__11409\,
            I => \c0.data_in_1_Z0Z_6\
        );

    \I__1749\ : Odrv12
    port map (
            O => \N__11406\,
            I => \c0.data_in_1_Z0Z_6\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__11403\,
            I => \c0.data_in_1_Z0Z_6\
        );

    \I__1747\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11392\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11389\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__11392\,
            I => \N__11385\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__11389\,
            I => \N__11382\
        );

    \I__1743\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11379\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__11385\,
            I => \c0.data_in_3_Z0Z_5\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__11382\,
            I => \c0.data_in_3_Z0Z_5\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__11379\,
            I => \c0.data_in_3_Z0Z_5\
        );

    \I__1739\ : InMux
    port map (
            O => \N__11372\,
            I => \N__11368\
        );

    \I__1738\ : InMux
    port map (
            O => \N__11371\,
            I => \N__11365\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__11368\,
            I => \c0.data_in_5_Z0Z_2\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11365\,
            I => \c0.data_in_5_Z0Z_2\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11360\,
            I => \c0.tx2.un1_r_Clock_Count_cry_0\
        );

    \I__1734\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11354\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__11354\,
            I => \c0.tx2.r_Clock_Count_RNO_0_0_2\
        );

    \I__1732\ : InMux
    port map (
            O => \N__11351\,
            I => \c0.tx2.un1_r_Clock_Count_cry_1\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__11348\,
            I => \c0.g3_2_0_cascade_\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11342\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__11342\,
            I => \c0.g0_2\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__11336\,
            I => \N__11333\
        );

    \I__1726\ : Span4Mux_h
    port map (
            O => \N__11333\,
            I => \N__11329\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11326\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__11329\,
            I => \c0.rx_data_1\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__11326\,
            I => \c0.rx_data_1\
        );

    \I__1722\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11317\
        );

    \I__1721\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11314\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__11317\,
            I => \c0.data_in_4_Z0Z_0\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__11314\,
            I => \c0.data_in_4_Z0Z_0\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__11309\,
            I => \c0.g1_cascade_\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11306\,
            I => \N__11303\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__11303\,
            I => \c0.g0_3\
        );

    \I__1715\ : InMux
    port map (
            O => \N__11300\,
            I => \N__11297\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__11297\,
            I => \c0.byte_transmit_counter2_0_sqmuxa_0\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__11294\,
            I => \c0.g1_1_cascade_\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11291\,
            I => \N__11288\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__11288\,
            I => \c0.N_72_mux\
        );

    \I__1710\ : CascadeMux
    port map (
            O => \N__11285\,
            I => \c0.N_249_cascade_\
        );

    \I__1709\ : InMux
    port map (
            O => \N__11282\,
            I => \N__11278\
        );

    \I__1708\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11275\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__11278\,
            I => \c0.dataZ0Z_5\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__11275\,
            I => \c0.dataZ0Z_5\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11270\,
            I => \N__11266\
        );

    \I__1704\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11263\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__11266\,
            I => \c0.dataZ0Z_13\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11263\,
            I => \c0.dataZ0Z_13\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11258\,
            I => \N__11253\
        );

    \I__1700\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11250\
        );

    \I__1699\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11246\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__11253\,
            I => \N__11241\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__11250\,
            I => \N__11241\
        );

    \I__1696\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11238\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__11246\,
            I => \N__11235\
        );

    \I__1694\ : Span4Mux_h
    port map (
            O => \N__11241\,
            I => \N__11232\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__11238\,
            I => \N__11229\
        );

    \I__1692\ : Odrv12
    port map (
            O => \N__11235\,
            I => \c0.d_2_37\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__11232\,
            I => \c0.d_2_37\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__11229\,
            I => \c0.d_2_37\
        );

    \I__1689\ : InMux
    port map (
            O => \N__11222\,
            I => \N__11218\
        );

    \I__1688\ : InMux
    port map (
            O => \N__11221\,
            I => \N__11215\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__11218\,
            I => \c0.dataZ0Z_4\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__11215\,
            I => \c0.dataZ0Z_4\
        );

    \I__1685\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11206\
        );

    \I__1684\ : InMux
    port map (
            O => \N__11209\,
            I => \N__11203\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__11206\,
            I => \c0.dataZ0Z_9\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__11203\,
            I => \c0.dataZ0Z_9\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__1680\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11192\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__11192\,
            I => \c0.i12_7_and\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__11189\,
            I => \c0.tx_data_RNO_3Z0Z_4_cascade_\
        );

    \I__1677\ : InMux
    port map (
            O => \N__11186\,
            I => \N__11183\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__11183\,
            I => \N__11180\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__11180\,
            I => \c0.tx_data_1_0_i_ns_1_4\
        );

    \I__1674\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11174\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__11174\,
            I => \c0.tx_data_RNO_4Z0Z_4\
        );

    \I__1672\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11168\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__11168\,
            I => \N__11165\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__11165\,
            I => \c0.data_out_7_Z0Z_4\
        );

    \I__1669\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11158\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11155\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__11158\,
            I => \c0.dataZ0Z_7\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__11155\,
            I => \c0.dataZ0Z_7\
        );

    \I__1665\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11146\
        );

    \I__1664\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11143\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__11146\,
            I => \c0.dataZ0Z_3\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__11143\,
            I => \c0.dataZ0Z_3\
        );

    \I__1661\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11134\
        );

    \I__1660\ : InMux
    port map (
            O => \N__11137\,
            I => \N__11131\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__11134\,
            I => \c0.dataZ0Z_10\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__11131\,
            I => \c0.dataZ0Z_10\
        );

    \I__1657\ : InMux
    port map (
            O => \N__11126\,
            I => \N__11122\
        );

    \I__1656\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11119\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__11122\,
            I => \c0.dataZ0Z_6\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__11119\,
            I => \c0.dataZ0Z_6\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11114\,
            I => \N__11110\
        );

    \I__1652\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11107\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__11110\,
            I => \c0.dataZ0Z_2\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__11107\,
            I => \c0.dataZ0Z_2\
        );

    \I__1649\ : InMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__1647\ : Span4Mux_v
    port map (
            O => \N__11096\,
            I => \N__11093\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__11093\,
            I => \c0.data_out_7_Z0Z_2\
        );

    \I__1645\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__1643\ : Span4Mux_h
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__11081\,
            I => \c0.tx_data_RNO_0Z0Z_5\
        );

    \I__1641\ : InMux
    port map (
            O => \N__11078\,
            I => \N__11071\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11077\,
            I => \N__11071\
        );

    \I__1639\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11068\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__11071\,
            I => \N__11065\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__11068\,
            I => \N__11059\
        );

    \I__1636\ : Span4Mux_h
    port map (
            O => \N__11065\,
            I => \N__11059\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__11064\,
            I => \N__11056\
        );

    \I__1634\ : Span4Mux_h
    port map (
            O => \N__11059\,
            I => \N__11053\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11050\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__11053\,
            I => \c0.d_2_23\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__11050\,
            I => \c0.d_2_23\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11042\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__11042\,
            I => \c0.tx_data_RNO_0Z0Z_7\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__11039\,
            I => \N__11036\
        );

    \I__1627\ : InMux
    port map (
            O => \N__11036\,
            I => \N__11033\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__11033\,
            I => \N__11030\
        );

    \I__1625\ : Span4Mux_h
    port map (
            O => \N__11030\,
            I => \N__11027\
        );

    \I__1624\ : Span4Mux_h
    port map (
            O => \N__11027\,
            I => \N__11024\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__11024\,
            I => \c0.tx_data_RNO_1Z0Z_1\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__11021\,
            I => \N__11018\
        );

    \I__1621\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11015\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__11015\,
            I => \c0.tx_data_RNO_1Z0Z_2\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__11012\,
            I => \c0.nextCRC16_3_0_a2_1_15_cascade_\
        );

    \I__1618\ : InMux
    port map (
            O => \N__11009\,
            I => \N__11006\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__11006\,
            I => \N__11003\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__11003\,
            I => \c0.m115_amcf1\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__11000\,
            I => \c0.N_293_cascade_\
        );

    \I__1614\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10994\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__10994\,
            I => \N__10991\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__10991\,
            I => \c0.tx_data_1_0_i_1_6\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__10988\,
            I => \c0.tx_data_RNO_1Z0Z_6_cascade_\
        );

    \I__1610\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10982\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__10982\,
            I => \N__10979\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__10979\,
            I => \N__10976\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__10976\,
            I => \c0.tx.r_Tx_DataZ0Z_6\
        );

    \I__1606\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10970\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__10970\,
            I => \N__10967\
        );

    \I__1604\ : Span4Mux_h
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__10964\,
            I => \c0.tx.r_Tx_DataZ0Z_2\
        );

    \I__1602\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10958\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__10958\,
            I => \c0.tx_data_1_0_i_ns_1_7\
        );

    \I__1600\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10952\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__10952\,
            I => \N__10949\
        );

    \I__1598\ : Span4Mux_h
    port map (
            O => \N__10949\,
            I => \N__10946\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__10946\,
            I => \c0.tx.r_Tx_DataZ0Z_7\
        );

    \I__1596\ : CEMux
    port map (
            O => \N__10943\,
            I => \N__10937\
        );

    \I__1595\ : CEMux
    port map (
            O => \N__10942\,
            I => \N__10934\
        );

    \I__1594\ : CEMux
    port map (
            O => \N__10941\,
            I => \N__10931\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__10940\,
            I => \N__10928\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__10937\,
            I => \N__10925\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__10934\,
            I => \N__10922\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__10931\,
            I => \N__10918\
        );

    \I__1589\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10915\
        );

    \I__1588\ : Span4Mux_h
    port map (
            O => \N__10925\,
            I => \N__10912\
        );

    \I__1587\ : Span4Mux_h
    port map (
            O => \N__10922\,
            I => \N__10909\
        );

    \I__1586\ : InMux
    port map (
            O => \N__10921\,
            I => \N__10906\
        );

    \I__1585\ : Span4Mux_v
    port map (
            O => \N__10918\,
            I => \N__10901\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__10915\,
            I => \N__10901\
        );

    \I__1583\ : Span4Mux_h
    port map (
            O => \N__10912\,
            I => \N__10898\
        );

    \I__1582\ : Span4Mux_h
    port map (
            O => \N__10909\,
            I => \N__10895\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__10906\,
            I => \N__10892\
        );

    \I__1580\ : Span4Mux_h
    port map (
            O => \N__10901\,
            I => \N__10889\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__10898\,
            I => \c0.tx.r_Tx_Data_0_sqmuxa\
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__10895\,
            I => \c0.tx.r_Tx_Data_0_sqmuxa\
        );

    \I__1577\ : Odrv12
    port map (
            O => \N__10892\,
            I => \c0.tx.r_Tx_Data_0_sqmuxa\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__10889\,
            I => \c0.tx.r_Tx_Data_0_sqmuxa\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__10880\,
            I => \N__10877\
        );

    \I__1574\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10874\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__10874\,
            I => \N__10871\
        );

    \I__1572\ : Span4Mux_h
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__10868\,
            I => \c0.tx_data_RNO_1Z0Z_4\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__1569\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10859\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__10859\,
            I => \N__10856\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__10853\,
            I => \c0.data_out_6_Z0Z_1\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__10850\,
            I => \N__10846\
        );

    \I__1564\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10843\
        );

    \I__1563\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10840\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__10843\,
            I => \N__10837\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__10840\,
            I => \N__10834\
        );

    \I__1560\ : Odrv12
    port map (
            O => \N__10837\,
            I => \c0.rx.un1_r_Rx_Byte_7\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__10834\,
            I => \c0.rx.un1_r_Rx_Byte_7\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__10829\,
            I => \c0.tx2.o_Tx_Serial12_cascade_\
        );

    \I__1557\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10823\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__1555\ : Span4Mux_h
    port map (
            O => \N__10820\,
            I => \N__10817\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__10817\,
            I => \c0.tx_data_RNO_3Z0Z_3\
        );

    \I__1553\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10808\
        );

    \I__1552\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10805\
        );

    \I__1551\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10802\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10799\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__10808\,
            I => \N__10796\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__10805\,
            I => \c0.d_2_38\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__10802\,
            I => \c0.d_2_38\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__10799\,
            I => \c0.d_2_38\
        );

    \I__1545\ : Odrv4
    port map (
            O => \N__10796\,
            I => \c0.d_2_38\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__10784\,
            I => \N__10780\
        );

    \I__1542\ : InMux
    port map (
            O => \N__10783\,
            I => \N__10777\
        );

    \I__1541\ : Odrv12
    port map (
            O => \N__10780\,
            I => \c0.rx_data_5\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__10777\,
            I => \c0.rx_data_5\
        );

    \I__1539\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10769\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__10769\,
            I => \c0.tx2_data_RNO_4Z0Z_2\
        );

    \I__1537\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__10763\,
            I => \c0.tx2_data_RNO_1Z0Z_2\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__10760\,
            I => \c0.tx2_data_RNO_0Z0Z_2_cascade_\
        );

    \I__1534\ : InMux
    port map (
            O => \N__10757\,
            I => \N__10754\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__10754\,
            I => \c0.tx2_data_1_0_i_ns_1_2\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10751\,
            I => \N__10748\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__10745\,
            I => \c0.tx2_data_1_iv_4_3\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10736\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__10736\,
            I => \c0.i12_4_and\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__10733\,
            I => \N__10730\
        );

    \I__1525\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10727\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__1523\ : Odrv4
    port map (
            O => \N__10724\,
            I => \c0.i12_6_and\
        );

    \I__1522\ : CascadeMux
    port map (
            O => \N__10721\,
            I => \N__10718\
        );

    \I__1521\ : InMux
    port map (
            O => \N__10718\,
            I => \N__10715\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__10715\,
            I => \c0.i12_5_and\
        );

    \I__1519\ : InMux
    port map (
            O => \N__10712\,
            I => \bfn_10_18_0_\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__10709\,
            I => \N__10706\
        );

    \I__1517\ : InMux
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__10703\,
            I => \c0.i12_1_and\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__1514\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10694\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__10694\,
            I => \c0.i12_3_and\
        );

    \I__1512\ : InMux
    port map (
            O => \N__10691\,
            I => \c0.data_cry_13\
        );

    \I__1511\ : InMux
    port map (
            O => \N__10688\,
            I => \c0.data_cry_14\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__1509\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10679\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__10679\,
            I => \c0.i12_0_and\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10670\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__10670\,
            I => \c0.i12_2_and\
        );

    \I__1504\ : InMux
    port map (
            O => \N__10667\,
            I => \c0.data_cry_5\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10664\,
            I => \c0.data_cry_6\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10661\,
            I => \bfn_9_28_0_\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10658\,
            I => \c0.data_cry_8\
        );

    \I__1500\ : InMux
    port map (
            O => \N__10655\,
            I => \c0.data_cry_9\
        );

    \I__1499\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10649\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__1497\ : Span4Mux_h
    port map (
            O => \N__10646\,
            I => \N__10642\
        );

    \I__1496\ : InMux
    port map (
            O => \N__10645\,
            I => \N__10639\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__10642\,
            I => \c0.dataZ0Z_11\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__10639\,
            I => \c0.dataZ0Z_11\
        );

    \I__1493\ : InMux
    port map (
            O => \N__10634\,
            I => \c0.data_cry_10\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10628\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10628\,
            I => \N__10624\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10621\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__10624\,
            I => \c0.dataZ0Z_12\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__10621\,
            I => \c0.dataZ0Z_12\
        );

    \I__1487\ : InMux
    port map (
            O => \N__10616\,
            I => \c0.data_cry_11\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10613\,
            I => \c0.data_cry_12\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10607\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__10607\,
            I => \N__10603\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10606\,
            I => \N__10600\
        );

    \I__1482\ : Odrv12
    port map (
            O => \N__10603\,
            I => \c0.dataZ0Z_14\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__10600\,
            I => \c0.dataZ0Z_14\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__10595\,
            I => \c0.N_74_cascade_\
        );

    \I__1479\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10588\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10585\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__10588\,
            I => \c0.d_2_19\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10585\,
            I => \c0.d_2_19\
        );

    \I__1475\ : InMux
    port map (
            O => \N__10580\,
            I => \bfn_9_27_0_\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10574\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__10574\,
            I => \N__10570\
        );

    \I__1472\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10567\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__10570\,
            I => \c0.dataZ0Z_1\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__10567\,
            I => \c0.dataZ0Z_1\
        );

    \I__1469\ : InMux
    port map (
            O => \N__10562\,
            I => \c0.data_cry_0\
        );

    \I__1468\ : InMux
    port map (
            O => \N__10559\,
            I => \c0.data_cry_1\
        );

    \I__1467\ : InMux
    port map (
            O => \N__10556\,
            I => \c0.data_cry_2\
        );

    \I__1466\ : InMux
    port map (
            O => \N__10553\,
            I => \c0.data_cry_3\
        );

    \I__1465\ : InMux
    port map (
            O => \N__10550\,
            I => \c0.data_cry_4\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__10547\,
            I => \c0.tx_data_RNO_4Z0Z_1_cascade_\
        );

    \I__1463\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__10541\,
            I => \N__10538\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__10538\,
            I => \c0.tx_data_1_0_i_ns_1_1\
        );

    \I__1460\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10532\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__10532\,
            I => \N__10529\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__10529\,
            I => \N__10526\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__10526\,
            I => \c0.tx_data_RNO_0Z0Z_3\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__10523\,
            I => \c0.nextCRC16_3_0_a2_1_11_cascade_\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__10520\,
            I => \N__10517\
        );

    \I__1454\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10514\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__10514\,
            I => \c0.data_out_6_Z0Z_3\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10511\,
            I => \N__10507\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10504\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__10507\,
            I => \N__10501\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__10504\,
            I => \N__10498\
        );

    \I__1448\ : Odrv12
    port map (
            O => \N__10501\,
            I => \c0.d_2_7\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__10498\,
            I => \c0.d_2_7\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__10493\,
            I => \c0.tx_data_RNO_3Z0Z_7_cascade_\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10487\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__10487\,
            I => \c0.tx_data_RNO_4Z0Z_7\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10481\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__1441\ : Span4Mux_h
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__10475\,
            I => \c0.N_74\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10465\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10462\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10459\
        );

    \I__1436\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10454\
        );

    \I__1435\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10454\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__10465\,
            I => \N__10450\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10445\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__10459\,
            I => \N__10445\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__10454\,
            I => \N__10442\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10453\,
            I => \N__10436\
        );

    \I__1429\ : Span4Mux_v
    port map (
            O => \N__10450\,
            I => \N__10431\
        );

    \I__1428\ : Span4Mux_v
    port map (
            O => \N__10445\,
            I => \N__10431\
        );

    \I__1427\ : Span4Mux_v
    port map (
            O => \N__10442\,
            I => \N__10428\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10441\,
            I => \N__10423\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10423\
        );

    \I__1424\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10420\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__10436\,
            I => \c0.tx.r_SM_MainZ0Z_0\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__10431\,
            I => \c0.tx.r_SM_MainZ0Z_0\
        );

    \I__1421\ : Odrv4
    port map (
            O => \N__10428\,
            I => \c0.tx.r_SM_MainZ0Z_0\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10423\,
            I => \c0.tx.r_SM_MainZ0Z_0\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__10420\,
            I => \c0.tx.r_SM_MainZ0Z_0\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__10409\,
            I => \N__10404\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__10408\,
            I => \N__10399\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10394\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10391\
        );

    \I__1414\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10388\
        );

    \I__1413\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10385\
        );

    \I__1412\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10382\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10379\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10375\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__10394\,
            I => \N__10370\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__10391\,
            I => \N__10370\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__10388\,
            I => \N__10363\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10363\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__10382\,
            I => \N__10358\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__10379\,
            I => \N__10358\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10355\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__10375\,
            I => \N__10350\
        );

    \I__1401\ : Span4Mux_v
    port map (
            O => \N__10370\,
            I => \N__10350\
        );

    \I__1400\ : InMux
    port map (
            O => \N__10369\,
            I => \N__10345\
        );

    \I__1399\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10345\
        );

    \I__1398\ : Span4Mux_h
    port map (
            O => \N__10363\,
            I => \N__10342\
        );

    \I__1397\ : Span4Mux_h
    port map (
            O => \N__10358\,
            I => \N__10339\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__10355\,
            I => \c0.tx.r_SM_MainZ0Z_1\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__10350\,
            I => \c0.tx.r_SM_MainZ0Z_1\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__10345\,
            I => \c0.tx.r_SM_MainZ0Z_1\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__10342\,
            I => \c0.tx.r_SM_MainZ0Z_1\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__10339\,
            I => \c0.tx.r_SM_MainZ0Z_1\
        );

    \I__1391\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10324\
        );

    \I__1390\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10321\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__10324\,
            I => \N__10313\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__10321\,
            I => \N__10313\
        );

    \I__1387\ : InMux
    port map (
            O => \N__10320\,
            I => \N__10310\
        );

    \I__1386\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10307\
        );

    \I__1385\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10297\
        );

    \I__1384\ : Span4Mux_h
    port map (
            O => \N__10313\,
            I => \N__10294\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__10310\,
            I => \N__10289\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__10307\,
            I => \N__10289\
        );

    \I__1381\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10282\
        );

    \I__1380\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10282\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10282\
        );

    \I__1378\ : InMux
    port map (
            O => \N__10303\,
            I => \N__10273\
        );

    \I__1377\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10273\
        );

    \I__1376\ : InMux
    port map (
            O => \N__10301\,
            I => \N__10273\
        );

    \I__1375\ : InMux
    port map (
            O => \N__10300\,
            I => \N__10273\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__10297\,
            I => \c0.tx.r_Clock_Count12_THRU_CO\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__10294\,
            I => \c0.tx.r_Clock_Count12_THRU_CO\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__10289\,
            I => \c0.tx.r_Clock_Count12_THRU_CO\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__10282\,
            I => \c0.tx.r_Clock_Count12_THRU_CO\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__10273\,
            I => \c0.tx.r_Clock_Count12_THRU_CO\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__10262\,
            I => \N__10256\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10261\,
            I => \N__10250\
        );

    \I__1367\ : InMux
    port map (
            O => \N__10260\,
            I => \N__10247\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__10259\,
            I => \N__10241\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10256\,
            I => \N__10236\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__10255\,
            I => \N__10233\
        );

    \I__1363\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10228\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10228\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__10250\,
            I => \N__10225\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__10247\,
            I => \N__10222\
        );

    \I__1359\ : InMux
    port map (
            O => \N__10246\,
            I => \N__10213\
        );

    \I__1358\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10213\
        );

    \I__1357\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10213\
        );

    \I__1356\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10213\
        );

    \I__1355\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10210\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__10239\,
            I => \N__10206\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__10236\,
            I => \N__10203\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10200\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__10228\,
            I => \N__10197\
        );

    \I__1350\ : Span4Mux_h
    port map (
            O => \N__10225\,
            I => \N__10190\
        );

    \I__1349\ : Span4Mux_v
    port map (
            O => \N__10222\,
            I => \N__10190\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__10213\,
            I => \N__10190\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__10210\,
            I => \N__10187\
        );

    \I__1346\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10182\
        );

    \I__1345\ : InMux
    port map (
            O => \N__10206\,
            I => \N__10182\
        );

    \I__1344\ : Span4Mux_v
    port map (
            O => \N__10203\,
            I => \N__10175\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__10200\,
            I => \N__10175\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__10197\,
            I => \N__10175\
        );

    \I__1341\ : Span4Mux_h
    port map (
            O => \N__10190\,
            I => \N__10172\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__10187\,
            I => \c0.tx.r_SM_MainZ0Z_2\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__10182\,
            I => \c0.tx.r_SM_MainZ0Z_2\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__10175\,
            I => \c0.tx.r_SM_MainZ0Z_2\
        );

    \I__1337\ : Odrv4
    port map (
            O => \N__10172\,
            I => \c0.tx.r_SM_MainZ0Z_2\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__10163\,
            I => \c0.nextCRC16_3_3_12_cascade_\
        );

    \I__1335\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__10157\,
            I => \c0.nextCRC16_3_4_12\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10151\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__10148\,
            I => \c0.data_out_6_Z0Z_4\
        );

    \I__1330\ : InMux
    port map (
            O => \N__10145\,
            I => \N__10142\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__10142\,
            I => \N__10139\
        );

    \I__1328\ : Span4Mux_v
    port map (
            O => \N__10139\,
            I => \N__10136\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__10136\,
            I => \c0.tx_data_RNO_0Z0Z_4\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__10133\,
            I => \c0.rx.r_Rx_Bytece_0_3_cascade_\
        );

    \I__1325\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10126\
        );

    \I__1324\ : InMux
    port map (
            O => \N__10129\,
            I => \N__10123\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__10126\,
            I => \c0.rx_data_3\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__10123\,
            I => \c0.rx_data_3\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__10118\,
            I => \c0.tx2_data_RNO_3Z0Z_2_cascade_\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__10115\,
            I => \c0.tx_data_RNO_1Z0Z_0_cascade_\
        );

    \I__1319\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__1317\ : Odrv4
    port map (
            O => \N__10106\,
            I => \c0.tx.r_Tx_DataZ0Z_0\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__1315\ : InMux
    port map (
            O => \N__10100\,
            I => \N__10097\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__10097\,
            I => \c0.tx.r_Tx_DataZ0Z_4\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10091\,
            I => \N__10088\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__1310\ : Span4Mux_h
    port map (
            O => \N__10085\,
            I => \N__10082\
        );

    \I__1309\ : Odrv4
    port map (
            O => \N__10082\,
            I => \c0.data_out_7_Z0Z_5\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__10079\,
            I => \c0.tx_data_1_0_i_ns_1_3_cascade_\
        );

    \I__1307\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__10073\,
            I => \c0.tx.r_Tx_DataZ0Z_3\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__10070\,
            I => \N__10067\
        );

    \I__1304\ : InMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__10064\,
            I => \c0.tx_data_RNO_1Z0Z_5\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__10061\,
            I => \N__10058\
        );

    \I__1301\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10055\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__10055\,
            I => \c0.tx.r_Tx_DataZ0Z_5\
        );

    \I__1299\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10049\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__10049\,
            I => \c0.tx_data_RNO_4Z0Z_3\
        );

    \I__1297\ : InMux
    port map (
            O => \N__10046\,
            I => \N__10040\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10045\,
            I => \N__10037\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10044\,
            I => \N__10034\
        );

    \I__1294\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10031\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__10040\,
            I => \c0.tx.r_Bit_IndexZ0Z_2\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__10037\,
            I => \c0.tx.r_Bit_IndexZ0Z_2\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__10034\,
            I => \c0.tx.r_Bit_IndexZ0Z_2\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__10031\,
            I => \c0.tx.r_Bit_IndexZ0Z_2\
        );

    \I__1289\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10012\
        );

    \I__1288\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10012\
        );

    \I__1287\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10007\
        );

    \I__1286\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10007\
        );

    \I__1285\ : InMux
    port map (
            O => \N__10018\,
            I => \N__10002\
        );

    \I__1284\ : InMux
    port map (
            O => \N__10017\,
            I => \N__10002\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__10012\,
            I => \c0.tx.r_Bit_IndexZ0Z_1\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__10007\,
            I => \c0.tx.r_Bit_IndexZ0Z_1\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__10002\,
            I => \c0.tx.r_Bit_IndexZ0Z_1\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__9995\,
            I => \c0.tx.r_Tx_Data_pmux_3_i_m2_ns_1_cascade_\
        );

    \I__1279\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__9989\,
            I => \c0.tx.N_354\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__9986\,
            I => \N__9982\
        );

    \I__1276\ : InMux
    port map (
            O => \N__9985\,
            I => \N__9977\
        );

    \I__1275\ : InMux
    port map (
            O => \N__9982\,
            I => \N__9974\
        );

    \I__1274\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9969\
        );

    \I__1273\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9969\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__9977\,
            I => \N__9966\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__9974\,
            I => \c0.tx.r_Bit_IndexZ0Z_0\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__9969\,
            I => \c0.tx.r_Bit_IndexZ0Z_0\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__9966\,
            I => \c0.tx.r_Bit_IndexZ0Z_0\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__9959\,
            I => \c0.tx.N_357_cascade_\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__1265\ : Odrv12
    port map (
            O => \N__9950\,
            I => \c0.tx.N_320\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__9947\,
            I => \c0.tx_data_RNO_3Z0Z_5_cascade_\
        );

    \I__1263\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__9941\,
            I => \c0.tx_data_1_0_i_ns_1_5\
        );

    \I__1261\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9934\
        );

    \I__1260\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9931\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__9934\,
            I => \N__9928\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__9931\,
            I => \N__9925\
        );

    \I__1257\ : Span4Mux_h
    port map (
            O => \N__9928\,
            I => \N__9919\
        );

    \I__1256\ : Span4Mux_v
    port map (
            O => \N__9925\,
            I => \N__9919\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9916\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__9919\,
            I => \c0.rx.r_Rx_DV6\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__9916\,
            I => \c0.rx.r_Rx_DV6\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__9911\,
            I => \c0.tx.r_Tx_Active_1_sqmuxa_cascade_\
        );

    \I__1251\ : InMux
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__9905\,
            I => \c0.tx_data_RNO_0Z0Z_1\
        );

    \I__1249\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__9899\,
            I => \c0.tx.r_Tx_DataZ0Z_1\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__9896\,
            I => \c0.tx.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__9893\,
            I => \c0.rx.r_Rx_Bytece_1_1_cascade_\
        );

    \I__1245\ : InMux
    port map (
            O => \N__9890\,
            I => \N__9887\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__9887\,
            I => \c0.rx.r_Rx_Bytece_1_5\
        );

    \I__1243\ : InMux
    port map (
            O => \N__9884\,
            I => \N__9880\
        );

    \I__1242\ : InMux
    port map (
            O => \N__9883\,
            I => \N__9877\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__9880\,
            I => \c0.tx.r_Clock_Count_i_0\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__9877\,
            I => \c0.tx.r_Clock_Count_i_0\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9868\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9865\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__9868\,
            I => \c0.tx.r_Clock_CountZ0Z_1\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__9865\,
            I => \c0.tx.r_Clock_CountZ0Z_1\
        );

    \I__1235\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__9857\,
            I => \c0.tx.r_Clock_Count_i_1\
        );

    \I__1233\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9850\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9853\,
            I => \N__9847\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__9850\,
            I => \c0.tx.r_Clock_CountZ0Z_2\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__9847\,
            I => \c0.tx.r_Clock_CountZ0Z_2\
        );

    \I__1229\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9839\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__9839\,
            I => \c0.tx.r_Clock_Count_i_2\
        );

    \I__1227\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9832\
        );

    \I__1226\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9829\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__9832\,
            I => \c0.tx.r_Clock_CountZ0Z_3\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__9829\,
            I => \c0.tx.r_Clock_CountZ0Z_3\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9821\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__9821\,
            I => \c0.tx.r_Clock_Count_i_3\
        );

    \I__1221\ : InMux
    port map (
            O => \N__9818\,
            I => \c0.tx.r_Clock_Count12\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9815\,
            I => blink_counter_cry_24
        );

    \I__1219\ : InMux
    port map (
            O => \N__9812\,
            I => \N__9808\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9811\,
            I => \N__9805\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__9808\,
            I => \N__9800\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__9805\,
            I => \N__9800\
        );

    \I__1215\ : Span4Mux_v
    port map (
            O => \N__9800\,
            I => \N__9796\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9799\,
            I => \N__9793\
        );

    \I__1213\ : Odrv4
    port map (
            O => \N__9796\,
            I => \blink_counterZ0Z_25\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__9793\,
            I => \blink_counterZ0Z_25\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__9788\,
            I => \c0.tx.N_287_cascade_\
        );

    \I__1210\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9782\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__9782\,
            I => \c0.tx.N_294\
        );

    \I__1208\ : SRMux
    port map (
            O => \N__9779\,
            I => \N__9774\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__9778\,
            I => \N__9770\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__9777\,
            I => \N__9767\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__9774\,
            I => \N__9763\
        );

    \I__1204\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9756\
        );

    \I__1203\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9756\
        );

    \I__1202\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9756\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__9766\,
            I => \N__9753\
        );

    \I__1200\ : Span4Mux_v
    port map (
            O => \N__9763\,
            I => \N__9749\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__9756\,
            I => \N__9746\
        );

    \I__1198\ : InMux
    port map (
            O => \N__9753\,
            I => \N__9743\
        );

    \I__1197\ : InMux
    port map (
            O => \N__9752\,
            I => \N__9740\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__9749\,
            I => \c0.tx.o_Tx_Serial12\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__9746\,
            I => \c0.tx.o_Tx_Serial12\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__9743\,
            I => \c0.tx.o_Tx_Serial12\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__9740\,
            I => \c0.tx.o_Tx_Serial12\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__9731\,
            I => \c0.tx.N_294_cascade_\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9725\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__9725\,
            I => \c0.tx.m5_0_0\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9718\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9715\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9718\,
            I => \c0.tx.N_287\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9715\,
            I => \c0.tx.N_287\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__9710\,
            I => \c0.tx.N_288_cascade_\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__9704\,
            I => \blink_counterZ0Z_17\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9701\,
            I => blink_counter_cry_16
        );

    \I__1181\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9695\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__9695\,
            I => \blink_counterZ0Z_18\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9692\,
            I => blink_counter_cry_17
        );

    \I__1178\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__9686\,
            I => \blink_counterZ0Z_19\
        );

    \I__1176\ : InMux
    port map (
            O => \N__9683\,
            I => blink_counter_cry_18
        );

    \I__1175\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9677\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__9677\,
            I => \blink_counterZ0Z_20\
        );

    \I__1173\ : InMux
    port map (
            O => \N__9674\,
            I => blink_counter_cry_19
        );

    \I__1172\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9668\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__1170\ : Span4Mux_h
    port map (
            O => \N__9665\,
            I => \N__9661\
        );

    \I__1169\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9658\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__9661\,
            I => \blink_counterZ0Z_21\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__9658\,
            I => \blink_counterZ0Z_21\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9653\,
            I => blink_counter_cry_20
        );

    \I__1165\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9644\
        );

    \I__1164\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9644\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__9641\,
            I => \N__9637\
        );

    \I__1161\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9634\
        );

    \I__1160\ : Odrv4
    port map (
            O => \N__9637\,
            I => \blink_counterZ0Z_22\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__9634\,
            I => \blink_counterZ0Z_22\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9629\,
            I => blink_counter_cry_21
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__9626\,
            I => \N__9623\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9620\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1154\ : Span4Mux_v
    port map (
            O => \N__9617\,
            I => \N__9613\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9610\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__9613\,
            I => \blink_counterZ0Z_23\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__9610\,
            I => \blink_counterZ0Z_23\
        );

    \I__1150\ : InMux
    port map (
            O => \N__9605\,
            I => blink_counter_cry_22
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__9602\,
            I => \N__9599\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9593\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9598\,
            I => \N__9593\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9593\,
            I => \N__9590\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__9590\,
            I => \N__9586\
        );

    \I__1144\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9583\
        );

    \I__1143\ : Odrv4
    port map (
            O => \N__9586\,
            I => \blink_counterZ0Z_24\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9583\,
            I => \blink_counterZ0Z_24\
        );

    \I__1141\ : InMux
    port map (
            O => \N__9578\,
            I => \bfn_6_23_0_\
        );

    \I__1140\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9572\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__9572\,
            I => \blink_counterZ0Z_9\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9569\,
            I => blink_counter_cry_8
        );

    \I__1137\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9563\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__9563\,
            I => \blink_counterZ0Z_10\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9560\,
            I => blink_counter_cry_9
        );

    \I__1134\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9554\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9554\,
            I => \blink_counterZ0Z_11\
        );

    \I__1132\ : InMux
    port map (
            O => \N__9551\,
            I => blink_counter_cry_10
        );

    \I__1131\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9545\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__9545\,
            I => \blink_counterZ0Z_12\
        );

    \I__1129\ : InMux
    port map (
            O => \N__9542\,
            I => blink_counter_cry_11
        );

    \I__1128\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__9536\,
            I => \blink_counterZ0Z_13\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9533\,
            I => blink_counter_cry_12
        );

    \I__1125\ : InMux
    port map (
            O => \N__9530\,
            I => \N__9527\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__9527\,
            I => \blink_counterZ0Z_14\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9524\,
            I => blink_counter_cry_13
        );

    \I__1122\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9518\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__9518\,
            I => \blink_counterZ0Z_15\
        );

    \I__1120\ : InMux
    port map (
            O => \N__9515\,
            I => blink_counter_cry_14
        );

    \I__1119\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9509\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__9509\,
            I => \blink_counterZ0Z_16\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9506\,
            I => \bfn_6_22_0_\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__9500\,
            I => \blink_counterZ0Z_0\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9497\,
            I => \bfn_6_20_0_\
        );

    \I__1113\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__9491\,
            I => \blink_counterZ0Z_1\
        );

    \I__1111\ : InMux
    port map (
            O => \N__9488\,
            I => blink_counter_cry_0
        );

    \I__1110\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9482\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__9482\,
            I => \blink_counterZ0Z_2\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9479\,
            I => blink_counter_cry_1
        );

    \I__1107\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9473\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__9473\,
            I => \blink_counterZ0Z_3\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9470\,
            I => blink_counter_cry_2
        );

    \I__1104\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__9464\,
            I => \blink_counterZ0Z_4\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9461\,
            I => blink_counter_cry_3
        );

    \I__1101\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__9455\,
            I => \blink_counterZ0Z_5\
        );

    \I__1099\ : InMux
    port map (
            O => \N__9452\,
            I => blink_counter_cry_4
        );

    \I__1098\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__9446\,
            I => \blink_counterZ0Z_6\
        );

    \I__1096\ : InMux
    port map (
            O => \N__9443\,
            I => blink_counter_cry_5
        );

    \I__1095\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__9437\,
            I => \blink_counterZ0Z_7\
        );

    \I__1093\ : InMux
    port map (
            O => \N__9434\,
            I => blink_counter_cry_6
        );

    \I__1092\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9428\,
            I => \blink_counterZ0Z_8\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9425\,
            I => \bfn_6_21_0_\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9422\,
            I => \c0.tx.un1_r_Clock_Count_cry_0\
        );

    \I__1088\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9416\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__9416\,
            I => \c0.tx.r_Clock_Count_RNO_0Z0Z_2\
        );

    \I__1086\ : InMux
    port map (
            O => \N__9413\,
            I => \c0.tx.un1_r_Clock_Count_cry_1\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9410\,
            I => \c0.tx.un1_r_Clock_Count_cry_2\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__9407\,
            I => \c0.tx.r_Clock_Count_RNO_0Z0Z_3_cascade_\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9401\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__9401\,
            I => \c0.tx.r_Clock_Count_RNO_0Z0Z_0\
        );

    \I__1081\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9394\
        );

    \I__1080\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9391\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__9394\,
            I => \c0.tx.r_Clock_CountZ0Z_0\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__9391\,
            I => \c0.tx.r_Clock_CountZ0Z_0\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__9386\,
            I => \N__9382\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9379\
        );

    \I__1075\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9376\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__9379\,
            I => \c0.tx.r_Clock_Count_0_sqmuxa\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9376\,
            I => \c0.tx.r_Clock_Count_0_sqmuxa\
        );

    \I__1072\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9368\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9368\,
            I => \c0.tx.r_Clock_Count_RNO_0Z0Z_1\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__9365\,
            I => \c0.rx.g0_i_a4_0_3_cascade_\
        );

    \I__1069\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9356\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9361\,
            I => \N__9353\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9348\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9348\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__9356\,
            I => \c0.rx.r_Clock_Count14_3\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9353\,
            I => \c0.rx.r_Clock_Count14_3\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9348\,
            I => \c0.rx.r_Clock_Count14_3\
        );

    \I__1062\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9338\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9338\,
            I => \c0.rx.N_13\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9331\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9328\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__9331\,
            I => \N__9322\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__9328\,
            I => \N__9322\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__9327\,
            I => \N__9316\
        );

    \I__1055\ : Span4Mux_h
    port map (
            O => \N__9322\,
            I => \N__9309\
        );

    \I__1054\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9306\
        );

    \I__1053\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9297\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9319\,
            I => \N__9297\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9316\,
            I => \N__9297\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9297\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9292\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9313\,
            I => \N__9292\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9312\,
            I => \N__9289\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__9309\,
            I => \c0.rx.r_Clock_Count26\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9306\,
            I => \c0.rx.r_Clock_Count26\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__9297\,
            I => \c0.rx.r_Clock_Count26\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9292\,
            I => \c0.rx.r_Clock_Count26\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__9289\,
            I => \c0.rx.r_Clock_Count26\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__9278\,
            I => \N__9272\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__9277\,
            I => \N__9269\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__9276\,
            I => \N__9266\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__9275\,
            I => \N__9259\
        );

    \I__1037\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9255\
        );

    \I__1036\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9252\
        );

    \I__1035\ : InMux
    port map (
            O => \N__9266\,
            I => \N__9249\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__9265\,
            I => \N__9244\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__9264\,
            I => \N__9236\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__9263\,
            I => \N__9229\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__9262\,
            I => \N__9226\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9259\,
            I => \N__9220\
        );

    \I__1029\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9220\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__9255\,
            I => \N__9217\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__9252\,
            I => \N__9214\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__9249\,
            I => \N__9211\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9204\
        );

    \I__1024\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9204\
        );

    \I__1023\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9204\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__9243\,
            I => \N__9201\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__9242\,
            I => \N__9197\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__9241\,
            I => \N__9192\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__9240\,
            I => \N__9188\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9185\
        );

    \I__1017\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9180\
        );

    \I__1016\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9180\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9175\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9175\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9166\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9166\
        );

    \I__1011\ : InMux
    port map (
            O => \N__9226\,
            I => \N__9166\
        );

    \I__1010\ : InMux
    port map (
            O => \N__9225\,
            I => \N__9166\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9220\,
            I => \N__9161\
        );

    \I__1008\ : Span4Mux_h
    port map (
            O => \N__9217\,
            I => \N__9161\
        );

    \I__1007\ : Span4Mux_h
    port map (
            O => \N__9214\,
            I => \N__9156\
        );

    \I__1006\ : Span4Mux_h
    port map (
            O => \N__9211\,
            I => \N__9156\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__9204\,
            I => \N__9153\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9201\,
            I => \N__9144\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9200\,
            I => \N__9144\
        );

    \I__1002\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9144\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9196\,
            I => \N__9144\
        );

    \I__1000\ : InMux
    port map (
            O => \N__9195\,
            I => \N__9135\
        );

    \I__999\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9135\
        );

    \I__998\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9135\
        );

    \I__997\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9135\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9185\,
            I => \c0.rx.r_SM_MainZ0Z_2\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__9180\,
            I => \c0.rx.r_SM_MainZ0Z_2\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__9175\,
            I => \c0.rx.r_SM_MainZ0Z_2\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__9166\,
            I => \c0.rx.r_SM_MainZ0Z_2\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__9161\,
            I => \c0.rx.r_SM_MainZ0Z_2\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__9156\,
            I => \c0.rx.r_SM_MainZ0Z_2\
        );

    \I__990\ : Odrv4
    port map (
            O => \N__9153\,
            I => \c0.rx.r_SM_MainZ0Z_2\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__9144\,
            I => \c0.rx.r_SM_MainZ0Z_2\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__9135\,
            I => \c0.rx.r_SM_MainZ0Z_2\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__9116\,
            I => \c0.rx.r_Rx_DV_1_sqmuxa_cascade_\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__9113\,
            I => \N__9110\
        );

    \I__985\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9104\
        );

    \I__984\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9101\
        );

    \I__983\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9098\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__9107\,
            I => \N__9089\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9085\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__9101\,
            I => \N__9079\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__9098\,
            I => \N__9079\
        );

    \I__978\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9065\
        );

    \I__977\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9065\
        );

    \I__976\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9062\
        );

    \I__975\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9051\
        );

    \I__974\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9051\
        );

    \I__973\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9051\
        );

    \I__972\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9051\
        );

    \I__971\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9051\
        );

    \I__970\ : Span4Mux_h
    port map (
            O => \N__9085\,
            I => \N__9048\
        );

    \I__969\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9045\
        );

    \I__968\ : Span4Mux_h
    port map (
            O => \N__9079\,
            I => \N__9042\
        );

    \I__967\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9031\
        );

    \I__966\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9031\
        );

    \I__965\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9031\
        );

    \I__964\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9031\
        );

    \I__963\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9031\
        );

    \I__962\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9022\
        );

    \I__961\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9022\
        );

    \I__960\ : InMux
    port map (
            O => \N__9071\,
            I => \N__9022\
        );

    \I__959\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9022\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9065\,
            I => \c0.rx.r_SM_MainZ0Z_1\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__9062\,
            I => \c0.rx.r_SM_MainZ0Z_1\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__9051\,
            I => \c0.rx.r_SM_MainZ0Z_1\
        );

    \I__955\ : Odrv4
    port map (
            O => \N__9048\,
            I => \c0.rx.r_SM_MainZ0Z_1\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9045\,
            I => \c0.rx.r_SM_MainZ0Z_1\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__9042\,
            I => \c0.rx.r_SM_MainZ0Z_1\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9031\,
            I => \c0.rx.r_SM_MainZ0Z_1\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__9022\,
            I => \c0.rx.r_SM_MainZ0Z_1\
        );

    \I__950\ : InMux
    port map (
            O => \N__9005\,
            I => \N__9000\
        );

    \I__949\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8997\
        );

    \I__948\ : InMux
    port map (
            O => \N__9003\,
            I => \N__8982\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__9000\,
            I => \N__8977\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__8997\,
            I => \N__8977\
        );

    \I__945\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8974\
        );

    \I__944\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8969\
        );

    \I__943\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8969\
        );

    \I__942\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8966\
        );

    \I__941\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8957\
        );

    \I__940\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8957\
        );

    \I__939\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8957\
        );

    \I__938\ : InMux
    port map (
            O => \N__8989\,
            I => \N__8957\
        );

    \I__937\ : InMux
    port map (
            O => \N__8988\,
            I => \N__8948\
        );

    \I__936\ : InMux
    port map (
            O => \N__8987\,
            I => \N__8948\
        );

    \I__935\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8948\
        );

    \I__934\ : InMux
    port map (
            O => \N__8985\,
            I => \N__8948\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__8982\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__932\ : Odrv4
    port map (
            O => \N__8977\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__8974\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__8969\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__8966\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__8957\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__8948\,
            I => \c0.rx.r_SM_MainZ0Z_0\
        );

    \I__926\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8925\
        );

    \I__925\ : InMux
    port map (
            O => \N__8932\,
            I => \N__8925\
        );

    \I__924\ : InMux
    port map (
            O => \N__8931\,
            I => \N__8922\
        );

    \I__923\ : InMux
    port map (
            O => \N__8930\,
            I => \N__8919\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__8925\,
            I => \c0.rx.r_Clock_Count14\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__8922\,
            I => \c0.rx.r_Clock_Count14\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__8919\,
            I => \c0.rx.r_Clock_Count14\
        );

    \I__919\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__8909\,
            I => \c0.rx.N_9\
        );

    \I__917\ : InMux
    port map (
            O => \N__8906\,
            I => \N__8902\
        );

    \I__916\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8896\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__8902\,
            I => \N__8890\
        );

    \I__914\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8883\
        );

    \I__913\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8883\
        );

    \I__912\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8883\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8896\,
            I => \N__8880\
        );

    \I__910\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8873\
        );

    \I__909\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8870\
        );

    \I__908\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8867\
        );

    \I__907\ : Span4Mux_s3_h
    port map (
            O => \N__8890\,
            I => \N__8860\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__8883\,
            I => \N__8860\
        );

    \I__905\ : Span4Mux_h
    port map (
            O => \N__8880\,
            I => \N__8860\
        );

    \I__904\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8855\
        );

    \I__903\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8855\
        );

    \I__902\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8852\
        );

    \I__901\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8849\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8873\,
            I => \c0.rx.r_Clock_CountZ0Z_0\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__8870\,
            I => \c0.rx.r_Clock_CountZ0Z_0\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__8867\,
            I => \c0.rx.r_Clock_CountZ0Z_0\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__8860\,
            I => \c0.rx.r_Clock_CountZ0Z_0\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__8855\,
            I => \c0.rx.r_Clock_CountZ0Z_0\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__8852\,
            I => \c0.rx.r_Clock_CountZ0Z_0\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__8849\,
            I => \c0.rx.r_Clock_CountZ0Z_0\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__8834\,
            I => \N__8828\
        );

    \I__892\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8822\
        );

    \I__891\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8818\
        );

    \I__890\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8813\
        );

    \I__889\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8813\
        );

    \I__888\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8808\
        );

    \I__887\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8808\
        );

    \I__886\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8802\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__8822\,
            I => \N__8799\
        );

    \I__884\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8796\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__8818\,
            I => \N__8789\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__8813\,
            I => \N__8789\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__8808\,
            I => \N__8789\
        );

    \I__880\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8784\
        );

    \I__879\ : InMux
    port map (
            O => \N__8806\,
            I => \N__8784\
        );

    \I__878\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8781\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__8802\,
            I => \c0.rx.r_Clock_CountZ0Z_1\
        );

    \I__876\ : Odrv4
    port map (
            O => \N__8799\,
            I => \c0.rx.r_Clock_CountZ0Z_1\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__8796\,
            I => \c0.rx.r_Clock_CountZ0Z_1\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__8789\,
            I => \c0.rx.r_Clock_CountZ0Z_1\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__8784\,
            I => \c0.rx.r_Clock_CountZ0Z_1\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__8781\,
            I => \c0.rx.r_Clock_CountZ0Z_1\
        );

    \I__871\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8765\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__8765\,
            I => \c0.rx.r_Clock_Count14_1\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__868\ : InMux
    port map (
            O => \N__8759\,
            I => \N__8756\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__8756\,
            I => \c0.rx.N_12_0\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__8753\,
            I => \c0.rx.N_9_0_cascade_\
        );

    \I__865\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8744\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__8744\,
            I => \c0.rx.N_11_i\
        );

    \I__862\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8737\
        );

    \I__861\ : InMux
    port map (
            O => \N__8740\,
            I => \N__8733\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__8737\,
            I => \N__8730\
        );

    \I__859\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8727\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__8733\,
            I => \c0.rx.r_Clock_CountZ0Z_6\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__8730\,
            I => \c0.rx.r_Clock_CountZ0Z_6\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__8727\,
            I => \c0.rx.r_Clock_CountZ0Z_6\
        );

    \I__855\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8716\
        );

    \I__854\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8713\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__8716\,
            I => \N__8710\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8713\,
            I => \N__8705\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__8710\,
            I => \N__8702\
        );

    \I__850\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8699\
        );

    \I__849\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8696\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__8705\,
            I => \c0.rx.r_Clock_CountZ0Z_5\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__8702\,
            I => \c0.rx.r_Clock_CountZ0Z_5\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__8699\,
            I => \c0.rx.r_Clock_CountZ0Z_5\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8696\,
            I => \c0.rx.r_Clock_CountZ0Z_5\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__843\ : InMux
    port map (
            O => \N__8684\,
            I => \N__8680\
        );

    \I__842\ : InMux
    port map (
            O => \N__8683\,
            I => \N__8677\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__8680\,
            I => \N__8674\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__8677\,
            I => \c0.rx.r_Clock_CountZ0Z_7\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__8674\,
            I => \c0.rx.r_Clock_CountZ0Z_7\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__8669\,
            I => \N__8663\
        );

    \I__837\ : InMux
    port map (
            O => \N__8668\,
            I => \N__8658\
        );

    \I__836\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8655\
        );

    \I__835\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8652\
        );

    \I__834\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8649\
        );

    \I__833\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8646\
        );

    \I__832\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8643\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8658\,
            I => \c0.rx.r_Clock_CountZ0Z_4\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8655\,
            I => \c0.rx.r_Clock_CountZ0Z_4\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__8652\,
            I => \c0.rx.r_Clock_CountZ0Z_4\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__8649\,
            I => \c0.rx.r_Clock_CountZ0Z_4\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__8646\,
            I => \c0.rx.r_Clock_CountZ0Z_4\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__8643\,
            I => \c0.rx.r_Clock_CountZ0Z_4\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__8630\,
            I => \c0.rx.r_Clock_Count14_3_cascade_\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__8627\,
            I => \c0.rx.r_Clock_Count26_cascade_\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__8624\,
            I => \N__8617\
        );

    \I__822\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8608\
        );

    \I__821\ : InMux
    port map (
            O => \N__8622\,
            I => \N__8605\
        );

    \I__820\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8602\
        );

    \I__819\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8599\
        );

    \I__818\ : InMux
    port map (
            O => \N__8617\,
            I => \N__8596\
        );

    \I__817\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8593\
        );

    \I__816\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8586\
        );

    \I__815\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8586\
        );

    \I__814\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8586\
        );

    \I__813\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8583\
        );

    \I__812\ : InMux
    port map (
            O => \N__8611\,
            I => \N__8580\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8608\,
            I => \c0.rx.r_Clock_CountZ0Z_2\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__8605\,
            I => \c0.rx.r_Clock_CountZ0Z_2\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__8602\,
            I => \c0.rx.r_Clock_CountZ0Z_2\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__8599\,
            I => \c0.rx.r_Clock_CountZ0Z_2\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8596\,
            I => \c0.rx.r_Clock_CountZ0Z_2\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8593\,
            I => \c0.rx.r_Clock_CountZ0Z_2\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__8586\,
            I => \c0.rx.r_Clock_CountZ0Z_2\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8583\,
            I => \c0.rx.r_Clock_CountZ0Z_2\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__8580\,
            I => \c0.rx.r_Clock_CountZ0Z_2\
        );

    \I__802\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8556\
        );

    \I__801\ : InMux
    port map (
            O => \N__8560\,
            I => \N__8550\
        );

    \I__800\ : InMux
    port map (
            O => \N__8559\,
            I => \N__8545\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8542\
        );

    \I__798\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8535\
        );

    \I__797\ : InMux
    port map (
            O => \N__8554\,
            I => \N__8535\
        );

    \I__796\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8535\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__8550\,
            I => \N__8532\
        );

    \I__794\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8529\
        );

    \I__793\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8524\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__8545\,
            I => \N__8513\
        );

    \I__791\ : Span4Mux_v
    port map (
            O => \N__8542\,
            I => \N__8513\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__8535\,
            I => \N__8513\
        );

    \I__789\ : Span4Mux_v
    port map (
            O => \N__8532\,
            I => \N__8513\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8513\
        );

    \I__787\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8508\
        );

    \I__786\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8508\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8524\,
            I => \c0.rx.r_Clock_CountZ0Z_3\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__8513\,
            I => \c0.rx.r_Clock_CountZ0Z_3\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__8508\,
            I => \c0.rx.r_Clock_CountZ0Z_3\
        );

    \I__782\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8495\
        );

    \I__781\ : InMux
    port map (
            O => \N__8500\,
            I => \N__8495\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__8495\,
            I => \c0.rx.r_Clock_Count_1_sqmuxa_0\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__8492\,
            I => \c0.rx.un1_r_Clock_Count_5_m_1_cascade_\
        );

    \I__778\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__8486\,
            I => \N_12\
        );

    \I__776\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__8480\,
            I => \N_8_0\
        );

    \I__774\ : IoInMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__8474\,
            I => \N__8471\
        );

    \I__772\ : Span4Mux_s0_v
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__771\ : Span4Mux_v
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__8465\,
            I => \LED_c\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__8462\,
            I => \c0.rx.CO1_cascade_\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__8459\,
            I => \c0.rx.g0_i_o3_0_4_cascade_\
        );

    \I__767\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__8453\,
            I => \c0.rx.N_10\
        );

    \I__765\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8447\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__8447\,
            I => \c0.rx.g1_4\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__8444\,
            I => \c0.rx.g1_5_cascade_\
        );

    \I__762\ : InMux
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__8438\,
            I => \c0.rx.g1\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__8435\,
            I => \c0.rx.g0_0_1_cascade_\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__8432\,
            I => \c0.rx.r_Clock_Count14_cascade_\
        );

    \I__758\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__8426\,
            I => \c0.rx.m6_ns_1\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__8423\,
            I => \c0.rx.un1_r_Clock_Count_5_m_0_cascade_\
        );

    \I__755\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8415\
        );

    \I__754\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8410\
        );

    \I__753\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8410\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__8415\,
            I => \c0.rx.un1_r_Clock_Count_2_sqmuxa_0\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8410\,
            I => \c0.rx.un1_r_Clock_Count_2_sqmuxa_0\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__8405\,
            I => \c0.rx.N_7_cascade_\
        );

    \I__749\ : SRMux
    port map (
            O => \N__8402\,
            I => \N__8399\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__8399\,
            I => \N__8396\
        );

    \I__747\ : Span4Mux_h
    port map (
            O => \N__8396\,
            I => \N__8392\
        );

    \I__746\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8389\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__8392\,
            I => \c0.rx.r_SM_Main_RNICMJF6_0Z0Z_1\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__8389\,
            I => \c0.rx.r_SM_Main_RNICMJF6_0Z0Z_1\
        );

    \I__743\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8381\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__8381\,
            I => \c0.rx.N_10_0\
        );

    \I__741\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8375\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__8375\,
            I => \c0.rx.N_13_0\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__8372\,
            I => \c0.rx.N_12_1_cascade_\
        );

    \I__738\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8366\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__8366\,
            I => \c0.rx.un1_r_Clock_Count_5_c2\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__8363\,
            I => \c0.rx.N_6_cascade_\
        );

    \I__735\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8354\
        );

    \I__734\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8354\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8354\,
            I => \c0.rx.r_Clock_Count_2_sqmuxa_0\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__8351\,
            I => \c0.rx.r_Clock_Count_2_sqmuxa_0_cascade_\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__8348\,
            I => \c0.rx.g0_i_o4_0_1_cascade_\
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__8345\,
            I => \c0.rx.g0_i_o2_2_3_cascade_\
        );

    \I__729\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__8339\,
            I => \c0.rx.g0_i_a4_1_1\
        );

    \I__727\ : IoInMux
    port map (
            O => \N__8336\,
            I => \N__8333\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__725\ : Span4Mux_s0_v
    port map (
            O => \N__8330\,
            I => \N__8326\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__8329\,
            I => \N__8323\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__8326\,
            I => \N__8320\
        );

    \I__722\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8317\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__8320\,
            I => \PIN_1_c\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__8317\,
            I => \PIN_1_c\
        );

    \I__719\ : CEMux
    port map (
            O => \N__8312\,
            I => \N__8309\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__8309\,
            I => \N__8306\
        );

    \I__717\ : Odrv4
    port map (
            O => \N__8306\,
            I => \c0.rx.un1_r_Rx_DV7_0\
        );

    \I__716\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8300\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__8300\,
            I => \c0.rx.g0_i_o2_5\
        );

    \I__714\ : InMux
    port map (
            O => \N__8297\,
            I => \N__8294\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__8294\,
            I => \c0.rx.g0_i_o2_4\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__8291\,
            I => \N__8288\
        );

    \I__711\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8285\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__8285\,
            I => \c0.rx.g0_i_o2_6\
        );

    \I__709\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8279\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__8279\,
            I => \c0.rx.g0_i_a4_1_3\
        );

    \I__707\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8273\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8270\
        );

    \I__705\ : Odrv12
    port map (
            O => \N__8270\,
            I => \PIN_2_c\
        );

    \I__704\ : InMux
    port map (
            O => \N__8267\,
            I => \N__8264\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__8264\,
            I => \c0.rx.r_Rx_Data_RZ0\
        );

    \I__702\ : IoInMux
    port map (
            O => \N__8261\,
            I => \N__8258\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__8258\,
            I => \N__8255\
        );

    \I__700\ : IoSpan4Mux
    port map (
            O => \N__8255\,
            I => \N__8252\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__8252\,
            I => \c0.rx.rx_data_ready\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__8249\,
            I => \c0.rx.un1_r_Clock_Count_5_c2_cascade_\
        );

    \I__697\ : IoInMux
    port map (
            O => \N__8246\,
            I => \N__8243\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__8243\,
            I => \N__8240\
        );

    \I__695\ : IoSpan4Mux
    port map (
            O => \N__8240\,
            I => \N__8237\
        );

    \I__694\ : IoSpan4Mux
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__693\ : IoSpan4Mux
    port map (
            O => \N__8234\,
            I => \N__8231\
        );

    \I__692\ : Odrv4
    port map (
            O => \N__8231\,
            I => \CLK_ibuf_gb_io_gb_input\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_6_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_25_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.i12\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_5_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_25_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.data_cry_7\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_6_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_20_0_\
        );

    \IN_MUX_bfv_6_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => blink_counter_cry_7,
            carryinitout => \bfn_6_21_0_\
        );

    \IN_MUX_bfv_6_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => blink_counter_cry_15,
            carryinitout => \bfn_6_22_0_\
        );

    \IN_MUX_bfv_6_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => blink_counter_cry_23,
            carryinitout => \bfn_6_23_0_\
        );

    \CLK_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8246\,
            GLOBALBUFFEROUTPUT => \CLK_c_g\
        );

    \c0.rx.r_Rx_DV_e_RNIHVG2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8261\,
            GLOBALBUFFEROUTPUT => \c0.rx_data_ready_g\
        );

    \c0.byte_transmit_counter_RNIA0ET3_0_2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__16949\,
            GLOBALBUFFEROUTPUT => \c0.data_out_0__1_sqmuxa_g\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12278\,
            GLOBALBUFFEROUTPUT => \c0.data_in_frame_0__0_sqmuxa_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8267\,
            lcout => \c0.rx.r_Rx_DataZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_R_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8276\,
            lcout => \c0.rx.r_Rx_Data_RZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_e_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__9005\,
            in1 => \N__9109\,
            in2 => \N__9277\,
            in3 => \N__9335\,
            lcout => \c0.rx.rx_data_ready\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21824\,
            ce => \N__8312\,
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_1_7_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__8906\,
            in1 => \N__8720\,
            in2 => \N__9278\,
            in3 => \N__8667\,
            lcout => \c0.rx.g0_i_o2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_2_7_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__8621\,
            in1 => \N__8741\,
            in2 => \N__9113\,
            in3 => \N__8832\,
            lcout => \c0.rx.g0_i_o2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_7_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8993\,
            in2 => \_gnd_net_\,
            in3 => \N__8548\,
            lcout => \c0.rx.g0_i_o2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNIPDG17_1_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8831\,
            in1 => \N__8901\,
            in2 => \_gnd_net_\,
            in3 => \N__8420\,
            lcout => \c0.rx.un1_r_Clock_Count_5_c2\,
            ltout => \c0.rx.un1_r_Clock_Count_5_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_3_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__8622\,
            in1 => \N__8395\,
            in2 => \N__8249\,
            in3 => \N__8555\,
            lcout => \c0.rx.r_Clock_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21827\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_3_4_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9248\,
            in2 => \_gnd_net_\,
            in3 => \N__8900\,
            lcout => OPEN,
            ltout => \c0.rx.g0_i_o4_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_4_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__8827\,
            in1 => \N__8615\,
            in2 => \N__8348\,
            in3 => \N__8554\,
            lcout => \c0.rx.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_4_4_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8826\,
            in1 => \N__8342\,
            in2 => \N__9265\,
            in3 => \N__8613\,
            lcout => \c0.rx.g0_i_a4_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_3_5_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__8614\,
            in1 => \N__8899\,
            in2 => \N__8834\,
            in3 => \N__9247\,
            lcout => OPEN,
            ltout => \c0.rx.g0_i_o2_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_1_5_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100101010101"
        )
    port map (
            in0 => \N__8719\,
            in1 => \N__8553\,
            in2 => \N__8345\,
            in3 => \N__8666\,
            lcout => \c0.rx.N_11_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_2_2_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8879\,
            in1 => \N__8616\,
            in2 => \N__21193\,
            in3 => \N__8821\,
            lcout => \c0.rx.g1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_5_4_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8878\,
            in2 => \_gnd_net_\,
            in3 => \N__8662\,
            lcout => \c0.rx.g0_i_a4_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__10261\,
            in1 => \N__9956\,
            in2 => \N__8329\,
            in3 => \N__10403\,
            lcout => \PIN_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21842\,
            ce => 'H',
            sr => \N__9779\
        );

    \c0.rx.r_Rx_DV_e_RNO_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100011001"
        )
    port map (
            in0 => \N__9108\,
            in1 => \N__9004\,
            in2 => \N__9276\,
            in3 => \N__9334\,
            lcout => \c0.rx.un1_r_Rx_DV7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_7_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000001"
        )
    port map (
            in0 => \N__8303\,
            in1 => \N__8297\,
            in2 => \N__8291\,
            in3 => \N__8683\,
            lcout => \c0.rx.r_Clock_CountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21828\,
            ce => 'H',
            sr => \N__8402\
        );

    \c0.rx.r_Clock_Count_RNO_2_4_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__8282\,
            in1 => \N__8559\,
            in2 => \N__9107\,
            in3 => \N__9361\,
            lcout => \c0.rx.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_8_1_0__m6_ns_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110001110111"
        )
    port map (
            in0 => \N__9320\,
            in1 => \N__9094\,
            in2 => \N__10850\,
            in3 => \N__8429\,
            lcout => OPEN,
            ltout => \c0.rx.N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_0_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__9232\,
            in1 => \_gnd_net_\,
            in2 => \N__8405\,
            in3 => \_gnd_net_\,
            lcout => \c0.rx.r_SM_MainZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNICMJF6_0_1_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__8359\,
            in1 => \N__9225\,
            in2 => \N__9327\,
            in3 => \N__9088\,
            lcout => \c0.rx.r_SM_Main_RNICMJF6_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_1_4_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__9093\,
            in1 => \N__8996\,
            in2 => \N__9263\,
            in3 => \N__9319\,
            lcout => OPEN,
            ltout => \c0.rx.N_12_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_4_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__8384\,
            in1 => \N__8378\,
            in2 => \N__8372\,
            in3 => \N__8668\,
            lcout => \c0.rx.r_Clock_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_2_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__9092\,
            in1 => \N__9315\,
            in2 => \N__9262\,
            in3 => \N__8360\,
            lcout => OPEN,
            ltout => \c0.rx.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_2_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101100000"
        )
    port map (
            in0 => \N__8623\,
            in1 => \N__8369\,
            in2 => \N__8363\,
            in3 => \N__8441\,
            lcout => \c0.rx.r_Clock_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNIHR7E3_1_0_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9070\,
            in1 => \N__8985\,
            in2 => \N__9240\,
            in3 => \N__8930\,
            lcout => \c0.rx.r_Clock_Count_2_sqmuxa_0\,
            ltout => \c0.rx.r_Clock_Count_2_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNICMJF6_1_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__9084\,
            in1 => \N__9191\,
            in2 => \N__8351\,
            in3 => \N__9312\,
            lcout => \c0.rx.un1_r_Clock_Count_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_3_2_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9072\,
            in1 => \N__8986\,
            in2 => \N__9241\,
            in3 => \N__8528\,
            lcout => OPEN,
            ltout => \c0.rx.g1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_1_2_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__8450\,
            in1 => \_gnd_net_\,
            in2 => \N__8444\,
            in3 => \N__9360\,
            lcout => \c0.rx.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNIGQSH_3_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8527\,
            in2 => \_gnd_net_\,
            in3 => \N__8805\,
            lcout => OPEN,
            ltout => \c0.rx.g0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNICMJ72_2_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8611\,
            in1 => \N__8877\,
            in2 => \N__8435\,
            in3 => \N__9359\,
            lcout => \c0.rx.r_Clock_Count14\,
            ltout => \c0.rx.r_Clock_Count14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_8_1_0__m6_ns_1_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__9071\,
            in1 => \N__21194\,
            in2 => \N__8432\,
            in3 => \N__8987\,
            lcout => \c0.rx.m6_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_RNIIGH91_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8988\,
            in1 => \N__9195\,
            in2 => \N__21213\,
            in3 => \N__9073\,
            lcout => \c0.rx.r_Clock_Count_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_0_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000110011"
        )
    port map (
            in0 => \N__9258\,
            in1 => \N__8418\,
            in2 => \_gnd_net_\,
            in3 => \N__8894\,
            lcout => OPEN,
            ltout => \c0.rx.un1_r_Clock_Count_5_m_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_0_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8500\,
            in2 => \N__8423\,
            in3 => \N__8932\,
            lcout => \c0.rx.r_Clock_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_1_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000100100010"
        )
    port map (
            in0 => \N__8895\,
            in1 => \N__8419\,
            in2 => \N__9275\,
            in3 => \N__8825\,
            lcout => OPEN,
            ltout => \c0.rx.un1_r_Clock_Count_5_m_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_1_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8501\,
            in2 => \N__8492\,
            in3 => \N__8933\,
            lcout => \c0.rx.r_Clock_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_obuf_RNO_0_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__9649\,
            in1 => \N__9598\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_obuf_RNO_1_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__9811\,
            in1 => \N__9650\,
            in2 => \N__9602\,
            in3 => \N__9671\,
            lcout => \N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_obuf_RNO_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100010101"
        )
    port map (
            in0 => \N__8489\,
            in1 => \N__8483\,
            in2 => \N__9626\,
            in3 => \N__9812\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_RNO_0_2_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21410\,
            in1 => \N__21304\,
            in2 => \_gnd_net_\,
            in3 => \N__21096\,
            lcout => OPEN,
            ltout => \c0.rx.CO1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_2_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9924\,
            in2 => \N__8462\,
            in3 => \N__21452\,
            lcout => \c0.rx.r_Bit_IndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_6_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110000100011"
        )
    port map (
            in0 => \N__9234\,
            in1 => \N__8456\,
            in2 => \N__8762\,
            in3 => \N__8740\,
            lcout => \c0.rx.r_Clock_CountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_2_6_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__8905\,
            in1 => \N__8709\,
            in2 => \N__8669\,
            in3 => \N__9233\,
            lcout => OPEN,
            ltout => \c0.rx.g0_i_o3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_6_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__8620\,
            in1 => \N__8561\,
            in2 => \N__8459\,
            in3 => \N__8833\,
            lcout => \c0.rx.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNI55K61_0_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__8991\,
            in1 => \_gnd_net_\,
            in2 => \N__9242\,
            in3 => \N__9075\,
            lcout => \c0.rx.r_Rx_DV6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_1_6_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8990\,
            lcout => \c0.rx.N_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_2_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__9314\,
            in1 => \N__9078\,
            in2 => \N__9243\,
            in3 => \N__9003\,
            lcout => \c0.rx.r_SM_MainZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_0_5_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9077\,
            in1 => \N__8992\,
            in2 => \_gnd_net_\,
            in3 => \N__9313\,
            lcout => OPEN,
            ltout => \c0.rx.N_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_5_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__9200\,
            in1 => \N__9341\,
            in2 => \N__8753\,
            in3 => \N__8750\,
            lcout => \c0.rx.r_Clock_CountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNIE3Q31_7_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8736\,
            in1 => \N__8708\,
            in2 => \N__8687\,
            in3 => \N__8661\,
            lcout => \c0.rx.r_Clock_Count14_3\,
            ltout => \c0.rx.r_Clock_Count14_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNICMJ72_3_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__8612\,
            in1 => \N__8768\,
            in2 => \N__8630\,
            in3 => \N__8549\,
            lcout => \c0.rx.r_Clock_Count26\,
            ltout => \c0.rx.r_Clock_Count26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNIHR7E3_0_0_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__9074\,
            in1 => \N__9196\,
            in2 => \N__8627\,
            in3 => \N__8989\,
            lcout => \c0.rx.r_Rx_Byte_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_4_5_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8807\,
            in1 => \N__8893\,
            in2 => \N__8624\,
            in3 => \N__8560\,
            lcout => OPEN,
            ltout => \c0.rx.g0_i_a4_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNO_2_5_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9235\,
            in1 => \N__9095\,
            in2 => \N__9365\,
            in3 => \N__9362\,
            lcout => \c0.rx.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_RNIHR7E3_0_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__9096\,
            in1 => \N__8994\,
            in2 => \N__9264\,
            in3 => \N__9321\,
            lcout => OPEN,
            ltout => \c0.rx.r_Rx_DV_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_1_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000100"
        )
    port map (
            in0 => \N__9239\,
            in1 => \N__9097\,
            in2 => \N__9116\,
            in3 => \N__8912\,
            lcout => \c0.rx.r_SM_MainZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_8_1_0__m8_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8995\,
            in1 => \N__21214\,
            in2 => \_gnd_net_\,
            in3 => \N__8931\,
            lcout => \c0.rx.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count_RNIDNSH_1_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8876\,
            in2 => \_gnd_net_\,
            in3 => \N__8806\,
            lcout => \c0.rx.r_Clock_Count14_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_0_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__9728\,
            in1 => \N__10045\,
            in2 => \N__10409\,
            in3 => \N__9785\,
            lcout => \c0.tx.r_SM_MainZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_2_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__10260\,
            in1 => \N__9419\,
            in2 => \N__9766\,
            in3 => \N__10318\,
            lcout => \c0.tx.r_Clock_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_0_c_inv_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__13360\,
            in1 => \N__9397\,
            in2 => \_gnd_net_\,
            in3 => \N__9884\,
            lcout => \c0.tx.r_Clock_Count_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_RNO_0_0_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9398\,
            in2 => \N__9386\,
            in3 => \N__9385\,
            lcout => \c0.tx.r_Clock_Count_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_25_0_\,
            carryout => \c0.tx.un1_r_Clock_Count_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_RNO_0_1_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9872\,
            in2 => \_gnd_net_\,
            in3 => \N__9422\,
            lcout => \c0.tx.r_Clock_Count_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \c0.tx.un1_r_Clock_Count_cry_0\,
            carryout => \c0.tx.un1_r_Clock_Count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_RNO_0_2_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9854\,
            in2 => \_gnd_net_\,
            in3 => \N__9413\,
            lcout => \c0.tx.r_Clock_Count_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \c0.tx.un1_r_Clock_Count_cry_1\,
            carryout => \c0.tx.un1_r_Clock_Count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_RNO_0_3_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9836\,
            in2 => \_gnd_net_\,
            in3 => \N__9410\,
            lcout => OPEN,
            ltout => \c0.tx.r_Clock_Count_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_3_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__10246\,
            in1 => \N__9773\,
            in2 => \N__9407\,
            in3 => \N__10303\,
            lcout => \c0.tx.r_Clock_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_0_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__10301\,
            in1 => \N__10244\,
            in2 => \N__9777\,
            in3 => \N__9404\,
            lcout => \c0.tx.r_Clock_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNIFAME1_0_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__10402\,
            in1 => \N__10439\,
            in2 => \N__10259\,
            in3 => \N__10300\,
            lcout => \c0.tx.r_Clock_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count_1_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__10302\,
            in1 => \N__10245\,
            in2 => \N__9778\,
            in3 => \N__9371\,
            lcout => \c0.tx.r_Clock_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNID5VK2_21_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11587\,
            in1 => \N__11833\,
            in2 => \N__11064\,
            in3 => \N__11649\,
            lcout => \c0.nextCRC16_3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_5_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21395\,
            in1 => \N__21461\,
            in2 => \_gnd_net_\,
            in3 => \N__21295\,
            lcout => \c0.rx.r_Rx_Bytece_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_0_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9503\,
            in2 => \_gnd_net_\,
            in3 => \N__9497\,
            lcout => \blink_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_20_0_\,
            carryout => blink_counter_cry_0,
            clk => \N__21833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9494\,
            in2 => \_gnd_net_\,
            in3 => \N__9488\,
            lcout => \blink_counterZ0Z_1\,
            ltout => OPEN,
            carryin => blink_counter_cry_0,
            carryout => blink_counter_cry_1,
            clk => \N__21833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_2_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9485\,
            in2 => \_gnd_net_\,
            in3 => \N__9479\,
            lcout => \blink_counterZ0Z_2\,
            ltout => OPEN,
            carryin => blink_counter_cry_1,
            carryout => blink_counter_cry_2,
            clk => \N__21833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_3_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9476\,
            in2 => \_gnd_net_\,
            in3 => \N__9470\,
            lcout => \blink_counterZ0Z_3\,
            ltout => OPEN,
            carryin => blink_counter_cry_2,
            carryout => blink_counter_cry_3,
            clk => \N__21833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_4_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9467\,
            in2 => \_gnd_net_\,
            in3 => \N__9461\,
            lcout => \blink_counterZ0Z_4\,
            ltout => OPEN,
            carryin => blink_counter_cry_3,
            carryout => blink_counter_cry_4,
            clk => \N__21833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_5_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9458\,
            in2 => \_gnd_net_\,
            in3 => \N__9452\,
            lcout => \blink_counterZ0Z_5\,
            ltout => OPEN,
            carryin => blink_counter_cry_4,
            carryout => blink_counter_cry_5,
            clk => \N__21833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_6_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9449\,
            in2 => \_gnd_net_\,
            in3 => \N__9443\,
            lcout => \blink_counterZ0Z_6\,
            ltout => OPEN,
            carryin => blink_counter_cry_5,
            carryout => blink_counter_cry_6,
            clk => \N__21833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_7_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9440\,
            in2 => \_gnd_net_\,
            in3 => \N__9434\,
            lcout => \blink_counterZ0Z_7\,
            ltout => OPEN,
            carryin => blink_counter_cry_6,
            carryout => blink_counter_cry_7,
            clk => \N__21833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_8_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9431\,
            in2 => \_gnd_net_\,
            in3 => \N__9425\,
            lcout => \blink_counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_6_21_0_\,
            carryout => blink_counter_cry_8,
            clk => \N__21837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_9_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9575\,
            in2 => \_gnd_net_\,
            in3 => \N__9569\,
            lcout => \blink_counterZ0Z_9\,
            ltout => OPEN,
            carryin => blink_counter_cry_8,
            carryout => blink_counter_cry_9,
            clk => \N__21837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_10_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9566\,
            in2 => \_gnd_net_\,
            in3 => \N__9560\,
            lcout => \blink_counterZ0Z_10\,
            ltout => OPEN,
            carryin => blink_counter_cry_9,
            carryout => blink_counter_cry_10,
            clk => \N__21837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_11_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9557\,
            in2 => \_gnd_net_\,
            in3 => \N__9551\,
            lcout => \blink_counterZ0Z_11\,
            ltout => OPEN,
            carryin => blink_counter_cry_10,
            carryout => blink_counter_cry_11,
            clk => \N__21837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_12_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9548\,
            in2 => \_gnd_net_\,
            in3 => \N__9542\,
            lcout => \blink_counterZ0Z_12\,
            ltout => OPEN,
            carryin => blink_counter_cry_11,
            carryout => blink_counter_cry_12,
            clk => \N__21837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_13_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9539\,
            in2 => \_gnd_net_\,
            in3 => \N__9533\,
            lcout => \blink_counterZ0Z_13\,
            ltout => OPEN,
            carryin => blink_counter_cry_12,
            carryout => blink_counter_cry_13,
            clk => \N__21837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_14_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9530\,
            in2 => \_gnd_net_\,
            in3 => \N__9524\,
            lcout => \blink_counterZ0Z_14\,
            ltout => OPEN,
            carryin => blink_counter_cry_13,
            carryout => blink_counter_cry_14,
            clk => \N__21837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_15_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9521\,
            in2 => \_gnd_net_\,
            in3 => \N__9515\,
            lcout => \blink_counterZ0Z_15\,
            ltout => OPEN,
            carryin => blink_counter_cry_14,
            carryout => blink_counter_cry_15,
            clk => \N__21837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_16_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9512\,
            in2 => \_gnd_net_\,
            in3 => \N__9506\,
            lcout => \blink_counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_6_22_0_\,
            carryout => blink_counter_cry_16,
            clk => \N__21845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_17_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9707\,
            in2 => \_gnd_net_\,
            in3 => \N__9701\,
            lcout => \blink_counterZ0Z_17\,
            ltout => OPEN,
            carryin => blink_counter_cry_16,
            carryout => blink_counter_cry_17,
            clk => \N__21845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_18_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9698\,
            in2 => \_gnd_net_\,
            in3 => \N__9692\,
            lcout => \blink_counterZ0Z_18\,
            ltout => OPEN,
            carryin => blink_counter_cry_17,
            carryout => blink_counter_cry_18,
            clk => \N__21845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_19_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9689\,
            in2 => \_gnd_net_\,
            in3 => \N__9683\,
            lcout => \blink_counterZ0Z_19\,
            ltout => OPEN,
            carryin => blink_counter_cry_18,
            carryout => blink_counter_cry_19,
            clk => \N__21845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_20_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9680\,
            in2 => \_gnd_net_\,
            in3 => \N__9674\,
            lcout => \blink_counterZ0Z_20\,
            ltout => OPEN,
            carryin => blink_counter_cry_19,
            carryout => blink_counter_cry_20,
            clk => \N__21845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_21_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9664\,
            in2 => \_gnd_net_\,
            in3 => \N__9653\,
            lcout => \blink_counterZ0Z_21\,
            ltout => OPEN,
            carryin => blink_counter_cry_20,
            carryout => blink_counter_cry_21,
            clk => \N__21845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_22_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9640\,
            in2 => \_gnd_net_\,
            in3 => \N__9629\,
            lcout => \blink_counterZ0Z_22\,
            ltout => OPEN,
            carryin => blink_counter_cry_21,
            carryout => blink_counter_cry_22,
            clk => \N__21845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_23_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9616\,
            in2 => \_gnd_net_\,
            in3 => \N__9605\,
            lcout => \blink_counterZ0Z_23\,
            ltout => OPEN,
            carryin => blink_counter_cry_22,
            carryout => blink_counter_cry_23,
            clk => \N__21845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_24_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9589\,
            in2 => \_gnd_net_\,
            in3 => \N__9578\,
            lcout => \blink_counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_6_23_0_\,
            carryout => blink_counter_cry_24,
            clk => \N__21852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_25_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9799\,
            in2 => \_gnd_net_\,
            in3 => \N__9815\,
            lcout => \blink_counterZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_0_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000010100100"
        )
    port map (
            in0 => \N__9722\,
            in1 => \N__10369\,
            in2 => \N__9986\,
            in3 => \N__10328\,
            lcout => \c0.tx.r_Bit_IndexZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNIBPOV_0_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10240\,
            in1 => \N__10368\,
            in2 => \_gnd_net_\,
            in3 => \N__10453\,
            lcout => \c0.tx.o_Tx_Serial12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNIIR5L_0_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10253\,
            in2 => \_gnd_net_\,
            in3 => \N__10440\,
            lcout => \c0.tx.N_287\,
            ltout => \c0.tx.N_287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_7_1_0__m5_0_o2_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__9980\,
            in1 => \N__10021\,
            in2 => \N__9788\,
            in3 => \N__10304\,
            lcout => \c0.tx.N_294\,
            ltout => \c0.tx.N_294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_2_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9752\,
            in2 => \N__9731\,
            in3 => \N__10046\,
            lcout => \c0.tx.r_Bit_IndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_7_1_0__m5_0_0_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__10305\,
            in1 => \N__10254\,
            in2 => \N__10940\,
            in3 => \N__10441\,
            lcout => \c0.tx.m5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_RNO_0_1_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__9981\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10306\,
            lcout => OPEN,
            ltout => \c0.tx.N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_1_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100110001000"
        )
    port map (
            in0 => \N__10022\,
            in1 => \N__9721\,
            in2 => \N__9710\,
            in3 => \N__10407\,
            lcout => \c0.tx.r_Bit_IndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_5_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__19361\,
            in1 => \N__14558\,
            in2 => \N__10094\,
            in3 => \N__19238\,
            lcout => \c0.tx_data_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_0_c_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9883\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_25_0_\,
            carryout => \c0.tx.r_Clock_Count12_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_1_c_inv_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9860\,
            in2 => \N__13386\,
            in3 => \N__9871\,
            lcout => \c0.tx.r_Clock_Count_i_1\,
            ltout => OPEN,
            carryin => \c0.tx.r_Clock_Count12_cry_0\,
            carryout => \c0.tx.r_Clock_Count12_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_2_c_inv_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9842\,
            in2 => \N__13394\,
            in3 => \N__9853\,
            lcout => \c0.tx.r_Clock_Count_i_2\,
            ltout => OPEN,
            carryin => \c0.tx.r_Clock_Count12_cry_1\,
            carryout => \c0.tx.r_Clock_Count12_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_cry_3_c_inv_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9835\,
            in1 => \N__9824\,
            in2 => \N__13387\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx.r_Clock_Count_i_3\,
            ltout => OPEN,
            carryin => \c0.tx.r_Clock_Count12_cry_2\,
            carryout => \c0.tx.r_Clock_Count12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count12_THRU_LUT4_0_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9818\,
            lcout => \c0.tx.r_Clock_Count12_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__3_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21863\,
            ce => 'H',
            sr => \N__17347\
        );

    \c0.data_out_0__7_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13362\,
            lcout => \c0.d_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21863\,
            ce => 'H',
            sr => \N__17347\
        );

    \c0.data_out_3__3_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13363\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21863\,
            ce => 'H',
            sr => \N__17347\
        );

    \c0.data_out_0__2_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13388\,
            lcout => \c0.d_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21872\,
            ce => 'H',
            sr => \N__17346\
        );

    \c0.data_out_1__7_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13390\,
            lcout => \c0.d_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21872\,
            ce => 'H',
            sr => \N__17346\
        );

    \c0.data_out_1__3_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13389\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21872\,
            ce => 'H',
            sr => \N__17346\
        );

    \c0.data_out_2__2_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13391\,
            lcout => \c0.d_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21872\,
            ce => 'H',
            sr => \N__17346\
        );

    \c0.data_out_2__5_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13392\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21872\,
            ce => 'H',
            sr => \N__17346\
        );

    \c0.data_out_2__7_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13393\,
            lcout => \c0.d_2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21872\,
            ce => 'H',
            sr => \N__17346\
        );

    \c0.d_2_RNIIQK01_7_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16541\,
            in1 => \N__16494\,
            in2 => \_gnd_net_\,
            in3 => \N__10510\,
            lcout => \c0.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_1_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__21481\,
            in1 => \N__21396\,
            in2 => \_gnd_net_\,
            in3 => \N__21293\,
            lcout => OPEN,
            ltout => \c0.rx.r_Rx_Bytece_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_1_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__11332\,
            in1 => \N__21228\,
            in2 => \N__9893\,
            in3 => \N__21136\,
            lcout => \c0.rx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21838\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_5_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__21137\,
            in1 => \N__10783\,
            in2 => \N__21241\,
            in3 => \N__9890\,
            lcout => \c0.rx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21838\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_0_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9937\,
            in1 => \N__21294\,
            in2 => \_gnd_net_\,
            in3 => \N__21145\,
            lcout => \c0.rx.r_Bit_IndexZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_RNIRD3K_2_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21471\,
            in1 => \N__21363\,
            in2 => \_gnd_net_\,
            in3 => \N__21277\,
            lcout => \c0.rx.un1_r_Rx_Byte_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_1_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000110"
        )
    port map (
            in0 => \N__10397\,
            in1 => \N__10471\,
            in2 => \N__10262\,
            in3 => \N__10320\,
            lcout => \c0.tx.r_SM_MainZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_1_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__21278\,
            in1 => \N__9938\,
            in2 => \N__21390\,
            in3 => \N__21132\,
            lcout => \c0.rx.r_Bit_IndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_RNIFAME1_0_0_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__10378\,
            in1 => \N__10470\,
            in2 => \N__10255\,
            in3 => \N__10319\,
            lcout => OPEN,
            ltout => \c0.tx.r_Tx_Active_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10921\,
            in2 => \N__9911\,
            in3 => \N__14184\,
            lcout => \c0.tx_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_1_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__19398\,
            in1 => \N__19205\,
            in2 => \N__10865\,
            in3 => \N__14959\,
            lcout => \c0.tx_data_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_1_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__16876\,
            in1 => \N__9908\,
            in2 => \N__11039\,
            in3 => \N__10544\,
            lcout => \c0.tx.r_Tx_DataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21864\,
            ce => \N__10942\,
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_3_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__9902\,
            in1 => \N__10043\,
            in2 => \N__10061\,
            in3 => \N__10017\,
            lcout => OPEN,
            ltout => \c0.tx.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_1_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__10018\,
            in1 => \N__10955\,
            in2 => \N__9896\,
            in3 => \N__10076\,
            lcout => \c0.tx.N_354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_3_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__10052\,
            in1 => \N__17567\,
            in2 => \N__16882\,
            in3 => \N__10826\,
            lcout => OPEN,
            ltout => \c0.tx_data_1_0_i_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_3_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__16877\,
            in1 => \N__14705\,
            in2 => \N__10079\,
            in3 => \N__10535\,
            lcout => \c0.tx.r_Tx_DataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21864\,
            ce => \N__10942\,
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_5_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__16875\,
            in1 => \N__11090\,
            in2 => \N__10070\,
            in3 => \N__9944\,
            lcout => \c0.tx.r_Tx_DataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21864\,
            ce => \N__10942\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_3_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__19410\,
            in1 => \N__19209\,
            in2 => \N__11903\,
            in3 => \N__15332\,
            lcout => \c0.tx_data_RNO_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_4_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__10112\,
            in1 => \N__10044\,
            in2 => \N__10103\,
            in3 => \N__10019\,
            lcout => OPEN,
            ltout => \c0.tx.r_Tx_Data_pmux_3_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_2_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__10020\,
            in1 => \N__10985\,
            in2 => \N__9995\,
            in3 => \N__10973\,
            lcout => OPEN,
            ltout => \c0.tx.N_357_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_RNO_0_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000111"
        )
    port map (
            in0 => \N__9992\,
            in1 => \N__9985\,
            in2 => \N__9959\,
            in3 => \N__10472\,
            lcout => \c0.tx.N_320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_5_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__15170\,
            in1 => \N__11257\,
            in2 => \N__19232\,
            in3 => \N__19397\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_5_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__16868\,
            in1 => \N__17554\,
            in2 => \N__9947\,
            in3 => \N__12746\,
            lcout => \c0.tx_data_1_0_i_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_0_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__12839\,
            in1 => \N__17566\,
            in2 => \N__13436\,
            in3 => \N__16913\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_0_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110110011"
        )
    port map (
            in0 => \N__16883\,
            in1 => \N__11570\,
            in2 => \N__10115\,
            in3 => \N__11777\,
            lcout => \c0.tx.r_Tx_DataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21879\,
            ce => \N__10943\,
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_4_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__16881\,
            in1 => \N__10145\,
            in2 => \N__10880\,
            in3 => \N__11186\,
            lcout => \c0.tx.r_Tx_DataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21879\,
            ce => \N__10943\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__5_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10484\,
            in1 => \N__12038\,
            in2 => \_gnd_net_\,
            in3 => \N__12971\,
            lcout => \c0.data_out_7_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21887\,
            ce => \N__17298\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__3_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10652\,
            lcout => \c0.d_2_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21887\,
            ce => \N__17298\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__4_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10631\,
            lcout => \c0.d_2_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21897\,
            ce => \N__17297\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__3_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13927\,
            lcout => \c0.data_in_0_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21825\,
            ce => \N__22151\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_2_c_RNO_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13887\,
            in1 => \N__14082\,
            in2 => \N__12361\,
            in3 => \N__13659\,
            lcout => \c0.i12_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_1__4_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16197\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_1_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21834\,
            ce => \N__22150\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__7_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15946\,
            lcout => \c0.data_in_1_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21834\,
            ce => \N__22150\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__4_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11443\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_2_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21834\,
            ce => \N__22150\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_5_c_RNO_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18121\,
            in1 => \N__11419\,
            in2 => \N__16201\,
            in3 => \N__13755\,
            lcout => \c0.i12_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__0_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18301\,
            lcout => \c0.data_in_0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21839\,
            ce => \N__22152\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__1_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13847\,
            lcout => \c0.data_in_2_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21839\,
            ce => \N__22152\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__0_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18674\,
            lcout => \c0.data_in_2_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21839\,
            ce => \N__22152\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__5_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13867\,
            lcout => \c0.data_in_1_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21839\,
            ce => \N__22152\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__0_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13660\,
            lcout => \c0.data_in_1_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21839\,
            ce => \N__22152\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__5_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13891\,
            lcout => \c0.data_in_0_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21839\,
            ce => \N__22152\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__7_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12360\,
            lcout => \c0.data_in_0_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21847\,
            ce => \N__22155\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__2_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16227\,
            lcout => \c0.data_in_1_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21847\,
            ce => \N__22155\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__3_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15424\,
            lcout => \c0.data_in_1_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21847\,
            ce => \N__22155\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__3_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10130\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_7_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21847\,
            ce => \N__22155\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__1_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13756\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_1_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21847\,
            ce => \N__22155\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__2_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16645\,
            lcout => \c0.data_in_0_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21847\,
            ce => \N__22155\,
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_3_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21494\,
            in1 => \N__21411\,
            in2 => \_gnd_net_\,
            in3 => \N__21315\,
            lcout => OPEN,
            ltout => \c0.rx.r_Rx_Bytece_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_3_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__10129\,
            in1 => \N__21227\,
            in2 => \N__10133\,
            in3 => \N__21146\,
            lcout => \c0.rx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_2_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__16628\,
            in1 => \N__18925\,
            in2 => \N__19563\,
            in3 => \N__12500\,
            lcout => OPEN,
            ltout => \c0.tx2_data_RNO_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_2_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__10772\,
            in1 => \N__20354\,
            in2 => \N__10118\,
            in3 => \N__20939\,
            lcout => \c0.tx2_data_1_0_i_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__4_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13330\,
            lcout => \c0.d_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21865\,
            ce => 'H',
            sr => \N__17348\
        );

    \c0.tx.r_SM_Main_7_1_0__m5_0_a2_0_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10398\,
            in1 => \N__14207\,
            in2 => \N__10239\,
            in3 => \N__10468\,
            lcout => \c0.tx.r_Tx_Data_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_5_6_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__11703\,
            in1 => \N__19158\,
            in2 => \N__11995\,
            in3 => \N__17561\,
            lcout => \c0.m115_amcf1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_2_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__10469\,
            in1 => \N__10209\,
            in2 => \N__10408\,
            in3 => \N__10327\,
            lcout => \c0.tx.r_SM_MainZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_0_4_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11912\,
            in2 => \_gnd_net_\,
            in3 => \N__13016\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_3_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__4_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10160\,
            in1 => \N__12934\,
            in2 => \N__10163\,
            in3 => \N__12110\,
            lcout => \c0.data_out_6_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21880\,
            ce => \N__17300\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_1_4_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12144\,
            in1 => \N__14657\,
            in2 => \N__13432\,
            in3 => \N__10812\,
            lcout => \c0.nextCRC16_3_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_4_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__19362\,
            in1 => \N__10154\,
            in2 => \N__15017\,
            in3 => \N__19204\,
            lcout => \c0.tx_data_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_4__6_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10610\,
            lcout => \c0.d_2_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21880\,
            ce => \N__17300\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__1_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10577\,
            lcout => \c0.d_2_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21880\,
            ce => \N__17300\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_1_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__19203\,
            in1 => \N__12794\,
            in2 => \N__12148\,
            in3 => \N__19363\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_4Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_1_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__16867\,
            in1 => \N__17562\,
            in2 => \N__10547\,
            in3 => \N__12635\,
            lcout => \c0.tx_data_1_0_i_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_3_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__19402\,
            in1 => \N__19202\,
            in2 => \N__10520\,
            in3 => \N__10592\,
            lcout => \c0.tx_data_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_0_3_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11955\,
            in1 => \N__11076\,
            in2 => \_gnd_net_\,
            in3 => \N__12106\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_0_a2_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__3_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10813\,
            in1 => \N__12770\,
            in2 => \N__10523\,
            in3 => \N__11258\,
            lcout => \c0.data_out_6_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21888\,
            ce => \N__17299\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_7_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__19200\,
            in1 => \N__10511\,
            in2 => \N__12938\,
            in3 => \N__19403\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_7_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__16842\,
            in1 => \N__17553\,
            in2 => \N__10493\,
            in3 => \N__10490\,
            lcout => \c0.tx_data_1_0_i_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_7_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__19201\,
            in1 => \N__15286\,
            in2 => \N__15208\,
            in3 => \N__19401\,
            lcout => \c0.tx_data_RNO_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNI1DHT_19_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17418\,
            in1 => \N__17379\,
            in2 => \_gnd_net_\,
            in3 => \N__10591\,
            lcout => \c0.N_74\,
            ltout => \c0.N_74_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNITDBK1_47_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15195\,
            in2 => \N__10595\,
            in3 => \N__15166\,
            lcout => \c0.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_2__3_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13300\,
            lcout => \c0.d_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21898\,
            ce => 'H',
            sr => \N__17343\
        );

    \c0.d_2_RNINVK01_8_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10814\,
            in1 => \N__11249\,
            in2 => \_gnd_net_\,
            in3 => \N__11788\,
            lcout => \c0.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__0_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13299\,
            lcout => \c0.d_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21898\,
            ce => 'H',
            sr => \N__17343\
        );

    \c0.data_0_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11809\,
            in2 => \_gnd_net_\,
            in3 => \N__10580\,
            lcout => \c0.dataZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \c0.data_cry_0\,
            clk => \N__21906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_1_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10573\,
            in2 => \_gnd_net_\,
            in3 => \N__10562\,
            lcout => \c0.dataZ0Z_1\,
            ltout => OPEN,
            carryin => \c0.data_cry_0\,
            carryout => \c0.data_cry_1\,
            clk => \N__21906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_2_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11113\,
            in2 => \_gnd_net_\,
            in3 => \N__10559\,
            lcout => \c0.dataZ0Z_2\,
            ltout => OPEN,
            carryin => \c0.data_cry_1\,
            carryout => \c0.data_cry_2\,
            clk => \N__21906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_3_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11149\,
            in2 => \_gnd_net_\,
            in3 => \N__10556\,
            lcout => \c0.dataZ0Z_3\,
            ltout => OPEN,
            carryin => \c0.data_cry_2\,
            carryout => \c0.data_cry_3\,
            clk => \N__21906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_4_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11221\,
            in2 => \_gnd_net_\,
            in3 => \N__10553\,
            lcout => \c0.dataZ0Z_4\,
            ltout => OPEN,
            carryin => \c0.data_cry_3\,
            carryout => \c0.data_cry_4\,
            clk => \N__21906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_5_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11281\,
            in2 => \_gnd_net_\,
            in3 => \N__10550\,
            lcout => \c0.dataZ0Z_5\,
            ltout => OPEN,
            carryin => \c0.data_cry_4\,
            carryout => \c0.data_cry_5\,
            clk => \N__21906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_6_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11125\,
            in2 => \_gnd_net_\,
            in3 => \N__10667\,
            lcout => \c0.dataZ0Z_6\,
            ltout => OPEN,
            carryin => \c0.data_cry_5\,
            carryout => \c0.data_cry_6\,
            clk => \N__21906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_7_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11161\,
            in2 => \_gnd_net_\,
            in3 => \N__10664\,
            lcout => \c0.dataZ0Z_7\,
            ltout => OPEN,
            carryin => \c0.data_cry_6\,
            carryout => \c0.data_cry_7\,
            clk => \N__21906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_8_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11869\,
            in2 => \_gnd_net_\,
            in3 => \N__10661\,
            lcout => \c0.dataZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_28_0_\,
            carryout => \c0.data_cry_8\,
            clk => \N__21914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_9_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11209\,
            in2 => \_gnd_net_\,
            in3 => \N__10658\,
            lcout => \c0.dataZ0Z_9\,
            ltout => OPEN,
            carryin => \c0.data_cry_8\,
            carryout => \c0.data_cry_9\,
            clk => \N__21914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_10_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11137\,
            in2 => \_gnd_net_\,
            in3 => \N__10655\,
            lcout => \c0.dataZ0Z_10\,
            ltout => OPEN,
            carryin => \c0.data_cry_9\,
            carryout => \c0.data_cry_10\,
            clk => \N__21914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_11_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10645\,
            in2 => \_gnd_net_\,
            in3 => \N__10634\,
            lcout => \c0.dataZ0Z_11\,
            ltout => OPEN,
            carryin => \c0.data_cry_10\,
            carryout => \c0.data_cry_11\,
            clk => \N__21914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_12_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10627\,
            in2 => \_gnd_net_\,
            in3 => \N__10616\,
            lcout => \c0.dataZ0Z_12\,
            ltout => OPEN,
            carryin => \c0.data_cry_11\,
            carryout => \c0.data_cry_12\,
            clk => \N__21914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_13_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11269\,
            in2 => \_gnd_net_\,
            in3 => \N__10613\,
            lcout => \c0.dataZ0Z_13\,
            ltout => OPEN,
            carryin => \c0.data_cry_12\,
            carryout => \c0.data_cry_13\,
            clk => \N__21914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_14_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10606\,
            in2 => \_gnd_net_\,
            in3 => \N__10691\,
            lcout => \c0.dataZ0Z_14\,
            ltout => OPEN,
            carryin => \c0.data_cry_13\,
            carryout => \c0.data_cry_14\,
            clk => \N__21914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_15_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12244\,
            in2 => \_gnd_net_\,
            in3 => \N__10688\,
            lcout => \c0.dataZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21914\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__1_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.d_2_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21929\,
            ce => 'H',
            sr => \N__17339\
        );

    \c0.FRAME_MATCHER_i12_0_c_RNO_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12166\,
            in1 => \N__12373\,
            in2 => \N__13585\,
            in3 => \N__15472\,
            lcout => \c0.i12_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0__1_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15976\,
            lcout => \c0.data_in_0_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21829\,
            ce => \N__22154\,
            sr => \_gnd_net_\
        );

    \c0.data_in_0__4_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14086\,
            lcout => \c0.data_in_0_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21829\,
            ce => \N__22154\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_0_c_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10685\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \c0.i12_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_1_c_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10709\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_0\,
            carryout => \c0.i12_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_2_c_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10676\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_1\,
            carryout => \c0.i12_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_3_c_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10700\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_2\,
            carryout => \c0.i12_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_4_c_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10742\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_3\,
            carryout => \c0.i12_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_5_c_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10721\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_4\,
            carryout => \c0.i12_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_6_c_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10733\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_5\,
            carryout => \c0.i12_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_7_c_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11198\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.i12_6\,
            carryout => \c0.i12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_THRU_LUT4_0_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10712\,
            lcout => \c0.i12_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_3_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011101110"
        )
    port map (
            in0 => \N__20334\,
            in1 => \N__17759\,
            in2 => \N__14111\,
            in3 => \N__17870\,
            lcout => \c0.tx2_data_1_iv_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_1_c_RNO_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18297\,
            in1 => \N__15960\,
            in2 => \N__13923\,
            in3 => \N__17956\,
            lcout => \c0.i12_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_3_c_RNO_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15939\,
            in1 => \N__13863\,
            in2 => \N__16231\,
            in3 => \N__15423\,
            lcout => \c0.i12_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_3_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__20902\,
            in1 => \N__13550\,
            in2 => \_gnd_net_\,
            in3 => \N__15406\,
            lcout => \c0.tx2_data_1_iv_3_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_4_c_RNO_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16258\,
            in1 => \N__13678\,
            in2 => \N__12409\,
            in3 => \N__16644\,
            lcout => \c0.i12_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_2__2_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16737\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_2_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21848\,
            ce => \N__22156\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__3_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13804\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_2_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21848\,
            ce => \N__22156\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__5_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11396\,
            lcout => \c0.data_in_2_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21848\,
            ce => \N__22156\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__7_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12331\,
            lcout => \c0.data_in_2_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21848\,
            ce => \N__22156\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_6_c_RNO_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18666\,
            in1 => \N__13839\,
            in2 => \N__16741\,
            in3 => \N__13803\,
            lcout => \c0.i12_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_4__1_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13819\,
            lcout => \c0.data_in_4_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21855\,
            ce => \N__22158\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__3_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15844\,
            lcout => \c0.data_in_3_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21855\,
            ce => \N__22158\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__1_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16078\,
            lcout => \c0.data_in_3_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21855\,
            ce => \N__22158\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__0_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11320\,
            lcout => \c0.data_in_3_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21855\,
            ce => \N__22158\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__0_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15913\,
            lcout => \c0.data_in_4_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21855\,
            ce => \N__22158\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__0_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18782\,
            lcout => \c0.data_in_5_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21855\,
            ce => \N__22158\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__5_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10787\,
            lcout => \c0.data_in_7_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21855\,
            ce => \N__22158\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_2_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__22088\,
            in1 => \N__21992\,
            in2 => \N__19564\,
            in3 => \N__18923\,
            lcout => \c0.tx2_data_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_2_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__18921\,
            in1 => \N__16181\,
            in2 => \N__19539\,
            in3 => \N__16721\,
            lcout => \c0.tx2_data_RNO_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_2_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__18924\,
            in1 => \N__18411\,
            in2 => \N__19540\,
            in3 => \N__14165\,
            lcout => OPEN,
            ltout => \c0.tx2_data_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_2_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__20357\,
            in1 => \N__10766\,
            in2 => \N__10760\,
            in3 => \N__10757\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21861\,
            ce => \N__20745\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_1_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__16670\,
            in1 => \N__19523\,
            in2 => \N__22040\,
            in3 => \N__18922\,
            lcout => \c0.tx2_data_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_3_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100111111"
        )
    port map (
            in0 => \N__14120\,
            in1 => \N__10751\,
            in2 => \N__12188\,
            in3 => \N__20356\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21861\,
            ce => \N__20745\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_3_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__14435\,
            in1 => \N__16436\,
            in2 => \N__14292\,
            in3 => \N__11555\,
            lcout => \c0.tx2.r_Clock_CountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_7_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__10849\,
            in1 => \N__21122\,
            in2 => \N__18826\,
            in3 => \N__21218\,
            lcout => \c0.rx_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNI13HR_0_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__16366\,
            in1 => \N__14433\,
            in2 => \_gnd_net_\,
            in3 => \N__14354\,
            lcout => \c0.tx2.o_Tx_Serial12\,
            ltout => \c0.tx2.o_Tx_Serial12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_2_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__14434\,
            in1 => \N__11357\,
            in2 => \N__10829\,
            in3 => \N__16435\,
            lcout => \c0.tx2.r_Clock_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_3_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__12064\,
            in1 => \N__16516\,
            in2 => \N__19234\,
            in3 => \N__19411\,
            lcout => \c0.tx_data_RNO_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_2_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__21485\,
            in1 => \N__21391\,
            in2 => \_gnd_net_\,
            in3 => \N__21308\,
            lcout => \c0.rx.r_Rx_Bytece_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__6_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13249\,
            lcout => \c0.d_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21874\,
            ce => 'H',
            sr => \N__17345\
        );

    \c0.data_out_2__4_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13250\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21874\,
            ce => 'H',
            sr => \N__17345\
        );

    \c0.data_out_2__6_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13251\,
            lcout => \c0.d_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21874\,
            ce => 'H',
            sr => \N__17345\
        );

    \c0.tx_data_RNO_4_6_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15060\,
            in1 => \N__17540\,
            in2 => \_gnd_net_\,
            in3 => \N__10811\,
            lcout => OPEN,
            ltout => \c0.N_293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_6_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010111111111"
        )
    port map (
            in0 => \N__11009\,
            in1 => \N__19162\,
            in2 => \N__11000\,
            in3 => \N__19412\,
            lcout => \c0.tx_data_1_0_i_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_6_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__17563\,
            in1 => \N__14511\,
            in2 => \N__11748\,
            in3 => \N__16908\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_6_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110111011"
        )
    port map (
            in0 => \N__16869\,
            in1 => \N__10997\,
            in2 => \N__10988\,
            in3 => \N__16958\,
            lcout => \c0.tx.r_Tx_DataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21881\,
            ce => \N__10941\,
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_2_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__11615\,
            in1 => \N__16871\,
            in2 => \N__11021\,
            in3 => \N__14666\,
            lcout => \c0.tx.r_Tx_DataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21881\,
            ce => \N__10941\,
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_7_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__16870\,
            in1 => \N__11045\,
            in2 => \N__14681\,
            in3 => \N__10961\,
            lcout => \c0.tx.r_Tx_DataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21881\,
            ce => \N__10941\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_0_0_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__11739\,
            in1 => \N__11256\,
            in2 => \_gnd_net_\,
            in3 => \N__17435\,
            lcout => \c0.nextCRC16_3_0_a2_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_4_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__19372\,
            in1 => \N__11171\,
            in2 => \N__19237\,
            in3 => \N__13092\,
            lcout => \c0.tx_data_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__1_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11605\,
            in1 => \N__11849\,
            in2 => \N__11653\,
            in3 => \N__11078\,
            lcout => \c0.data_out_6_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21889\,
            ce => \N__17295\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_5_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__11604\,
            in1 => \N__19373\,
            in2 => \N__12887\,
            in3 => \N__19218\,
            lcout => \c0.tx_data_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_7_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__19374\,
            in1 => \N__12851\,
            in2 => \N__19235\,
            in3 => \N__11077\,
            lcout => \c0.tx_data_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_1_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__11956\,
            in1 => \N__19371\,
            in2 => \N__13127\,
            in3 => \N__19222\,
            lcout => \c0.tx_data_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_2_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__19375\,
            in1 => \N__11102\,
            in2 => \N__19236\,
            in3 => \N__13003\,
            lcout => \c0.tx_data_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__4_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13298\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21899\,
            ce => 'H',
            sr => \N__17342\
        );

    \c0.data_out_6__RNO_2_7_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14603\,
            in1 => \N__12124\,
            in2 => \N__13011\,
            in3 => \N__12098\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_0_a2_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_0_7_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11957\,
            in1 => \N__11907\,
            in2 => \N__11012\,
            in3 => \N__13046\,
            lcout => \c0.nextCRC16_3_0_a2_3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_3__2_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.d_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21899\,
            ce => 'H',
            sr => \N__17342\
        );

    \c0.tx_data_RNO_3_4_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__14860\,
            in1 => \N__16566\,
            in2 => \N__19233\,
            in3 => \N__19400\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_4_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__16843\,
            in1 => \N__17564\,
            in2 => \N__11189\,
            in3 => \N__11177\,
            lcout => \c0.tx_data_1_0_i_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_4_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__19213\,
            in1 => \N__12125\,
            in2 => \N__12020\,
            in3 => \N__19399\,
            lcout => \c0.tx_data_RNO_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__4_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12002\,
            in1 => \N__12838\,
            in2 => \N__14518\,
            in3 => \N__17378\,
            lcout => \c0.data_out_7_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21907\,
            ce => \N__17293\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__7_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11162\,
            lcout => \c0.d_2_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21907\,
            ce => \N__17293\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__3_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11150\,
            lcout => \c0.d_2_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21907\,
            ce => \N__17293\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__2_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11138\,
            lcout => \c0.d_2_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21907\,
            ce => \N__17293\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__6_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11126\,
            lcout => \c0.d_2_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21907\,
            ce => \N__17293\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__2_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11114\,
            lcout => \c0.d_2_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21907\,
            ce => \N__17293\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__2_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14557\,
            in1 => \N__14916\,
            in2 => \N__14519\,
            in3 => \N__12071\,
            lcout => \c0.data_out_7_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21907\,
            ce => \N__17293\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__5_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11282\,
            lcout => \c0.d_2_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21907\,
            ce => \N__17293\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__5_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11270\,
            lcout => \c0.d_2_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21915\,
            ce => \N__17291\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__4_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11222\,
            lcout => \c0.d_2_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21915\,
            ce => \N__17291\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__1_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11210\,
            lcout => \c0.d_2_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21915\,
            ce => \N__17291\,
            sr => \_gnd_net_\
        );

    \c0.data_out_1__6_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13349\,
            lcout => \c0.d_2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21923\,
            ce => 'H',
            sr => \N__17338\
        );

    \c0.data_in_0__6_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11418\,
            lcout => \c0.data_in_0_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21835\,
            ce => \N__22157\,
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNO_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11388\,
            in1 => \N__11436\,
            in2 => \N__13705\,
            in3 => \N__12324\,
            lcout => \c0.i12_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_3__4_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18511\,
            lcout => \c0.data_in_3_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21841\,
            ce => \N__22153\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__5_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20009\,
            lcout => \c0.data_in_3_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21841\,
            ce => \N__22153\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__6_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20555\,
            lcout => \c0.data_in_3_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21841\,
            ce => \N__22153\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__7_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18848\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_3_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21841\,
            ce => \N__22153\,
            sr => \_gnd_net_\
        );

    \c0.data_in_2__6_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13701\,
            lcout => \c0.data_in_2_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21841\,
            ce => \N__22153\,
            sr => \_gnd_net_\
        );

    \c0.data_in_1__6_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18114\,
            lcout => \c0.data_in_1_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21841\,
            ce => \N__22153\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__4_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18719\,
            lcout => \c0.data_in_4_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21841\,
            ce => \N__22153\,
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_2_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__19493\,
            in1 => \N__20333\,
            in2 => \N__20901\,
            in3 => \N__18896\,
            lcout => \c0.N_72_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNI0CLC_0_0_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__20332\,
            in1 => \N__20861\,
            in2 => \_gnd_net_\,
            in3 => \N__19488\,
            lcout => OPEN,
            ltout => \c0.g1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_active_RNIU1BT1_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19758\,
            in1 => \N__12232\,
            in2 => \N__11294\,
            in3 => \N__18895\,
            lcout => \c0.N_247_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_0_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12233\,
            in1 => \N__19759\,
            in2 => \_gnd_net_\,
            in3 => \N__11291\,
            lcout => OPEN,
            ltout => \c0.N_249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__19807\,
            in1 => \N__11300\,
            in2 => \N__11285\,
            in3 => \N__12284\,
            lcout => \c0.wait_for_transmissionZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21849\,
            ce => 'H',
            sr => \N__20045\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNI6ITQ_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__19793\,
            in1 => \N__17725\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_frame_0__0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_0_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__18910\,
            in1 => \N__15601\,
            in2 => \N__19502\,
            in3 => \N__15902\,
            lcout => \c0.tx2_data_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_1_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__18897\,
            in1 => \N__15782\,
            in2 => \N__16067\,
            in3 => \N__19492\,
            lcout => \c0.tx2_data_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIM5UG_0_19_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15595\,
            in1 => \N__15401\,
            in2 => \N__19961\,
            in3 => \N__17903\,
            lcout => \c0.g3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__0_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11321\,
            lcout => \c0.d_4_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21856\,
            ce => \N__21594\,
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_4_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__17744\,
            in1 => \N__18143\,
            in2 => \N__18536\,
            in3 => \N__17724\,
            lcout => \c0.g0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIM5UG_19_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17905\,
            in1 => \N__19954\,
            in2 => \N__15407\,
            in3 => \N__15597\,
            lcout => \c0.g3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_5_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001010000100"
        )
    port map (
            in0 => \N__15869\,
            in1 => \N__17691\,
            in2 => \N__13565\,
            in3 => \N__17660\,
            lcout => OPEN,
            ltout => \c0.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_1_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11345\,
            in2 => \N__11309\,
            in3 => \N__11306\,
            lcout => \c0.byte_transmit_counter2_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_6_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15596\,
            in1 => \N__15402\,
            in2 => \N__19962\,
            in3 => \N__17904\,
            lcout => OPEN,
            ltout => \c0.g3_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_3_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__15698\,
            in1 => \N__15734\,
            in2 => \N__11348\,
            in3 => \N__15818\,
            lcout => \c0.g0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_4__2_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11371\,
            lcout => \c0.data_in_4_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21862\,
            ce => \N__22159\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__3_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14065\,
            lcout => \c0.data_in_6_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21862\,
            ce => \N__22159\,
            sr => \_gnd_net_\
        );

    \c0.data_in_3__2_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13939\,
            lcout => \c0.data_in_3_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21862\,
            ce => \N__22159\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__1_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18809\,
            lcout => \c0.data_in_5_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21862\,
            ce => \N__22159\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__2_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22115\,
            lcout => \c0.data_in_5_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21862\,
            ce => \N__22159\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__1_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11339\,
            lcout => \c0.data_in_7_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21862\,
            ce => \N__22159\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__3_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14446\,
            lcout => \c0.data_in_4_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21862\,
            ce => \N__22159\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__3_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20631\,
            lcout => \c0.data_in_5_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21862\,
            ce => \N__22159\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIBANL_28_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17015\,
            in1 => \N__18956\,
            in2 => \N__14008\,
            in3 => \N__12598\,
            lcout => \c0.un1_data_in_7__2_0_a2_0_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__4_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11444\,
            lcout => \c0.d_4_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21867\,
            ce => \N__21599\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__6_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11420\,
            lcout => \c0.d_4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21867\,
            ce => \N__21599\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__5_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11395\,
            lcout => \c0.d_4_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21867\,
            ce => \N__21599\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI7BIA_29_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22200\,
            in1 => \_gnd_net_\,
            in2 => \N__17023\,
            in3 => \N__17127\,
            lcout => \c0.un1_data_in_6__7_0_a2_17_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__4_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18718\,
            lcout => \c0.d_4_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21867\,
            ce => \N__21599\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__2_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11372\,
            lcout => \c0.d_4_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21867\,
            ce => \N__21599\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_RNO_0_0_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11528\,
            in2 => \N__11549\,
            in3 => \N__11548\,
            lcout => \c0.tx2.r_Clock_Count_RNO_0_0_0\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \c0.tx2.un1_r_Clock_Count_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_RNO_0_1_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11498\,
            in2 => \_gnd_net_\,
            in3 => \N__11360\,
            lcout => \c0.tx2.r_Clock_Count_RNO_0_0_1\,
            ltout => OPEN,
            carryin => \c0.tx2.un1_r_Clock_Count_cry_0\,
            carryout => \c0.tx2.un1_r_Clock_Count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_RNO_0_2_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11480\,
            in2 => \_gnd_net_\,
            in3 => \N__11351\,
            lcout => \c0.tx2.r_Clock_Count_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \c0.tx2.un1_r_Clock_Count_cry_1\,
            carryout => \c0.tx2.un1_r_Clock_Count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_RNO_0_3_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11462\,
            in2 => \_gnd_net_\,
            in3 => \N__11558\,
            lcout => \c0.tx2.r_Clock_Count_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNINID81_0_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__16365\,
            in1 => \N__14350\,
            in2 => \N__14432\,
            in3 => \N__16420\,
            lcout => \c0.tx2.r_Clock_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_0_c_inv_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__13348\,
            in1 => \N__11527\,
            in2 => \_gnd_net_\,
            in3 => \N__11510\,
            lcout => \c0.tx2.r_Clock_Count_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_0_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__14419\,
            in1 => \N__11534\,
            in2 => \N__14293\,
            in3 => \N__16421\,
            lcout => \c0.tx2.r_Clock_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count_1_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__16422\,
            in1 => \N__14420\,
            in2 => \N__14291\,
            in3 => \N__11516\,
            lcout => \c0.tx2.r_Clock_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_0_c_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11509\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \c0.tx2.r_Clock_Count12_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_1_c_inv_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11486\,
            in2 => \N__13301\,
            in3 => \N__11497\,
            lcout => \c0.tx2.r_Clock_Count_i_1\,
            ltout => OPEN,
            carryin => \c0.tx2.r_Clock_Count12_cry_0\,
            carryout => \c0.tx2.r_Clock_Count12_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_2_c_inv_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11468\,
            in2 => \N__13303\,
            in3 => \N__11479\,
            lcout => \c0.tx2.r_Clock_Count_i_2\,
            ltout => OPEN,
            carryin => \c0.tx2.r_Clock_Count12_cry_1\,
            carryout => \c0.tx2.r_Clock_Count12_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_cry_3_c_inv_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11461\,
            in1 => \N__11450\,
            in2 => \N__13302\,
            in3 => \_gnd_net_\,
            lcout => \c0.tx2.r_Clock_Count_i_3\,
            ltout => OPEN,
            carryin => \c0.tx2.r_Clock_Count12_cry_2\,
            carryout => \c0.tx2.r_Clock_Count12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Clock_Count12_THRU_LUT4_0_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11657\,
            lcout => \c0.tx2.r_Clock_Count12_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__1_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13260\,
            lcout => \c0.d_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21882\,
            ce => 'H',
            sr => \N__17344\
        );

    \c0.data_out_1__2_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13261\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21882\,
            ce => 'H',
            sr => \N__17344\
        );

    \c0.data_out_6__2_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12932\,
            in1 => \N__12790\,
            in2 => \N__11762\,
            in3 => \N__11654\,
            lcout => \c0.data_out_6_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21890\,
            ce => \N__17296\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_2_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__15106\,
            in1 => \N__19185\,
            in2 => \N__11624\,
            in3 => \N__19370\,
            lcout => \c0.tx_data_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__7_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11709\,
            in1 => \N__11609\,
            in2 => \N__16478\,
            in3 => \N__11675\,
            lcout => \c0.data_out_7_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21890\,
            ce => \N__17296\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_0_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__15135\,
            in1 => \N__16808\,
            in2 => \N__12105\,
            in3 => \N__17521\,
            lcout => OPEN,
            ltout => \c0.tx_data_1_iv_i_m2_0_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_0_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__16809\,
            in1 => \N__11798\,
            in2 => \N__11576\,
            in3 => \N__11822\,
            lcout => OPEN,
            ltout => \c0.N_304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_0_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19396\,
            in2 => \N__11573\,
            in3 => \N__19214\,
            lcout => \c0.tx_data_1_iv_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__0_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15023\,
            in1 => \N__11723\,
            in2 => \N__11858\,
            in3 => \N__11848\,
            lcout => \c0.data_out_6_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21900\,
            ce => \N__17294\,
            sr => \_gnd_net_\
        );

    \c0.data_out_5__0_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11816\,
            lcout => \c0.d_2_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21900\,
            ce => \N__17294\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__0_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11768\,
            in1 => \N__12701\,
            in2 => \N__13190\,
            in3 => \N__13147\,
            lcout => \c0.data_out_7_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21900\,
            ce => \N__17294\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_0_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__11792\,
            in1 => \N__17565\,
            in2 => \N__13064\,
            in3 => \N__16909\,
            lcout => \c0.tx_data_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_0_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__15098\,
            in1 => \_gnd_net_\,
            in2 => \N__15246\,
            in3 => \N__12034\,
            lcout => \c0.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_0_2_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16568\,
            in1 => \N__11750\,
            in2 => \_gnd_net_\,
            in3 => \N__13418\,
            lcout => \c0.nextCRC16_3_0_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_2_0_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__15308\,
            in1 => \_gnd_net_\,
            in2 => \N__15062\,
            in3 => \N__12828\,
            lcout => \c0.nextCRC16_3_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIQ3DA1_20_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11749\,
            in1 => \N__15021\,
            in2 => \N__13425\,
            in3 => \N__11716\,
            lcout => OPEN,
            ltout => \c0.nextCRC16_3_0_a2_6_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIKDAK6_20_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12769\,
            in1 => \N__11687\,
            in2 => \N__11678\,
            in3 => \N__11671\,
            lcout => \c0.N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIM3JT_12_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12149\,
            in1 => \N__12123\,
            in2 => \_gnd_net_\,
            in3 => \N__12097\,
            lcout => \c0.N_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__RNO_1_7_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12967\,
            in1 => \N__14550\,
            in2 => \N__14921\,
            in3 => \N__14501\,
            lcout => \c0.nextCRC16_3_0_a2_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_2_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15055\,
            in1 => \N__12820\,
            in2 => \N__11996\,
            in3 => \N__13070\,
            lcout => \c0.nextCRC16_3_0_a2_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNI6EK01_3_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15126\,
            in1 => \N__15350\,
            in2 => \_gnd_net_\,
            in3 => \N__12065\,
            lcout => \c0.N_75\,
            ltout => \c0.N_75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIJ2812_44_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15247\,
            in1 => \N__15105\,
            in2 => \N__12023\,
            in3 => \N__12013\,
            lcout => \c0.N_95\,
            ltout => \c0.N_95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIJDOU2_14_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15056\,
            in1 => \N__11991\,
            in2 => \N__11960\,
            in3 => \N__12821\,
            lcout => \c0.nextCRC16_3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNII92R1_27_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11954\,
            in1 => \N__11911\,
            in2 => \N__14731\,
            in3 => \N__14569\,
            lcout => \c0.N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_4__0_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11873\,
            lcout => \c0.d_2_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21924\,
            ce => \N__17289\,
            sr => \_gnd_net_\
        );

    \c0.data_out_4__7_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12248\,
            lcout => \c0.d_2_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21924\,
            ce => \N__17289\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Active_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__20749\,
            in1 => \N__12231\,
            in2 => \_gnd_net_\,
            in3 => \N__12647\,
            lcout => \c0.tx2_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21840\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_5_7_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__20924\,
            in1 => \N__12206\,
            in2 => \_gnd_net_\,
            in3 => \N__18218\,
            lcout => \c0.tx2_data_1_iv_5_1_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_7_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101111111"
        )
    port map (
            in0 => \N__18044\,
            in1 => \N__20925\,
            in2 => \N__20411\,
            in3 => \N__18335\,
            lcout => OPEN,
            ltout => \c0.tx2_data_1_iv_5_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_7_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111110000"
        )
    port map (
            in0 => \N__12215\,
            in1 => \N__20408\,
            in2 => \N__12209\,
            in3 => \N__20339\,
            lcout => \c0.tx2_data_1_iv_5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__7_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22205\,
            lcout => \c0.data_in_frame_6_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21850\,
            ce => \N__21586\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_3_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__12200\,
            in1 => \N__20407\,
            in2 => \_gnd_net_\,
            in3 => \N__20338\,
            lcout => \c0.tx2_data_1_iv_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__3_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12173\,
            lcout => \c0.d_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21850\,
            ce => \N__21586\,
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNI94LS6_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__19792\,
            in1 => \N__12155\,
            in2 => \_gnd_net_\,
            in3 => \N__13478\,
            lcout => \c0.wait_for_transmission_RNI94LSZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIT2KP_20_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19726\,
            in1 => \N__18334\,
            in2 => \N__18781\,
            in3 => \N__14158\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__0_0_a2_5_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI2LMH1_6_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18004\,
            in1 => \N__18182\,
            in2 => \N__12308\,
            in3 => \N__15460\,
            lcout => \c0.un1_data_in_6__0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI4CPT_18_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13545\,
            in1 => \N__16180\,
            in2 => \N__21980\,
            in3 => \N__16063\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__4_0_a2_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIHG3O1_16_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12422\,
            in2 => \N__12305\,
            in3 => \N__12467\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__4_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIK1Q66_10_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__14132\,
            in1 => \N__15995\,
            in2 => \N__12302\,
            in3 => \N__12299\,
            lcout => \c0.wait_for_transmission4_12_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIF73E2_14_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17184\,
            in1 => \N__16717\,
            in2 => \N__14024\,
            in3 => \N__13783\,
            lcout => OPEN,
            ltout => \c0.d_4_RNIF73E2Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIMKFE3_14_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__12434\,
            in1 => \_gnd_net_\,
            in2 => \N__12293\,
            in3 => \N__14803\,
            lcout => OPEN,
            ltout => \c0.d_4_RNIMKFE3Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIOL9I8_10_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15550\,
            in1 => \N__16103\,
            in2 => \N__12290\,
            in3 => \N__15811\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIB4H0M_43_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17627\,
            in1 => \N__17605\,
            in2 => \N__12287\,
            in3 => \N__17587\,
            lcout => \c0.wait_for_transmission4_12\,
            ltout => \c0.wait_for_transmission4_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNI61KS81_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12265\,
            in1 => \N__13442\,
            in2 => \N__12251\,
            in3 => \N__13454\,
            lcout => \c0.tx2_transmit_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIFCG72_32_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15594\,
            in1 => \N__12386\,
            in2 => \_gnd_net_\,
            in3 => \N__12392\,
            lcout => \c0.N_129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI46QL_16_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13635\,
            in1 => \N__17128\,
            in2 => \N__13969\,
            in3 => \N__12491\,
            lcout => \c0.un1_data_in_7__4_0_a2_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__2_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12413\,
            lcout => \c0.d_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21868\,
            ce => \N__21595\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNID6K21_0_15_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17901\,
            in1 => \N__12487\,
            in2 => \N__17941\,
            in3 => \N__12600\,
            lcout => \c0.d_4_RNID6K21_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNID6K21_15_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12599\,
            in1 => \N__17937\,
            in2 => \N__12496\,
            in3 => \N__17902\,
            lcout => \c0.d_4_RNID6K21Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__1_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12380\,
            lcout => \c0.d_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21868\,
            ce => \N__21595\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__7_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12362\,
            lcout => \c0.d_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21868\,
            ce => \N__21595\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__7_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12332\,
            lcout => \c0.d_4_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21868\,
            ce => \N__21595\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI9UF4_32_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15593\,
            in2 => \_gnd_net_\,
            in3 => \N__17900\,
            lcout => \c0.N_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_7__RNI74HC_1_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22056\,
            in2 => \_gnd_net_\,
            in3 => \N__17125\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__1_0_a2_24_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI716J_16_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18412\,
            in1 => \N__13642\,
            in2 => \N__12503\,
            in3 => \N__17171\,
            lcout => \c0.wait_for_transmission4_13_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNID6C91_1_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12492\,
            in1 => \N__12463\,
            in2 => \N__15723\,
            in3 => \N__12601\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__1_0_a2_24_a2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI8S283_14_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14009\,
            in1 => \N__12452\,
            in2 => \N__12446\,
            in3 => \N__12440\,
            lcout => \c0.wait_for_transmission4_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIJ6E4_27_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18957\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__1_0_a2_24_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIVMA91_17_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13546\,
            in1 => \N__13738\,
            in2 => \N__12443\,
            in3 => \N__15618\,
            lcout => \c0.un1_data_in_7__1_0_a2_24_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNITCRC_29_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17126\,
            in1 => \N__22201\,
            in2 => \N__18423\,
            in3 => \N__17022\,
            lcout => \c0.d_4_RNITCRCZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_0_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__18928\,
            in1 => \N__18648\,
            in2 => \N__19574\,
            in3 => \N__13643\,
            lcout => OPEN,
            ltout => \c0.tx2_data_RNO_4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_0_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__20342\,
            in1 => \N__13601\,
            in2 => \N__12425\,
            in3 => \N__20941\,
            lcout => OPEN,
            ltout => \c0.tx2_data_1_0_i_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_0_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12539\,
            in1 => \N__12623\,
            in2 => \N__12611\,
            in3 => \N__20344\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21883\,
            ce => \N__20741\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_1_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__19572\,
            in1 => \N__18257\,
            in2 => \N__12608\,
            in3 => \N__18927\,
            lcout => OPEN,
            ltout => \c0.tx2_data_RNO_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_1_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__20942\,
            in1 => \N__12545\,
            in2 => \N__12575\,
            in3 => \N__20343\,
            lcout => OPEN,
            ltout => \c0.tx2_data_1_0_i_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_1_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__20345\,
            in1 => \N__12572\,
            in2 => \N__12560\,
            in3 => \N__12557\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21883\,
            ce => \N__20741\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_1_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__18926\,
            in1 => \N__13739\,
            in2 => \N__19573\,
            in3 => \N__16031\,
            lcout => \c0.tx2_data_RNO_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_0_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__16754\,
            in1 => \N__19568\,
            in2 => \N__16583\,
            in3 => \N__18929\,
            lcout => \c0.tx2_data_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_2_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__16306\,
            in1 => \N__12533\,
            in2 => \N__14744\,
            in3 => \N__12515\,
            lcout => \c0.tx2.N_349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_4_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__12521\,
            in1 => \N__14225\,
            in2 => \N__20768\,
            in3 => \N__16304\,
            lcout => \c0.tx2.r_Tx_Data_pmux_3_i_m2_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_3_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__16305\,
            in1 => \N__16982\,
            in2 => \N__14233\,
            in3 => \N__12509\,
            lcout => OPEN,
            ltout => \c0.tx2.r_Tx_Data_pmux_6_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_1_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__17081\,
            in1 => \N__12695\,
            in2 => \N__12683\,
            in3 => \N__16307\,
            lcout => OPEN,
            ltout => \c0.tx2.N_346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_RNO_0_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__16461\,
            in1 => \N__12680\,
            in2 => \N__12674\,
            in3 => \N__14343\,
            lcout => OPEN,
            ltout => \c0.tx2.N_279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.o_Tx_Serial_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__14408\,
            in1 => \N__12664\,
            in2 => \N__12671\,
            in3 => \N__16349\,
            lcout => \PIN_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21891\,
            ce => 'H',
            sr => \N__14287\
        );

    \c0.tx2.r_SM_Main_RNINID81_0_0_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__14342\,
            in1 => \N__16348\,
            in2 => \N__14429\,
            in3 => \N__16423\,
            lcout => \c0.tx2.r_Tx_Active_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_2_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__16352\,
            in1 => \N__14349\,
            in2 => \N__14431\,
            in3 => \N__16434\,
            lcout => \c0.tx2.r_SM_MainZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_1_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__19168\,
            in1 => \N__14889\,
            in2 => \N__17392\,
            in3 => \N__19322\,
            lcout => \c0.tx_data_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_7_1_0__m5_0_0_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__14409\,
            in1 => \N__14347\,
            in2 => \N__20715\,
            in3 => \N__16432\,
            lcout => OPEN,
            ltout => \c0.tx2.m5_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_0_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__14234\,
            in1 => \N__16350\,
            in2 => \N__12626\,
            in3 => \N__14300\,
            lcout => \c0.tx2.r_SM_MainZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_1_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000110"
        )
    port map (
            in0 => \N__16351\,
            in1 => \N__14348\,
            in2 => \N__14430\,
            in3 => \N__16433\,
            lcout => \c0.tx2.r_SM_MainZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21901\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIGMI01_10_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12933\,
            in1 => \N__14641\,
            in2 => \_gnd_net_\,
            in3 => \N__12786\,
            lcout => \c0.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_5_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__19321\,
            in1 => \N__19169\,
            in2 => \N__13037\,
            in3 => \N__12731\,
            lcout => \c0.tx_data_RNO_4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIFMJ01_45_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12730\,
            in1 => \N__14939\,
            in2 => \_gnd_net_\,
            in3 => \N__14843\,
            lcout => \c0.N_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__4_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13351\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => 'H',
            sr => \N__17341\
        );

    \c0.data_out_2__1_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13352\,
            lcout => \c0.d_2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => 'H',
            sr => \N__17341\
        );

    \c0.data_out_3__5_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13353\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => 'H',
            sr => \N__17341\
        );

    \c0.data_out_0__1_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13350\,
            lcout => \c0.d_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => 'H',
            sr => \N__17341\
        );

    \c0.data_out_3__6_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13354\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21908\,
            ce => 'H',
            sr => \N__17341\
        );

    \c0.data_out_7__RNO_1_0_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14899\,
            in1 => \N__12707\,
            in2 => \N__14505\,
            in3 => \N__12944\,
            lcout => \c0.nextCRC16_3_0_a2_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_2_RNIK3C71_13_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13094\,
            in1 => \N__13004\,
            in2 => \N__14629\,
            in3 => \N__13029\,
            lcout => \c0.nextCRC16_3_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_1__5_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21916\,
            ce => 'H',
            sr => \N__17340\
        );

    \c0.data_out_7__RNO_1_2_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13093\,
            in1 => \N__15360\,
            in2 => \N__14628\,
            in3 => \N__13060\,
            lcout => \c0.nextCRC16_3_0_a2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_0__0_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13355\,
            lcout => \c0.d_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21916\,
            ce => 'H',
            sr => \N__17340\
        );

    \c0.d_2_RNIIJMM_15_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15282\,
            in2 => \_gnd_net_\,
            in3 => \N__13059\,
            lcout => \c0.nextCRC16_3_4_0\,
            ltout => \c0.nextCRC16_3_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_3_0_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13030\,
            in1 => \N__13012\,
            in2 => \N__12974\,
            in3 => \N__12960\,
            lcout => \c0.nextCRC16_3_0_a2_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__5_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14618\,
            in1 => \N__12919\,
            in2 => \_gnd_net_\,
            in3 => \N__13179\,
            lcout => \c0.data_out_6_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21925\,
            ce => \N__17290\,
            sr => \_gnd_net_\
        );

    \c0.data_out_6__7_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__12872\,
            in1 => \N__13159\,
            in2 => \N__12866\,
            in3 => \N__13143\,
            lcout => \c0.data_out_6_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21925\,
            ce => \N__17290\,
            sr => \_gnd_net_\
        );

    \c0.data_out_2__0_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13358\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21930\,
            ce => 'H',
            sr => \N__17337\
        );

    \c0.data_out_3__7_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13359\,
            lcout => \c0.d_2_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21930\,
            ce => 'H',
            sr => \N__17337\
        );

    \c0.data_out_3__0_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.d_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21930\,
            ce => 'H',
            sr => \N__17337\
        );

    \c0.data_out_0__5_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13357\,
            lcout => \c0.d_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21930\,
            ce => 'H',
            sr => \N__17337\
        );

    \c0.data_out_7__1_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13186\,
            in1 => \N__13163\,
            in2 => \N__14825\,
            in3 => \N__13148\,
            lcout => \c0.data_out_7_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21931\,
            ce => \N__17287\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_5_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101111111"
        )
    port map (
            in0 => \N__17856\,
            in1 => \N__20926\,
            in2 => \N__13112\,
            in3 => \N__13510\,
            lcout => \c0.tx2_data_1_0_i_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__5_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19967\,
            lcout => \c0.data_in_frame_7_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21857\,
            ce => \N__21583\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__5_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19985\,
            lcout => \c0.d_4_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21857\,
            ce => \N__21583\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_7_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101101111111"
        )
    port map (
            in0 => \N__20927\,
            in1 => \N__17857\,
            in2 => \N__13103\,
            in3 => \N__15524\,
            lcout => \c0.tx2_data_1_0_i_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__7_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22238\,
            lcout => \c0.data_in_frame_7_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21857\,
            ce => \N__21583\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__7_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20666\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_4_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21857\,
            ce => \N__21583\,
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_10_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17999\,
            in1 => \N__15390\,
            in2 => \N__15527\,
            in3 => \N__15456\,
            lcout => OPEN,
            ltout => \c0.wait_for_transmission_RNOZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_8_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15557\,
            in1 => \N__16247\,
            in2 => \N__13568\,
            in3 => \N__18590\,
            lcout => \c0.g0_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI5L571_45_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13725\,
            in1 => \N__13544\,
            in2 => \N__13514\,
            in3 => \N__15628\,
            lcout => \c0.N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI8A8H_26_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18429\,
            in1 => \N__16716\,
            in2 => \N__13496\,
            in3 => \N__17188\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__7_0_a2_17_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI6CFJ4_26_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13782\,
            in1 => \N__14799\,
            in2 => \N__13481\,
            in3 => \N__15808\,
            lcout => \c0.un1_data_in_6__7_0_a2_17_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIU7HB6_19_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000100"
        )
    port map (
            in0 => \N__18062\,
            in1 => \N__15680\,
            in2 => \N__13472\,
            in3 => \N__15809\,
            lcout => \c0.g0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIIVJN_13_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15644\,
            in1 => \N__16715\,
            in2 => \N__15780\,
            in3 => \N__17062\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__0_0_a2_1_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIG1RP4_13_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13781\,
            in1 => \N__14798\,
            in2 => \N__13448\,
            in3 => \N__15807\,
            lcout => \c0.un1_data_in_7__0_0_a2_1_a2_5_0\,
            ltout => \c0.un1_data_in_7__0_0_a2_1_a2_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIN2KLB_14_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17705\,
            in2 => \N__13445\,
            in3 => \N__17692\,
            lcout => \c0.tx2_transmit_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIN7VG_17_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13962\,
            in1 => \N__13731\,
            in2 => \N__14064\,
            in3 => \N__15526\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_7__3_0_a2_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIORVS2_43_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17035\,
            in1 => \N__15671\,
            in2 => \N__13787\,
            in3 => \N__13784\,
            lcout => \c0.un1_data_in_7__3_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__1_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13763\,
            lcout => \c0.d_4_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21869\,
            ce => \N__21589\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__6_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13709\,
            lcout => \c0.d_4_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21869\,
            ce => \N__21589\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIA0HJ_0_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13961\,
            in1 => \N__13629\,
            in2 => \_gnd_net_\,
            in3 => \N__13609\,
            lcout => \c0.N_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__0_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13685\,
            lcout => \c0.d_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21869\,
            ce => \N__21589\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__0_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13667\,
            lcout => \c0.d_4_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21869\,
            ce => \N__21589\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_0_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__18281\,
            in1 => \N__19541\,
            in2 => \N__13613\,
            in3 => \N__18911\,
            lcout => \c0.tx2_data_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__4_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13589\,
            lcout => \c0.d_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__21592\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__2_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13943\,
            lcout => \c0.d_4_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__21592\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__3_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13928\,
            lcout => \c0.d_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__21592\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__5_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13898\,
            lcout => \c0.d_4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__21592\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__5_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13871\,
            lcout => \c0.d_4_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__21592\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__1_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13846\,
            lcout => \c0.d_4_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__21592\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__1_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13823\,
            lcout => \c0.d_4_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__21592\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__3_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13808\,
            lcout => \c0.d_4_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21876\,
            ce => \N__21592\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_6_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__20928\,
            in1 => \N__18092\,
            in2 => \_gnd_net_\,
            in3 => \N__15461\,
            lcout => OPEN,
            ltout => \c0.tx2_data_1_iv_3_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_6_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__20410\,
            in1 => \_gnd_net_\,
            in2 => \N__13790\,
            in3 => \N__20340\,
            lcout => \c0.tx2_data_1_iv_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI1VL6_13_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17055\,
            in1 => \N__15760\,
            in2 => \_gnd_net_\,
            in3 => \N__16691\,
            lcout => \c0.N_132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIH9JJ_4_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14150\,
            in1 => \N__16049\,
            in2 => \_gnd_net_\,
            in3 => \N__19687\,
            lcout => \c0.N_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNII9QU3_14_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__14022\,
            in1 => \N__15551\,
            in2 => \_gnd_net_\,
            in3 => \N__16099\,
            lcout => \c0.d_4_RNII9QU3Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI675O1_33_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14151\,
            in1 => \N__15497\,
            in2 => \N__16277\,
            in3 => \N__16050\,
            lcout => \c0.un1_data_in_7__7_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_3_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010111111111"
        )
    port map (
            in0 => \N__18005\,
            in1 => \N__20612\,
            in2 => \N__20940\,
            in3 => \N__20409\,
            lcout => \c0.tx2_data_1_0_i_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_5_3_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__20932\,
            in1 => \N__14030\,
            in2 => \_gnd_net_\,
            in3 => \N__15660\,
            lcout => \c0.tx2_data_1_iv_4_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__4_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14093\,
            lcout => \c0.d_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21892\,
            ce => \N__21597\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__3_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14066\,
            lcout => \c0.data_in_frame_7_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21892\,
            ce => \N__21597\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_6_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111110111111"
        )
    port map (
            in0 => \N__20933\,
            in1 => \N__14023\,
            in2 => \N__17869\,
            in3 => \N__13970\,
            lcout => OPEN,
            ltout => \c0.tx2_data_1_iv_4_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_6_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111110000"
        )
    port map (
            in0 => \N__18449\,
            in1 => \N__17865\,
            in2 => \N__14456\,
            in3 => \N__20341\,
            lcout => \c0.tx2_data_1_iv_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__3_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14453\,
            lcout => \c0.d_4_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21892\,
            ce => \N__21597\,
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_7_1_0__m5_0_a2_0_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__19763\,
            in1 => \N__16346\,
            in2 => \N__14421\,
            in3 => \N__14341\,
            lcout => \c0.tx2.r_Tx_Data_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_0_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011000010"
        )
    port map (
            in0 => \N__16347\,
            in1 => \N__16381\,
            in2 => \N__16463\,
            in3 => \N__16438\,
            lcout => \c0.tx2.r_Bit_IndexZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21902\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_RNIMCBI_0_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14398\,
            in2 => \_gnd_net_\,
            in3 => \N__14340\,
            lcout => \c0.tx2.N_257\,
            ltout => \c0.tx2.N_257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_SM_Main_7_1_0__m5_0_o2_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__16457\,
            in1 => \N__16302\,
            in2 => \N__14303\,
            in3 => \N__16437\,
            lcout => \c0.tx2.N_261\,
            ltout => \c0.tx2.N_261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_2_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14294\,
            in2 => \N__14237\,
            in3 => \N__14232\,
            lcout => \c0.tx2.r_Bit_IndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21902\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14200\,
            in2 => \_gnd_net_\,
            in3 => \N__14186\,
            lcout => \c0.tx_transmitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21902\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_active_RNI6GJO_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14199\,
            in2 => \_gnd_net_\,
            in3 => \N__14185\,
            lcout => \c0.byte_transmit_counter15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_6_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100111111"
        )
    port map (
            in0 => \N__20600\,
            in1 => \N__14765\,
            in2 => \N__14756\,
            in3 => \N__20355\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21909\,
            ce => \N__20750\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_3_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__19312\,
            in1 => \N__14465\,
            in2 => \N__14735\,
            in3 => \N__19172\,
            lcout => \c0.tx_data_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_1_7_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__19313\,
            in1 => \N__19173\,
            in2 => \N__14693\,
            in3 => \N__15365\,
            lcout => \c0.tx_data_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_2_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__19170\,
            in1 => \N__17434\,
            in2 => \N__15257\,
            in3 => \N__19314\,
            lcout => OPEN,
            ltout => \c0.tx_data_RNO_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_2_2_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__17520\,
            in1 => \N__16782\,
            in2 => \N__14669\,
            in3 => \N__14582\,
            lcout => \c0.tx_data_1_0_i_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_4_2_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__19171\,
            in1 => \N__14653\,
            in2 => \N__14630\,
            in3 => \N__19311\,
            lcout => \c0.tx_data_RNO_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_RNIRD6P_0_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16781\,
            in2 => \_gnd_net_\,
            in3 => \N__17475\,
            lcout => \c0.N_201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_6__6_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15331\,
            in1 => \N__14974\,
            in2 => \_gnd_net_\,
            in3 => \N__14576\,
            lcout => \c0.data_out_6_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21917\,
            ce => \N__17292\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__3_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14546\,
            in1 => \N__14500\,
            in2 => \N__14912\,
            in3 => \N__15176\,
            lcout => \c0.data_out_7_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21917\,
            ce => \N__17292\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_1_3_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15142\,
            in1 => \N__15361\,
            in2 => \N__15330\,
            in3 => \N__15287\,
            lcout => OPEN,
            ltout => \c0.un105_newcrc_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_3_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15239\,
            in1 => \N__15209\,
            in2 => \N__15179\,
            in3 => \N__14940\,
            lcout => \c0.un105_newcrc_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_1_6_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__15159\,
            in1 => \N__15143\,
            in2 => \N__15110\,
            in3 => \N__14856\,
            lcout => \c0.un144_newcrc_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_6_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15061\,
            in1 => \N__15022\,
            in2 => \_gnd_net_\,
            in3 => \N__16515\,
            lcout => \c0.un144_newcrc_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_1_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14978\,
            in1 => \N__14960\,
            in2 => \N__14920\,
            in3 => \N__14861\,
            lcout => \c0.nextCRC16_3_0_a2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI22UN_24_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18649\,
            in1 => \N__20534\,
            in2 => \N__14816\,
            in3 => \N__16132\,
            lcout => \c0.un1_data_in_6__4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_6__RNIFRNC_4_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16619\,
            in1 => \N__15781\,
            in2 => \N__22271\,
            in3 => \N__16708\,
            lcout => \c0.un1_data_in_6__4_0_a2_5_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI9IAQ1_31_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18347\,
            in1 => \N__14807\,
            in2 => \N__14780\,
            in3 => \N__17917\,
            lcout => OPEN,
            ltout => \c0.wait_for_transmission4_12_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI7HDA4_24_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__15563\,
            in1 => \N__15638\,
            in2 => \N__15632\,
            in3 => \N__15629\,
            lcout => \c0.wait_for_transmission4_12_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_7__RNIBJH41_6_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16151\,
            in1 => \N__17995\,
            in2 => \N__19877\,
            in3 => \N__15605\,
            lcout => \c0.un1_data_in_7__6_0_a2_5_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_11_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__16620\,
            in1 => \N__16030\,
            in2 => \_gnd_net_\,
            in3 => \N__18253\,
            lcout => \c0.wait_for_transmission_RNOZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI4SA91_10_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16029\,
            in1 => \N__18252\,
            in2 => \N__16627\,
            in3 => \N__15490\,
            lcout => \c0.un1_data_in_6__7_0_a2_17_a2_4_1\,
            ltout => \c0.un1_data_in_6__7_0_a2_17_a2_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIV4MJ3_24_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16150\,
            in1 => \N__18572\,
            in2 => \N__15530\,
            in3 => \N__15862\,
            lcout => \c0.N_136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIJLQL_47_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17991\,
            in1 => \N__15383\,
            in2 => \N__15525\,
            in3 => \N__15452\,
            lcout => \c0.N_125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__6_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15479\,
            lcout => \c0.d_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21870\,
            ce => \N__21584\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__3_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15431\,
            lcout => \c0.d_4_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21870\,
            ce => \N__21584\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIQCTH_24_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20533\,
            in1 => \N__18178\,
            in2 => \N__18650\,
            in3 => \N__16124\,
            lcout => \c0.un1_data_in_6__7_0_a2_17_a2_4_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__3_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15851\,
            lcout => \c0.d_4_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21870\,
            ce => \N__21584\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIO7RC_28_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20588\,
            in1 => \N__18967\,
            in2 => \N__15898\,
            in3 => \N__15670\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__6_0_a2_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI15AH_12_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__17180\,
            in1 => \_gnd_net_\,
            in2 => \N__15833\,
            in3 => \N__18431\,
            lcout => \c0.un1_data_in_6__6_0_a2_0_a2_3\,
            ltout => \c0.un1_data_in_6__6_0_a2_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNITU3G2_19_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__15830\,
            in1 => \N__15732\,
            in2 => \N__15821\,
            in3 => \N__15810\,
            lcout => \c0.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIN4PC_27_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__16018\,
            in1 => \N__15761\,
            in2 => \N__19928\,
            in3 => \N__17800\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__5_0_a2_5_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI23VN_12_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18430\,
            in1 => \N__17179\,
            in2 => \N__15737\,
            in3 => \N__16125\,
            lcout => \c0.un1_data_in_6__5\,
            ltout => \c0.un1_data_in_6__5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIOEM13_24_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001001"
        )
    port map (
            in0 => \N__15733\,
            in1 => \N__15694\,
            in2 => \N__15683\,
            in3 => \N__18188\,
            lcout => \c0.g0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIH0UG_27_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__17799\,
            in1 => \N__15669\,
            in2 => \N__18746\,
            in3 => \N__17178\,
            lcout => \c0.un1_data_in_7__0_0_a2_1_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI21N6_11_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__15890\,
            in1 => \N__18209\,
            in2 => \_gnd_net_\,
            in3 => \N__17770\,
            lcout => \c0.d_4_RNI21N6Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIQ7PC_23_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18036\,
            in1 => \N__20532\,
            in2 => \N__20641\,
            in3 => \N__20158\,
            lcout => OPEN,
            ltout => \c0.un1_data_in_6__3_0_a2_5_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIRKQ41_10_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15983\,
            in1 => \N__16615\,
            in2 => \N__16034\,
            in3 => \N__16025\,
            lcout => \c0.un1_data_in_6__3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIPIKJ_39_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18248\,
            in1 => \N__15891\,
            in2 => \_gnd_net_\,
            in3 => \N__18211\,
            lcout => \c0.un1_data_in_6__3_0_a2_5_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__1_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15977\,
            lcout => \c0.d_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21884\,
            ce => \N__21590\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__7_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15947\,
            lcout => \c0.d_4_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21884\,
            ce => \N__21590\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__7_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18841\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_4_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21884\,
            ce => \N__21590\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__0_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15917\,
            lcout => \c0.d_4_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21884\,
            ce => \N__21590\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__5_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20002\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_4_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21884\,
            ce => \N__21590\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI6FQT_21_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20470\,
            in1 => \N__20430\,
            in2 => \N__22227\,
            in3 => \N__18492\,
            lcout => \c0.un1_data_in_7__7_0_a2_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__5_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16268\,
            lcout => \c0.d_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21893\,
            ce => \N__21593\,
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_9_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19713\,
            in1 => \N__20469\,
            in2 => \N__18371\,
            in3 => \N__16167\,
            lcout => \c0.wait_for_transmission_RNOZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__2_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16235\,
            lcout => \c0.d_4_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21893\,
            ce => \N__21593\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__4_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16208\,
            lcout => \c0.d_4_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21893\,
            ce => \N__21593\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_5__6_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19895\,
            lcout => \c0.d_4_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21893\,
            ce => \N__21593\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIABPL_18_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19712\,
            in1 => \N__20468\,
            in2 => \N__18370\,
            in3 => \N__16166\,
            lcout => \c0.N_124\,
            ltout => \c0.N_124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIPF9J2_37_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18680\,
            in1 => \N__18582\,
            in2 => \N__16136\,
            in3 => \N__16133\,
            lcout => \c0.d_4_RNIPF9J2Z0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__1_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16085\,
            lcout => \c0.d_4_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21903\,
            ce => \N__21596\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__0_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18765\,
            lcout => \c0.data_in_frame_6_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21903\,
            ce => \N__21596\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__2_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16745\,
            lcout => \c0.d_4_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21903\,
            ce => \N__21596\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__1_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18801\,
            lcout => \c0.data_in_frame_6_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21903\,
            ce => \N__21596\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__2_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16655\,
            lcout => \c0.d_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21903\,
            ce => \N__21596\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__0_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18738\,
            lcout => \c0.data_in_frame_7_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21903\,
            ce => \N__21596\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__RNO_0_7_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16567\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16523\,
            lcout => \c0.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_6_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__21413\,
            in1 => \N__21497\,
            in2 => \_gnd_net_\,
            in3 => \N__21324\,
            lcout => \c0.rx.r_Rx_Bytece_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_RNO_0_1_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16462\,
            in2 => \_gnd_net_\,
            in3 => \N__16439\,
            lcout => OPEN,
            ltout => \c0.tx2.N_258_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Bit_Index_1_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100110001000"
        )
    port map (
            in0 => \N__16382\,
            in1 => \N__16303\,
            in2 => \N__16370\,
            in3 => \N__16367\,
            lcout => \c0.tx2.r_Bit_IndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_3_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21918\,
            ce => \N__19030\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_6_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21918\,
            ce => \N__19030\,
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_3_6_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19077\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19287\,
            lcout => OPEN,
            ltout => \c0.N_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_data_RNO_0_6_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101011111"
        )
    port map (
            in0 => \N__16967\,
            in1 => \N__17357\,
            in2 => \N__16961\,
            in3 => \N__17503\,
            lcout => \c0.N_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_RNIA0ET3_2_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__19019\,
            in1 => \N__19423\,
            in2 => \N__19114\,
            in3 => \N__19286\,
            lcout => \c0.data_out_0__1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_RNI3M6P_3_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16931\,
            in2 => \_gnd_net_\,
            in3 => \N__16925\,
            lcout => OPEN,
            ltout => \c0.m2_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_RNIQP0V1_4_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__19040\,
            in1 => \N__18695\,
            in2 => \N__16919\,
            in3 => \N__17573\,
            lcout => \c0.N_129_mux\,
            ltout => \c0.N_129_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_RNI92KB2_2_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16916\,
            in3 => \N__19076\,
            lcout => \c0.N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__16807\,
            in1 => \N__17505\,
            in2 => \_gnd_net_\,
            in3 => \N__19319\,
            lcout => \c0.byte_transmit_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21926\,
            ce => \N__19034\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_4_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21926\,
            ce => \N__19034\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17504\,
            in2 => \_gnd_net_\,
            in3 => \N__19318\,
            lcout => \c0.byte_transmit_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21926\,
            ce => \N__19034\,
            sr => \_gnd_net_\
        );

    \c0.data_out_7__6_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17441\,
            in1 => \N__17433\,
            in2 => \N__17402\,
            in3 => \N__17393\,
            lcout => \c0.data_out_7_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21932\,
            ce => \N__17288\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_4_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111110111111"
        )
    port map (
            in0 => \N__20327\,
            in1 => \N__17192\,
            in2 => \N__17858\,
            in3 => \N__17138\,
            lcout => \c0.tx2_data_1_0_i_1_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_7_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101110111"
        )
    port map (
            in0 => \N__17102\,
            in1 => \N__17876\,
            in2 => \N__17093\,
            in3 => \N__20277\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21871\,
            ce => \N__20734\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_5_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__20845\,
            in1 => \N__17835\,
            in2 => \N__20326\,
            in3 => \N__17066\,
            lcout => OPEN,
            ltout => \c0.data_in_frame_1__m_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_5_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__17042\,
            in1 => \N__20275\,
            in2 => \N__16997\,
            in3 => \N__18985\,
            lcout => OPEN,
            ltout => \c0.tx2_data_1_iv_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_5_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__20276\,
            in1 => \N__16994\,
            in2 => \N__16985\,
            in3 => \N__20189\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21871\,
            ce => \N__20734\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_7_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17945\,
            in1 => \N__20270\,
            in2 => \N__17850\,
            in3 => \N__20844\,
            lcout => OPEN,
            ltout => \c0.data_in_frame_1__m_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_1_7_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__20274\,
            in1 => \N__18986\,
            in2 => \N__17921\,
            in3 => \N__17918\,
            lcout => \c0.tx2_data_1_iv_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNIJBBP_6_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__19480\,
            in1 => \N__19607\,
            in2 => \N__19648\,
            in3 => \N__19738\,
            lcout => \c0.N_205\,
            ltout => \c0.N_205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_3_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111101111111"
        )
    port map (
            in0 => \N__20846\,
            in1 => \N__17807\,
            in2 => \N__17780\,
            in3 => \N__17777\,
            lcout => \c0.tx2_data_1_iv_4_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNI25GA4_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__18011\,
            in1 => \N__18139\,
            in2 => \N__17743\,
            in3 => \N__17726\,
            lcout => OPEN,
            ltout => \c0.g1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i12_7_c_RNIP740G_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001000000"
        )
    port map (
            in0 => \N__17704\,
            in1 => \N__17693\,
            in2 => \N__17663\,
            in3 => \N__17653\,
            lcout => OPEN,
            ltout => \c0.i12_7_c_RNIP740G_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIM68GI_19_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17636\,
            in3 => \N__17633\,
            lcout => OPEN,
            ltout => \c0.g1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI9LFUV_43_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__17620\,
            in1 => \N__17609\,
            in2 => \N__17591\,
            in3 => \N__17588\,
            lcout => \c0.d_4_RNI9LFUVZ0Z_43\,
            ltout => \c0.d_4_RNI9LFUVZ0Z_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNI9PP5B1_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010101011"
        )
    port map (
            in0 => \N__19803\,
            in1 => \N__19849\,
            in2 => \N__18068\,
            in3 => \N__19825\,
            lcout => \c0.wait_for_transmission_RNI9PP5BZ0Z1\,
            ltout => \c0.wait_for_transmission_RNI9PP5BZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_0_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18065\,
            in3 => \N__19486\,
            lcout => \c0.byte_transmit_counter2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21877\,
            ce => 'H',
            sr => \N__20053\
        );

    \c0.byte_transmit_counter2_1_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19485\,
            in1 => \N__20859\,
            in2 => \_gnd_net_\,
            in3 => \N__20078\,
            lcout => \c0.byte_transmit_counter2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21877\,
            ce => 'H',
            sr => \N__20053\
        );

    \c0.byte_transmit_counter2_2_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__20860\,
            in1 => \N__20289\,
            in2 => \N__20087\,
            in3 => \N__19487\,
            lcout => \c0.byte_transmit_counter2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21877\,
            ce => 'H',
            sr => \N__20053\
        );

    \c0.d_4_RNIBUMH1_0_37_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18550\,
            in1 => \N__20159\,
            in2 => \N__18500\,
            in3 => \N__18050\,
            lcout => \c0.un1_data_in_6__1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNINGK21_0_21_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18322\,
            in1 => \N__18035\,
            in2 => \N__18280\,
            in3 => \N__20443\,
            lcout => \c0.g0_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNINGK21_21_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20442\,
            in1 => \N__18272\,
            in2 => \N__18040\,
            in3 => \N__18321\,
            lcout => \c0.N_126\,
            ltout => \c0.N_126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIBUMH1_37_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20160\,
            in1 => \N__18496\,
            in2 => \N__18014\,
            in3 => \N__18549\,
            lcout => \c0.un1_data_in_6__1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_6__RNI15IA_1_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18003\,
            in1 => \N__20528\,
            in2 => \_gnd_net_\,
            in3 => \N__18805\,
            lcout => \c0.un1_data_in_6__1_0_a2_4_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__7_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17960\,
            lcout => \c0.d_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21885\,
            ce => \N__21585\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_1__0_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18308\,
            lcout => \c0.d_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21885\,
            ce => \N__21585\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNISRG61_39_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18273\,
            in1 => \N__18241\,
            in2 => \N__22110\,
            in3 => \N__18210\,
            lcout => \c0.un1_data_in_6__2_0_a2_6_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIK7NH1_0_24_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18155\,
            in1 => \N__20506\,
            in2 => \N__18644\,
            in3 => \N__18177\,
            lcout => \c0.un1_data_in_6__2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI76N6_22_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20156\,
            in1 => \N__18482\,
            in2 => \_gnd_net_\,
            in3 => \N__18083\,
            lcout => \c0.N_107\,
            ltout => \c0.N_107_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIK7NH1_24_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__18154\,
            in1 => \N__18627\,
            in2 => \N__18146\,
            in3 => \N__20507\,
            lcout => \c0.un1_data_in_6__2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_2__6_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18122\,
            lcout => \c0.d_4_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21894\,
            ce => \N__21587\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIU6U8_22_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18084\,
            in1 => \N__18626\,
            in2 => \N__18495\,
            in3 => \N__20504\,
            lcout => \c0.d_4_RNIU6U8Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIU6U8_0_22_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20505\,
            in1 => \N__18486\,
            in2 => \N__18640\,
            in3 => \N__18085\,
            lcout => OPEN,
            ltout => \c0.d_4_RNIU6U8_0Z0Z_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.d_4_RNIMI4K_37_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18689\,
            in2 => \N__18683\,
            in3 => \N__20157\,
            lcout => \c0.d_4_RNIMI4KZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_3__0_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_4_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21894\,
            ce => \N__21587\,
            sr => \_gnd_net_\
        );

    \c0.wait_for_transmission_RNO_7_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__20161\,
            in1 => \N__18493\,
            in2 => \N__18589\,
            in3 => \N__18554\,
            lcout => \c0.un1_data_in_6__1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__4_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18521\,
            lcout => \c0.d_4_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21904\,
            ce => \N__21591\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_4_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__18455\,
            in1 => \N__18494\,
            in2 => \_gnd_net_\,
            in3 => \N__20919\,
            lcout => \c0.tx2_data_1_iv_5_1_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__4_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22263\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_frame_6_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21904\,
            ce => \N__21591\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_5_6_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__20920\,
            in1 => \N__18437\,
            in2 => \_gnd_net_\,
            in3 => \N__18369\,
            lcout => \c0.tx2_data_1_iv_4_1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__6_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19870\,
            lcout => \c0.data_in_frame_7_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21904\,
            ce => \N__21591\,
            sr => \_gnd_net_\
        );

    \c0.d_4_RNI09QE_46_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22017\,
            in1 => \N__18419\,
            in2 => \_gnd_net_\,
            in3 => \N__18368\,
            lcout => \c0.un1_data_in_7__2_0_a2_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_7__4_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21509\,
            lcout => \c0.data_in_7_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21911\,
            ce => \N__22161\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__2_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21526\,
            lcout => \c0.data_in_7_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21911\,
            ce => \N__22161\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__7_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20665\,
            lcout => \c0.data_in_4_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21911\,
            ce => \N__22161\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__7_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18827\,
            lcout => \c0.data_in_7_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21911\,
            ce => \N__22161\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__1_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22069\,
            lcout => \c0.data_in_6_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21911\,
            ce => \N__22161\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__0_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18742\,
            lcout => \c0.data_in_6_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21911\,
            ce => \N__22161\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__0_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21071\,
            lcout => \c0.data_in_7_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21911\,
            ce => \N__22161\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__4_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22270\,
            lcout => \c0.data_in_5_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21911\,
            ce => \N__22161\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21919\,
            ce => \N__19029\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_2_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__19113\,
            in1 => \N__19430\,
            in2 => \_gnd_net_\,
            in3 => \N__19320\,
            lcout => \c0.byte_transmit_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21919\,
            ce => \N__19029\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_7_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \c0.byte_transmit_counterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21919\,
            ce => \N__19029\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__5_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19927\,
            lcout => \c0.data_in_frame_6_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21927\,
            ce => \N__21598\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_3_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21059\,
            in1 => \N__21039\,
            in2 => \_gnd_net_\,
            in3 => \N__20082\,
            lcout => \c0.byte_transmit_counter2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21878\,
            ce => 'H',
            sr => \N__20046\
        );

    \c0.tx2_data_RNO_2_4_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__20388\,
            in1 => \N__19676\,
            in2 => \N__18998\,
            in3 => \N__20279\,
            lcout => \c0.tx2_data_1_iv_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNIJFIT_0_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20831\,
            in1 => \N__19482\,
            in2 => \_gnd_net_\,
            in3 => \N__18873\,
            lcout => \c0.N_207\,
            ltout => \c0.N_207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_4_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101111111"
        )
    port map (
            in0 => \N__21944\,
            in1 => \N__20278\,
            in2 => \N__18971\,
            in3 => \N__18968\,
            lcout => \c0.tx2_data_1_0_i_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNIBNLC_7_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__21032\,
            in1 => \N__19666\,
            in2 => \_gnd_net_\,
            in3 => \N__21005\,
            lcout => \c0.m2_e_0_2\,
            ltout => \c0.m2_e_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNIK84L_6_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19630\,
            in2 => \N__18932\,
            in3 => \N__19599\,
            lcout => \c0.N_71_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_transmit_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000111001"
        )
    port map (
            in0 => \N__19850\,
            in1 => \N__19826\,
            in2 => \N__19811\,
            in3 => \N__19769\,
            lcout => \c0.tx2_transmitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNIJBBP_0_6_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__19481\,
            in1 => \N__19739\,
            in2 => \N__19649\,
            in3 => \N__19600\,
            lcout => \c0.N_203\,
            ltout => \c0.N_203_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_3_4_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111101111111"
        )
    port map (
            in0 => \N__20832\,
            in1 => \N__19727\,
            in2 => \N__19697\,
            in3 => \N__19694\,
            lcout => \c0.tx2_data_1_iv_5_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNO_1_7_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20858\,
            in1 => \N__21009\,
            in2 => \N__20325\,
            in3 => \N__21040\,
            lcout => OPEN,
            ltout => \c0.un1_m4_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_7_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__19655\,
            in1 => \N__19667\,
            in2 => \N__19670\,
            in3 => \N__20086\,
            lcout => \c0.byte_transmit_counter2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21895\,
            ce => 'H',
            sr => \N__20054\
        );

    \c0.byte_transmit_counter2_RNO_0_7_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19484\,
            in1 => \N__19637\,
            in2 => \_gnd_net_\,
            in3 => \N__19604\,
            lcout => \c0.un1_m4_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_6_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__20983\,
            in1 => \N__19606\,
            in2 => \N__19647\,
            in3 => \N__20085\,
            lcout => \c0.byte_transmit_counter2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21895\,
            ce => 'H',
            sr => \N__20054\
        );

    \c0.byte_transmit_counter2_5_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__19605\,
            in1 => \_gnd_net_\,
            in2 => \N__20984\,
            in3 => \N__20084\,
            lcout => \c0.byte_transmit_counter2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21895\,
            ce => 'H',
            sr => \N__20054\
        );

    \c0.byte_transmit_counter2_RNI0CLC_0_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__19483\,
            in1 => \_gnd_net_\,
            in2 => \N__20324\,
            in3 => \N__20843\,
            lcout => \c0.un1_byte_transmit_counter2_1_ac0_3_out\,
            ltout => \c0.un1_byte_transmit_counter2_1_ac0_3_out_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_4_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__21041\,
            in1 => \N__21010\,
            in2 => \N__20090\,
            in3 => \N__20083\,
            lcout => \c0.byte_transmit_counter2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21895\,
            ce => 'H',
            sr => \N__20054\
        );

    \c0.data_in_4__5_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19978\,
            lcout => \c0.data_in_4_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21905\,
            ce => \N__22160\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__5_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19914\,
            lcout => \c0.data_in_5_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21905\,
            ce => \N__22160\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__5_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19963\,
            lcout => \c0.data_in_6_Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21905\,
            ce => \N__22160\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__2_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22018\,
            lcout => \c0.data_in_6_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21905\,
            ce => \N__22160\,
            sr => \_gnd_net_\
        );

    \c0.data_in_4__6_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19888\,
            lcout => \c0.data_in_4_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21905\,
            ce => \N__22160\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__6_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20583\,
            lcout => \c0.data_in_5_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21905\,
            ce => \N__22160\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__6_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19869\,
            lcout => \c0.data_in_6_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21905\,
            ce => \N__22160\,
            sr => \_gnd_net_\
        );

    \c0.data_in_7__6_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20108\,
            lcout => \c0.data_in_7_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21905\,
            ce => \N__22160\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__3_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20642\,
            lcout => \c0.data_in_frame_6_Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21912\,
            ce => \N__21588\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_0_6_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101101111111"
        )
    port map (
            in0 => \N__20923\,
            in1 => \N__20390\,
            in2 => \N__20564\,
            in3 => \N__20515\,
            lcout => \c0.tx2_data_1_0_i_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__6_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20584\,
            lcout => \c0.data_in_frame_6_Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21912\,
            ce => \N__21588\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_4__6_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20545\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.d_4_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21912\,
            ce => \N__21588\,
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_4_5_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101110111"
        )
    port map (
            in0 => \N__20389\,
            in1 => \N__20474\,
            in2 => \N__20450\,
            in3 => \N__20922\,
            lcout => OPEN,
            ltout => \c0.tx2_data_1_iv_5_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_2_5_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111110000"
        )
    port map (
            in0 => \N__20126\,
            in1 => \N__20391\,
            in2 => \N__20360\,
            in3 => \N__20328\,
            lcout => \c0.tx2_data_1_iv_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2_data_RNO_5_5_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__20177\,
            in1 => \N__20921\,
            in2 => \_gnd_net_\,
            in3 => \N__20168\,
            lcout => \c0.tx2_data_1_iv_5_1_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_6_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__21245\,
            in1 => \N__20120\,
            in2 => \N__20107\,
            in3 => \N__21144\,
            lcout => \c0.rx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21920\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_2_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__21142\,
            in1 => \N__21536\,
            in2 => \N__21527\,
            in3 => \N__21243\,
            lcout => \c0.rx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21920\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_4_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__21326\,
            in1 => \_gnd_net_\,
            in2 => \N__21412\,
            in3 => \N__21496\,
            lcout => OPEN,
            ltout => \c0.rx.r_Rx_Bytece_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_4_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__21143\,
            in1 => \N__21508\,
            in2 => \N__21512\,
            in3 => \N__21244\,
            lcout => \c0.rx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21920\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_RNO_0_0_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__21495\,
            in1 => \N__21403\,
            in2 => \_gnd_net_\,
            in3 => \N__21325\,
            lcout => OPEN,
            ltout => \c0.rx.r_Rx_Bytece_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_0_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__21242\,
            in1 => \N__21070\,
            in2 => \N__21149\,
            in3 => \N__21141\,
            lcout => \c0.rx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21920\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter2_RNI5P3L_4_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21058\,
            in1 => \N__21033\,
            in2 => \_gnd_net_\,
            in3 => \N__21011\,
            lcout => \c0.un1_byte_transmit_counter2_1_ac0_7_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx2.r_Tx_Data_4_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__20969\,
            in1 => \N__20963\,
            in2 => \N__20957\,
            in3 => \N__20878\,
            lcout => \c0.tx2.r_Tx_DataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21896\,
            ce => \N__20733\,
            sr => \_gnd_net_\
        );

    \c0.data_in_5__7_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22190\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.data_in_5_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21913\,
            ce => \N__22162\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__4_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21975\,
            lcout => \c0.data_in_6_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21921\,
            ce => \N__22163\,
            sr => \_gnd_net_\
        );

    \c0.data_in_6__7_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22234\,
            lcout => \c0.data_in_6_Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21921\,
            ce => \N__22163\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_6__2_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22111\,
            lcout => \c0.data_in_frame_6_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21922\,
            ce => \N__21581\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__1_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22073\,
            lcout => \c0.data_in_frame_7_Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21928\,
            ce => \N__21582\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__2_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22022\,
            lcout => \c0.data_in_frame_7_Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21928\,
            ce => \N__21582\,
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_7__4_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21976\,
            lcout => \c0.data_in_frame_7_Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21928\,
            ce => \N__21582\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
