// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 12 2019 13:57:57

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    inout PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    inout PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    inout PIN_1;
    output LED;
    input CLK;

    wire N__37526;
    wire N__37525;
    wire N__37524;
    wire N__37517;
    wire N__37516;
    wire N__37515;
    wire N__37508;
    wire N__37507;
    wire N__37506;
    wire N__37499;
    wire N__37498;
    wire N__37497;
    wire N__37490;
    wire N__37489;
    wire N__37488;
    wire N__37481;
    wire N__37480;
    wire N__37479;
    wire N__37462;
    wire N__37461;
    wire N__37456;
    wire N__37453;
    wire N__37452;
    wire N__37449;
    wire N__37446;
    wire N__37441;
    wire N__37438;
    wire N__37437;
    wire N__37432;
    wire N__37429;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37417;
    wire N__37414;
    wire N__37413;
    wire N__37410;
    wire N__37405;
    wire N__37402;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37390;
    wire N__37387;
    wire N__37384;
    wire N__37383;
    wire N__37378;
    wire N__37375;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37351;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37339;
    wire N__37338;
    wire N__37335;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37291;
    wire N__37290;
    wire N__37289;
    wire N__37286;
    wire N__37285;
    wire N__37282;
    wire N__37281;
    wire N__37280;
    wire N__37279;
    wire N__37278;
    wire N__37277;
    wire N__37276;
    wire N__37275;
    wire N__37274;
    wire N__37273;
    wire N__37272;
    wire N__37271;
    wire N__37270;
    wire N__37269;
    wire N__37268;
    wire N__37267;
    wire N__37266;
    wire N__37265;
    wire N__37262;
    wire N__37261;
    wire N__37258;
    wire N__37251;
    wire N__37250;
    wire N__37243;
    wire N__37232;
    wire N__37231;
    wire N__37230;
    wire N__37229;
    wire N__37228;
    wire N__37227;
    wire N__37226;
    wire N__37223;
    wire N__37222;
    wire N__37219;
    wire N__37218;
    wire N__37215;
    wire N__37214;
    wire N__37213;
    wire N__37212;
    wire N__37209;
    wire N__37208;
    wire N__37207;
    wire N__37204;
    wire N__37203;
    wire N__37202;
    wire N__37201;
    wire N__37200;
    wire N__37199;
    wire N__37196;
    wire N__37195;
    wire N__37194;
    wire N__37191;
    wire N__37190;
    wire N__37189;
    wire N__37188;
    wire N__37187;
    wire N__37186;
    wire N__37185;
    wire N__37184;
    wire N__37181;
    wire N__37176;
    wire N__37171;
    wire N__37168;
    wire N__37167;
    wire N__37166;
    wire N__37165;
    wire N__37164;
    wire N__37163;
    wire N__37162;
    wire N__37161;
    wire N__37158;
    wire N__37155;
    wire N__37154;
    wire N__37153;
    wire N__37152;
    wire N__37151;
    wire N__37150;
    wire N__37149;
    wire N__37148;
    wire N__37147;
    wire N__37146;
    wire N__37145;
    wire N__37144;
    wire N__37143;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37132;
    wire N__37129;
    wire N__37128;
    wire N__37127;
    wire N__37126;
    wire N__37125;
    wire N__37124;
    wire N__37123;
    wire N__37120;
    wire N__37117;
    wire N__37116;
    wire N__37111;
    wire N__37106;
    wire N__37099;
    wire N__37090;
    wire N__37089;
    wire N__37088;
    wire N__37087;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37079;
    wire N__37074;
    wire N__37071;
    wire N__37070;
    wire N__37069;
    wire N__37068;
    wire N__37061;
    wire N__37060;
    wire N__37059;
    wire N__37058;
    wire N__37055;
    wire N__37054;
    wire N__37053;
    wire N__37050;
    wire N__37045;
    wire N__37042;
    wire N__37033;
    wire N__37026;
    wire N__37021;
    wire N__37010;
    wire N__37009;
    wire N__37008;
    wire N__37007;
    wire N__37006;
    wire N__37005;
    wire N__37004;
    wire N__37003;
    wire N__37002;
    wire N__37001;
    wire N__37000;
    wire N__36999;
    wire N__36998;
    wire N__36997;
    wire N__36996;
    wire N__36993;
    wire N__36992;
    wire N__36991;
    wire N__36990;
    wire N__36989;
    wire N__36984;
    wire N__36977;
    wire N__36966;
    wire N__36957;
    wire N__36956;
    wire N__36955;
    wire N__36954;
    wire N__36953;
    wire N__36952;
    wire N__36951;
    wire N__36950;
    wire N__36945;
    wire N__36938;
    wire N__36937;
    wire N__36934;
    wire N__36927;
    wire N__36922;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36902;
    wire N__36895;
    wire N__36894;
    wire N__36893;
    wire N__36890;
    wire N__36889;
    wire N__36888;
    wire N__36885;
    wire N__36882;
    wire N__36881;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36865;
    wire N__36862;
    wire N__36857;
    wire N__36854;
    wire N__36849;
    wire N__36848;
    wire N__36847;
    wire N__36846;
    wire N__36845;
    wire N__36842;
    wire N__36837;
    wire N__36826;
    wire N__36823;
    wire N__36816;
    wire N__36815;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36807;
    wire N__36806;
    wire N__36805;
    wire N__36804;
    wire N__36803;
    wire N__36802;
    wire N__36799;
    wire N__36798;
    wire N__36795;
    wire N__36792;
    wire N__36791;
    wire N__36788;
    wire N__36787;
    wire N__36786;
    wire N__36785;
    wire N__36782;
    wire N__36775;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36757;
    wire N__36752;
    wire N__36745;
    wire N__36742;
    wire N__36739;
    wire N__36734;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36716;
    wire N__36711;
    wire N__36706;
    wire N__36705;
    wire N__36704;
    wire N__36699;
    wire N__36692;
    wire N__36691;
    wire N__36686;
    wire N__36681;
    wire N__36678;
    wire N__36673;
    wire N__36666;
    wire N__36663;
    wire N__36654;
    wire N__36651;
    wire N__36650;
    wire N__36649;
    wire N__36640;
    wire N__36639;
    wire N__36638;
    wire N__36637;
    wire N__36636;
    wire N__36635;
    wire N__36630;
    wire N__36627;
    wire N__36622;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36608;
    wire N__36607;
    wire N__36606;
    wire N__36605;
    wire N__36604;
    wire N__36599;
    wire N__36592;
    wire N__36587;
    wire N__36584;
    wire N__36579;
    wire N__36574;
    wire N__36567;
    wire N__36562;
    wire N__36557;
    wire N__36542;
    wire N__36537;
    wire N__36532;
    wire N__36529;
    wire N__36524;
    wire N__36513;
    wire N__36510;
    wire N__36509;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36501;
    wire N__36500;
    wire N__36497;
    wire N__36496;
    wire N__36495;
    wire N__36494;
    wire N__36491;
    wire N__36486;
    wire N__36483;
    wire N__36482;
    wire N__36479;
    wire N__36466;
    wire N__36455;
    wire N__36446;
    wire N__36441;
    wire N__36438;
    wire N__36437;
    wire N__36430;
    wire N__36425;
    wire N__36416;
    wire N__36413;
    wire N__36402;
    wire N__36399;
    wire N__36392;
    wire N__36387;
    wire N__36380;
    wire N__36377;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36357;
    wire N__36350;
    wire N__36331;
    wire N__36330;
    wire N__36329;
    wire N__36328;
    wire N__36327;
    wire N__36324;
    wire N__36323;
    wire N__36322;
    wire N__36321;
    wire N__36320;
    wire N__36319;
    wire N__36316;
    wire N__36315;
    wire N__36314;
    wire N__36313;
    wire N__36312;
    wire N__36311;
    wire N__36310;
    wire N__36309;
    wire N__36302;
    wire N__36299;
    wire N__36294;
    wire N__36293;
    wire N__36292;
    wire N__36291;
    wire N__36290;
    wire N__36289;
    wire N__36282;
    wire N__36277;
    wire N__36274;
    wire N__36273;
    wire N__36272;
    wire N__36271;
    wire N__36270;
    wire N__36267;
    wire N__36266;
    wire N__36265;
    wire N__36264;
    wire N__36263;
    wire N__36262;
    wire N__36261;
    wire N__36258;
    wire N__36257;
    wire N__36256;
    wire N__36255;
    wire N__36254;
    wire N__36253;
    wire N__36252;
    wire N__36251;
    wire N__36244;
    wire N__36241;
    wire N__36236;
    wire N__36235;
    wire N__36232;
    wire N__36231;
    wire N__36230;
    wire N__36229;
    wire N__36228;
    wire N__36227;
    wire N__36226;
    wire N__36225;
    wire N__36224;
    wire N__36223;
    wire N__36222;
    wire N__36219;
    wire N__36218;
    wire N__36217;
    wire N__36216;
    wire N__36215;
    wire N__36212;
    wire N__36209;
    wire N__36208;
    wire N__36207;
    wire N__36206;
    wire N__36205;
    wire N__36204;
    wire N__36203;
    wire N__36202;
    wire N__36201;
    wire N__36200;
    wire N__36199;
    wire N__36198;
    wire N__36197;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36193;
    wire N__36190;
    wire N__36183;
    wire N__36176;
    wire N__36175;
    wire N__36174;
    wire N__36173;
    wire N__36172;
    wire N__36171;
    wire N__36170;
    wire N__36169;
    wire N__36168;
    wire N__36167;
    wire N__36164;
    wire N__36163;
    wire N__36162;
    wire N__36161;
    wire N__36160;
    wire N__36159;
    wire N__36154;
    wire N__36147;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36130;
    wire N__36123;
    wire N__36120;
    wire N__36113;
    wire N__36102;
    wire N__36101;
    wire N__36096;
    wire N__36091;
    wire N__36088;
    wire N__36087;
    wire N__36086;
    wire N__36085;
    wire N__36084;
    wire N__36083;
    wire N__36082;
    wire N__36081;
    wire N__36076;
    wire N__36073;
    wire N__36064;
    wire N__36063;
    wire N__36062;
    wire N__36061;
    wire N__36060;
    wire N__36059;
    wire N__36058;
    wire N__36057;
    wire N__36050;
    wire N__36045;
    wire N__36042;
    wire N__36041;
    wire N__36040;
    wire N__36039;
    wire N__36038;
    wire N__36037;
    wire N__36036;
    wire N__36035;
    wire N__36034;
    wire N__36033;
    wire N__36032;
    wire N__36031;
    wire N__36030;
    wire N__36027;
    wire N__36026;
    wire N__36025;
    wire N__36024;
    wire N__36019;
    wire N__36018;
    wire N__36017;
    wire N__36014;
    wire N__36013;
    wire N__36012;
    wire N__36011;
    wire N__36010;
    wire N__36007;
    wire N__36006;
    wire N__36005;
    wire N__36000;
    wire N__35997;
    wire N__35996;
    wire N__35993;
    wire N__35992;
    wire N__35991;
    wire N__35990;
    wire N__35989;
    wire N__35988;
    wire N__35987;
    wire N__35986;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35970;
    wire N__35967;
    wire N__35966;
    wire N__35965;
    wire N__35964;
    wire N__35961;
    wire N__35956;
    wire N__35951;
    wire N__35944;
    wire N__35939;
    wire N__35930;
    wire N__35925;
    wire N__35922;
    wire N__35917;
    wire N__35904;
    wire N__35901;
    wire N__35896;
    wire N__35887;
    wire N__35878;
    wire N__35875;
    wire N__35870;
    wire N__35865;
    wire N__35864;
    wire N__35863;
    wire N__35862;
    wire N__35861;
    wire N__35860;
    wire N__35859;
    wire N__35858;
    wire N__35857;
    wire N__35846;
    wire N__35839;
    wire N__35838;
    wire N__35837;
    wire N__35832;
    wire N__35825;
    wire N__35818;
    wire N__35809;
    wire N__35800;
    wire N__35797;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35781;
    wire N__35772;
    wire N__35769;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35755;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35730;
    wire N__35727;
    wire N__35722;
    wire N__35717;
    wire N__35706;
    wire N__35701;
    wire N__35698;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35674;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35653;
    wire N__35652;
    wire N__35651;
    wire N__35650;
    wire N__35649;
    wire N__35648;
    wire N__35647;
    wire N__35646;
    wire N__35645;
    wire N__35644;
    wire N__35643;
    wire N__35642;
    wire N__35641;
    wire N__35640;
    wire N__35639;
    wire N__35636;
    wire N__35633;
    wire N__35628;
    wire N__35625;
    wire N__35620;
    wire N__35615;
    wire N__35606;
    wire N__35603;
    wire N__35600;
    wire N__35595;
    wire N__35590;
    wire N__35583;
    wire N__35574;
    wire N__35571;
    wire N__35566;
    wire N__35559;
    wire N__35556;
    wire N__35549;
    wire N__35546;
    wire N__35543;
    wire N__35536;
    wire N__35529;
    wire N__35524;
    wire N__35517;
    wire N__35512;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35494;
    wire N__35481;
    wire N__35476;
    wire N__35469;
    wire N__35440;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35410;
    wire N__35409;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35405;
    wire N__35404;
    wire N__35403;
    wire N__35402;
    wire N__35401;
    wire N__35400;
    wire N__35399;
    wire N__35398;
    wire N__35397;
    wire N__35396;
    wire N__35395;
    wire N__35394;
    wire N__35393;
    wire N__35392;
    wire N__35391;
    wire N__35390;
    wire N__35389;
    wire N__35388;
    wire N__35387;
    wire N__35386;
    wire N__35385;
    wire N__35384;
    wire N__35383;
    wire N__35382;
    wire N__35381;
    wire N__35380;
    wire N__35379;
    wire N__35378;
    wire N__35377;
    wire N__35376;
    wire N__35375;
    wire N__35374;
    wire N__35373;
    wire N__35372;
    wire N__35371;
    wire N__35370;
    wire N__35369;
    wire N__35368;
    wire N__35367;
    wire N__35366;
    wire N__35365;
    wire N__35364;
    wire N__35363;
    wire N__35362;
    wire N__35361;
    wire N__35360;
    wire N__35359;
    wire N__35358;
    wire N__35357;
    wire N__35356;
    wire N__35355;
    wire N__35354;
    wire N__35353;
    wire N__35352;
    wire N__35351;
    wire N__35350;
    wire N__35349;
    wire N__35348;
    wire N__35347;
    wire N__35346;
    wire N__35345;
    wire N__35344;
    wire N__35343;
    wire N__35342;
    wire N__35341;
    wire N__35340;
    wire N__35339;
    wire N__35338;
    wire N__35337;
    wire N__35336;
    wire N__35335;
    wire N__35334;
    wire N__35333;
    wire N__35332;
    wire N__35331;
    wire N__35330;
    wire N__35329;
    wire N__35328;
    wire N__35327;
    wire N__35326;
    wire N__35325;
    wire N__35324;
    wire N__35323;
    wire N__35322;
    wire N__35321;
    wire N__35320;
    wire N__35319;
    wire N__35318;
    wire N__35317;
    wire N__35316;
    wire N__35315;
    wire N__35314;
    wire N__35313;
    wire N__35312;
    wire N__35311;
    wire N__35310;
    wire N__35309;
    wire N__35308;
    wire N__35307;
    wire N__35306;
    wire N__35305;
    wire N__35304;
    wire N__35303;
    wire N__35302;
    wire N__35301;
    wire N__35300;
    wire N__35299;
    wire N__35298;
    wire N__35297;
    wire N__35296;
    wire N__35295;
    wire N__35294;
    wire N__35293;
    wire N__35292;
    wire N__35291;
    wire N__35290;
    wire N__35289;
    wire N__35288;
    wire N__35287;
    wire N__35286;
    wire N__35285;
    wire N__35284;
    wire N__35283;
    wire N__35282;
    wire N__35281;
    wire N__35280;
    wire N__35279;
    wire N__35278;
    wire N__35277;
    wire N__35276;
    wire N__35275;
    wire N__35274;
    wire N__35273;
    wire N__35272;
    wire N__35271;
    wire N__35270;
    wire N__35269;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34843;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34831;
    wire N__34830;
    wire N__34829;
    wire N__34828;
    wire N__34827;
    wire N__34822;
    wire N__34821;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34813;
    wire N__34812;
    wire N__34811;
    wire N__34808;
    wire N__34807;
    wire N__34806;
    wire N__34805;
    wire N__34804;
    wire N__34801;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34763;
    wire N__34762;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34748;
    wire N__34747;
    wire N__34744;
    wire N__34735;
    wire N__34730;
    wire N__34727;
    wire N__34722;
    wire N__34717;
    wire N__34714;
    wire N__34707;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34651;
    wire N__34648;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34617;
    wire N__34614;
    wire N__34613;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34598;
    wire N__34591;
    wire N__34588;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34576;
    wire N__34573;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34557;
    wire N__34554;
    wire N__34553;
    wire N__34552;
    wire N__34551;
    wire N__34550;
    wire N__34549;
    wire N__34548;
    wire N__34547;
    wire N__34546;
    wire N__34545;
    wire N__34544;
    wire N__34543;
    wire N__34542;
    wire N__34541;
    wire N__34540;
    wire N__34539;
    wire N__34538;
    wire N__34537;
    wire N__34536;
    wire N__34535;
    wire N__34534;
    wire N__34533;
    wire N__34532;
    wire N__34531;
    wire N__34530;
    wire N__34529;
    wire N__34528;
    wire N__34527;
    wire N__34526;
    wire N__34525;
    wire N__34524;
    wire N__34523;
    wire N__34514;
    wire N__34509;
    wire N__34506;
    wire N__34505;
    wire N__34502;
    wire N__34501;
    wire N__34500;
    wire N__34499;
    wire N__34498;
    wire N__34497;
    wire N__34496;
    wire N__34495;
    wire N__34494;
    wire N__34493;
    wire N__34492;
    wire N__34491;
    wire N__34490;
    wire N__34487;
    wire N__34482;
    wire N__34479;
    wire N__34478;
    wire N__34475;
    wire N__34474;
    wire N__34473;
    wire N__34468;
    wire N__34467;
    wire N__34466;
    wire N__34465;
    wire N__34464;
    wire N__34461;
    wire N__34460;
    wire N__34459;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34451;
    wire N__34450;
    wire N__34449;
    wire N__34448;
    wire N__34447;
    wire N__34446;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34428;
    wire N__34427;
    wire N__34426;
    wire N__34425;
    wire N__34424;
    wire N__34423;
    wire N__34422;
    wire N__34421;
    wire N__34418;
    wire N__34417;
    wire N__34416;
    wire N__34415;
    wire N__34414;
    wire N__34413;
    wire N__34412;
    wire N__34409;
    wire N__34408;
    wire N__34407;
    wire N__34406;
    wire N__34403;
    wire N__34398;
    wire N__34391;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34379;
    wire N__34378;
    wire N__34375;
    wire N__34368;
    wire N__34367;
    wire N__34364;
    wire N__34363;
    wire N__34362;
    wire N__34361;
    wire N__34354;
    wire N__34349;
    wire N__34342;
    wire N__34337;
    wire N__34334;
    wire N__34329;
    wire N__34324;
    wire N__34321;
    wire N__34320;
    wire N__34319;
    wire N__34310;
    wire N__34307;
    wire N__34302;
    wire N__34297;
    wire N__34296;
    wire N__34295;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34287;
    wire N__34286;
    wire N__34285;
    wire N__34284;
    wire N__34283;
    wire N__34282;
    wire N__34281;
    wire N__34280;
    wire N__34279;
    wire N__34278;
    wire N__34273;
    wire N__34268;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34252;
    wire N__34247;
    wire N__34232;
    wire N__34221;
    wire N__34220;
    wire N__34219;
    wire N__34218;
    wire N__34217;
    wire N__34216;
    wire N__34215;
    wire N__34212;
    wire N__34203;
    wire N__34196;
    wire N__34189;
    wire N__34186;
    wire N__34181;
    wire N__34172;
    wire N__34169;
    wire N__34168;
    wire N__34167;
    wire N__34166;
    wire N__34163;
    wire N__34158;
    wire N__34153;
    wire N__34152;
    wire N__34151;
    wire N__34148;
    wire N__34147;
    wire N__34142;
    wire N__34141;
    wire N__34140;
    wire N__34139;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34127;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34103;
    wire N__34100;
    wire N__34095;
    wire N__34090;
    wire N__34083;
    wire N__34082;
    wire N__34081;
    wire N__34078;
    wire N__34077;
    wire N__34076;
    wire N__34075;
    wire N__34074;
    wire N__34073;
    wire N__34068;
    wire N__34061;
    wire N__34058;
    wire N__34051;
    wire N__34038;
    wire N__34037;
    wire N__34036;
    wire N__34035;
    wire N__34032;
    wire N__34031;
    wire N__34030;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34016;
    wire N__34015;
    wire N__34014;
    wire N__34013;
    wire N__34012;
    wire N__34011;
    wire N__34010;
    wire N__34009;
    wire N__34000;
    wire N__33993;
    wire N__33988;
    wire N__33983;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33941;
    wire N__33934;
    wire N__33931;
    wire N__33926;
    wire N__33923;
    wire N__33922;
    wire N__33921;
    wire N__33920;
    wire N__33919;
    wire N__33918;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33886;
    wire N__33885;
    wire N__33884;
    wire N__33883;
    wire N__33882;
    wire N__33881;
    wire N__33880;
    wire N__33879;
    wire N__33878;
    wire N__33877;
    wire N__33876;
    wire N__33875;
    wire N__33874;
    wire N__33873;
    wire N__33872;
    wire N__33865;
    wire N__33862;
    wire N__33855;
    wire N__33852;
    wire N__33847;
    wire N__33842;
    wire N__33837;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33817;
    wire N__33812;
    wire N__33805;
    wire N__33794;
    wire N__33787;
    wire N__33784;
    wire N__33775;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33753;
    wire N__33746;
    wire N__33739;
    wire N__33734;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33714;
    wire N__33701;
    wire N__33692;
    wire N__33683;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33651;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33634;
    wire N__33631;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33619;
    wire N__33616;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33558;
    wire N__33555;
    wire N__33552;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33535;
    wire N__33532;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33518;
    wire N__33513;
    wire N__33510;
    wire N__33505;
    wire N__33502;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33490;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33478;
    wire N__33477;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33455;
    wire N__33454;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33433;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33403;
    wire N__33402;
    wire N__33399;
    wire N__33398;
    wire N__33395;
    wire N__33394;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33368;
    wire N__33361;
    wire N__33360;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33328;
    wire N__33325;
    wire N__33316;
    wire N__33315;
    wire N__33312;
    wire N__33311;
    wire N__33310;
    wire N__33309;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33299;
    wire N__33298;
    wire N__33295;
    wire N__33294;
    wire N__33291;
    wire N__33290;
    wire N__33289;
    wire N__33288;
    wire N__33287;
    wire N__33286;
    wire N__33285;
    wire N__33282;
    wire N__33277;
    wire N__33276;
    wire N__33275;
    wire N__33274;
    wire N__33273;
    wire N__33272;
    wire N__33271;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33247;
    wire N__33246;
    wire N__33241;
    wire N__33238;
    wire N__33237;
    wire N__33236;
    wire N__33233;
    wire N__33228;
    wire N__33223;
    wire N__33222;
    wire N__33221;
    wire N__33218;
    wire N__33213;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33202;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33190;
    wire N__33187;
    wire N__33186;
    wire N__33185;
    wire N__33184;
    wire N__33183;
    wire N__33182;
    wire N__33181;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33139;
    wire N__33138;
    wire N__33135;
    wire N__33128;
    wire N__33123;
    wire N__33118;
    wire N__33117;
    wire N__33116;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33104;
    wire N__33101;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33079;
    wire N__33076;
    wire N__33067;
    wire N__33062;
    wire N__33053;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33033;
    wire N__33024;
    wire N__33017;
    wire N__33014;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32994;
    wire N__32991;
    wire N__32990;
    wire N__32987;
    wire N__32986;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32972;
    wire N__32965;
    wire N__32964;
    wire N__32961;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32950;
    wire N__32947;
    wire N__32942;
    wire N__32939;
    wire N__32938;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32924;
    wire N__32921;
    wire N__32914;
    wire N__32913;
    wire N__32910;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32893;
    wire N__32890;
    wire N__32889;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32875;
    wire N__32872;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32854;
    wire N__32853;
    wire N__32852;
    wire N__32849;
    wire N__32844;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32830;
    wire N__32829;
    wire N__32826;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32809;
    wire N__32806;
    wire N__32801;
    wire N__32798;
    wire N__32791;
    wire N__32790;
    wire N__32789;
    wire N__32786;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32778;
    wire N__32777;
    wire N__32776;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32756;
    wire N__32755;
    wire N__32750;
    wire N__32741;
    wire N__32736;
    wire N__32735;
    wire N__32734;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32720;
    wire N__32717;
    wire N__32714;
    wire N__32713;
    wire N__32712;
    wire N__32709;
    wire N__32702;
    wire N__32699;
    wire N__32698;
    wire N__32697;
    wire N__32696;
    wire N__32691;
    wire N__32688;
    wire N__32685;
    wire N__32680;
    wire N__32679;
    wire N__32678;
    wire N__32675;
    wire N__32674;
    wire N__32671;
    wire N__32668;
    wire N__32667;
    wire N__32666;
    wire N__32663;
    wire N__32660;
    wire N__32659;
    wire N__32658;
    wire N__32657;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32643;
    wire N__32634;
    wire N__32631;
    wire N__32630;
    wire N__32629;
    wire N__32628;
    wire N__32627;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32599;
    wire N__32596;
    wire N__32595;
    wire N__32594;
    wire N__32593;
    wire N__32590;
    wire N__32589;
    wire N__32588;
    wire N__32587;
    wire N__32586;
    wire N__32583;
    wire N__32582;
    wire N__32581;
    wire N__32580;
    wire N__32577;
    wire N__32576;
    wire N__32573;
    wire N__32572;
    wire N__32571;
    wire N__32570;
    wire N__32565;
    wire N__32564;
    wire N__32561;
    wire N__32554;
    wire N__32547;
    wire N__32546;
    wire N__32545;
    wire N__32544;
    wire N__32543;
    wire N__32540;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32527;
    wire N__32526;
    wire N__32525;
    wire N__32524;
    wire N__32523;
    wire N__32522;
    wire N__32519;
    wire N__32518;
    wire N__32517;
    wire N__32516;
    wire N__32513;
    wire N__32508;
    wire N__32507;
    wire N__32506;
    wire N__32505;
    wire N__32504;
    wire N__32503;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32484;
    wire N__32483;
    wire N__32480;
    wire N__32477;
    wire N__32476;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32465;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32447;
    wire N__32446;
    wire N__32445;
    wire N__32444;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32434;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32418;
    wire N__32413;
    wire N__32412;
    wire N__32407;
    wire N__32404;
    wire N__32401;
    wire N__32396;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32373;
    wire N__32366;
    wire N__32361;
    wire N__32356;
    wire N__32351;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32334;
    wire N__32329;
    wire N__32326;
    wire N__32321;
    wire N__32320;
    wire N__32319;
    wire N__32318;
    wire N__32317;
    wire N__32316;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32297;
    wire N__32286;
    wire N__32281;
    wire N__32278;
    wire N__32267;
    wire N__32262;
    wire N__32251;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32221;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32203;
    wire N__32192;
    wire N__32189;
    wire N__32170;
    wire N__32167;
    wire N__32166;
    wire N__32163;
    wire N__32162;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32149;
    wire N__32140;
    wire N__32137;
    wire N__32134;
    wire N__32131;
    wire N__32128;
    wire N__32125;
    wire N__32124;
    wire N__32123;
    wire N__32122;
    wire N__32119;
    wire N__32116;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32108;
    wire N__32103;
    wire N__32100;
    wire N__32099;
    wire N__32098;
    wire N__32097;
    wire N__32092;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32079;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32061;
    wire N__32058;
    wire N__32047;
    wire N__32044;
    wire N__32041;
    wire N__32038;
    wire N__32035;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32011;
    wire N__32010;
    wire N__32007;
    wire N__32006;
    wire N__32003;
    wire N__32000;
    wire N__31999;
    wire N__31996;
    wire N__31993;
    wire N__31990;
    wire N__31987;
    wire N__31978;
    wire N__31975;
    wire N__31972;
    wire N__31969;
    wire N__31968;
    wire N__31967;
    wire N__31964;
    wire N__31959;
    wire N__31954;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31936;
    wire N__31933;
    wire N__31932;
    wire N__31931;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31906;
    wire N__31903;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31884;
    wire N__31883;
    wire N__31880;
    wire N__31875;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31858;
    wire N__31855;
    wire N__31854;
    wire N__31853;
    wire N__31850;
    wire N__31845;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31825;
    wire N__31824;
    wire N__31823;
    wire N__31820;
    wire N__31815;
    wire N__31810;
    wire N__31807;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31799;
    wire N__31796;
    wire N__31791;
    wire N__31786;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31768;
    wire N__31767;
    wire N__31764;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31731;
    wire N__31730;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31714;
    wire N__31711;
    wire N__31710;
    wire N__31709;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31693;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31672;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31652;
    wire N__31647;
    wire N__31644;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31623;
    wire N__31622;
    wire N__31619;
    wire N__31614;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31599;
    wire N__31598;
    wire N__31595;
    wire N__31590;
    wire N__31585;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31575;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31560;
    wire N__31555;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31543;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31517;
    wire N__31514;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31501;
    wire N__31496;
    wire N__31489;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31481;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31459;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31441;
    wire N__31440;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31417;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31402;
    wire N__31399;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31348;
    wire N__31345;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31331;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31313;
    wire N__31306;
    wire N__31305;
    wire N__31300;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31288;
    wire N__31285;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31252;
    wire N__31251;
    wire N__31248;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31237;
    wire N__31234;
    wire N__31229;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31204;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31190;
    wire N__31185;
    wire N__31184;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31156;
    wire N__31155;
    wire N__31154;
    wire N__31151;
    wire N__31146;
    wire N__31141;
    wire N__31138;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31121;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31107;
    wire N__31106;
    wire N__31103;
    wire N__31098;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31072;
    wire N__31069;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31049;
    wire N__31048;
    wire N__31045;
    wire N__31042;
    wire N__31037;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30992;
    wire N__30987;
    wire N__30984;
    wire N__30979;
    wire N__30976;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30940;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30930;
    wire N__30929;
    wire N__30926;
    wire N__30921;
    wire N__30916;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30908;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30896;
    wire N__30893;
    wire N__30886;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30865;
    wire N__30862;
    wire N__30857;
    wire N__30854;
    wire N__30851;
    wire N__30850;
    wire N__30849;
    wire N__30844;
    wire N__30841;
    wire N__30836;
    wire N__30833;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30811;
    wire N__30808;
    wire N__30807;
    wire N__30806;
    wire N__30803;
    wire N__30798;
    wire N__30793;
    wire N__30792;
    wire N__30789;
    wire N__30788;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30764;
    wire N__30757;
    wire N__30754;
    wire N__30753;
    wire N__30750;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30742;
    wire N__30739;
    wire N__30736;
    wire N__30733;
    wire N__30730;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30714;
    wire N__30713;
    wire N__30710;
    wire N__30705;
    wire N__30700;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30686;
    wire N__30681;
    wire N__30678;
    wire N__30673;
    wire N__30672;
    wire N__30669;
    wire N__30668;
    wire N__30665;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30626;
    wire N__30623;
    wire N__30616;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30580;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30572;
    wire N__30571;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30556;
    wire N__30547;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30530;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30518;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30497;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30468;
    wire N__30463;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30451;
    wire N__30450;
    wire N__30449;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30409;
    wire N__30406;
    wire N__30405;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30382;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30367;
    wire N__30358;
    wire N__30355;
    wire N__30354;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30284;
    wire N__30279;
    wire N__30276;
    wire N__30271;
    wire N__30268;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30260;
    wire N__30259;
    wire N__30258;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30243;
    wire N__30240;
    wire N__30233;
    wire N__30230;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30203;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30187;
    wire N__30186;
    wire N__30185;
    wire N__30182;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30164;
    wire N__30157;
    wire N__30154;
    wire N__30153;
    wire N__30150;
    wire N__30149;
    wire N__30148;
    wire N__30145;
    wire N__30142;
    wire N__30137;
    wire N__30134;
    wire N__30127;
    wire N__30124;
    wire N__30123;
    wire N__30120;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30100;
    wire N__30097;
    wire N__30092;
    wire N__30089;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30013;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29994;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29929;
    wire N__29928;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29911;
    wire N__29910;
    wire N__29907;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29890;
    wire N__29889;
    wire N__29886;
    wire N__29885;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29875;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29857;
    wire N__29854;
    wire N__29849;
    wire N__29846;
    wire N__29839;
    wire N__29838;
    wire N__29837;
    wire N__29834;
    wire N__29829;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29799;
    wire N__29796;
    wire N__29795;
    wire N__29794;
    wire N__29791;
    wire N__29790;
    wire N__29787;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29757;
    wire N__29752;
    wire N__29743;
    wire N__29740;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29713;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29703;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29676;
    wire N__29675;
    wire N__29674;
    wire N__29671;
    wire N__29666;
    wire N__29663;
    wire N__29656;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29645;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29629;
    wire N__29626;
    wire N__29625;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29608;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29551;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29539;
    wire N__29536;
    wire N__29535;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29527;
    wire N__29524;
    wire N__29519;
    wire N__29516;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29495;
    wire N__29488;
    wire N__29485;
    wire N__29484;
    wire N__29483;
    wire N__29480;
    wire N__29475;
    wire N__29472;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29457;
    wire N__29456;
    wire N__29455;
    wire N__29452;
    wire N__29447;
    wire N__29444;
    wire N__29437;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29399;
    wire N__29398;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29367;
    wire N__29366;
    wire N__29365;
    wire N__29362;
    wire N__29361;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29335;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29302;
    wire N__29299;
    wire N__29298;
    wire N__29295;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29284;
    wire N__29281;
    wire N__29276;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29250;
    wire N__29247;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29218;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29195;
    wire N__29194;
    wire N__29191;
    wire N__29188;
    wire N__29183;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29152;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29140;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29115;
    wire N__29114;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29102;
    wire N__29095;
    wire N__29092;
    wire N__29091;
    wire N__29088;
    wire N__29085;
    wire N__29082;
    wire N__29079;
    wire N__29078;
    wire N__29073;
    wire N__29070;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29044;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29032;
    wire N__29031;
    wire N__29030;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29019;
    wire N__29016;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28984;
    wire N__28975;
    wire N__28974;
    wire N__28973;
    wire N__28970;
    wire N__28965;
    wire N__28960;
    wire N__28959;
    wire N__28956;
    wire N__28955;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28917;
    wire N__28916;
    wire N__28915;
    wire N__28914;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28854;
    wire N__28853;
    wire N__28850;
    wire N__28849;
    wire N__28848;
    wire N__28845;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28813;
    wire N__28810;
    wire N__28809;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28793;
    wire N__28790;
    wire N__28789;
    wire N__28788;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28726;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28714;
    wire N__28711;
    wire N__28708;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28669;
    wire N__28666;
    wire N__28665;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28655;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28643;
    wire N__28636;
    wire N__28635;
    wire N__28632;
    wire N__28631;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28609;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28563;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28550;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28523;
    wire N__28518;
    wire N__28515;
    wire N__28510;
    wire N__28509;
    wire N__28506;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28458;
    wire N__28457;
    wire N__28456;
    wire N__28453;
    wire N__28448;
    wire N__28445;
    wire N__28438;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28424;
    wire N__28419;
    wire N__28416;
    wire N__28411;
    wire N__28410;
    wire N__28409;
    wire N__28406;
    wire N__28401;
    wire N__28396;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28382;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28367;
    wire N__28366;
    wire N__28361;
    wire N__28356;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28306;
    wire N__28305;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28273;
    wire N__28270;
    wire N__28261;
    wire N__28258;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28250;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28178;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28148;
    wire N__28145;
    wire N__28140;
    wire N__28137;
    wire N__28132;
    wire N__28131;
    wire N__28130;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28108;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28078;
    wire N__28075;
    wire N__28074;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28050;
    wire N__28047;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28035;
    wire N__28030;
    wire N__28029;
    wire N__28026;
    wire N__28025;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28004;
    wire N__28003;
    wire N__28000;
    wire N__27995;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27966;
    wire N__27963;
    wire N__27960;
    wire N__27957;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27928;
    wire N__27927;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27919;
    wire N__27916;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27899;
    wire N__27892;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27869;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27857;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27837;
    wire N__27836;
    wire N__27835;
    wire N__27832;
    wire N__27825;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27779;
    wire N__27772;
    wire N__27769;
    wire N__27768;
    wire N__27763;
    wire N__27760;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27748;
    wire N__27745;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27721;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27706;
    wire N__27703;
    wire N__27698;
    wire N__27695;
    wire N__27688;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27661;
    wire N__27658;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27650;
    wire N__27645;
    wire N__27642;
    wire N__27641;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27613;
    wire N__27612;
    wire N__27609;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27586;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27578;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27550;
    wire N__27547;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27529;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27517;
    wire N__27514;
    wire N__27513;
    wire N__27510;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27493;
    wire N__27490;
    wire N__27489;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27456;
    wire N__27455;
    wire N__27454;
    wire N__27451;
    wire N__27446;
    wire N__27443;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27426;
    wire N__27425;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27414;
    wire N__27411;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27354;
    wire N__27353;
    wire N__27350;
    wire N__27345;
    wire N__27340;
    wire N__27337;
    wire N__27336;
    wire N__27335;
    wire N__27334;
    wire N__27331;
    wire N__27324;
    wire N__27319;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27311;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27297;
    wire N__27296;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27240;
    wire N__27239;
    wire N__27236;
    wire N__27231;
    wire N__27226;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27218;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27180;
    wire N__27179;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27161;
    wire N__27154;
    wire N__27151;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27139;
    wire N__27138;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27130;
    wire N__27127;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27099;
    wire N__27094;
    wire N__27085;
    wire N__27082;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27042;
    wire N__27039;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27016;
    wire N__27013;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26999;
    wire N__26998;
    wire N__26993;
    wire N__26988;
    wire N__26983;
    wire N__26982;
    wire N__26979;
    wire N__26978;
    wire N__26975;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26946;
    wire N__26945;
    wire N__26942;
    wire N__26937;
    wire N__26936;
    wire N__26931;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26878;
    wire N__26875;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26835;
    wire N__26832;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26816;
    wire N__26809;
    wire N__26808;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26796;
    wire N__26795;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26764;
    wire N__26763;
    wire N__26760;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26748;
    wire N__26745;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26730;
    wire N__26729;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26664;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26656;
    wire N__26655;
    wire N__26652;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26574;
    wire N__26571;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26538;
    wire N__26537;
    wire N__26534;
    wire N__26529;
    wire N__26524;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26510;
    wire N__26505;
    wire N__26502;
    wire N__26497;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26457;
    wire N__26456;
    wire N__26453;
    wire N__26448;
    wire N__26443;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26395;
    wire N__26394;
    wire N__26393;
    wire N__26390;
    wire N__26385;
    wire N__26380;
    wire N__26379;
    wire N__26376;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26365;
    wire N__26364;
    wire N__26361;
    wire N__26356;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26329;
    wire N__26326;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26307;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26295;
    wire N__26292;
    wire N__26289;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26264;
    wire N__26261;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26247;
    wire N__26242;
    wire N__26237;
    wire N__26234;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26218;
    wire N__26215;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26199;
    wire N__26196;
    wire N__26195;
    wire N__26190;
    wire N__26187;
    wire N__26182;
    wire N__26179;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26167;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26155;
    wire N__26154;
    wire N__26151;
    wire N__26150;
    wire N__26147;
    wire N__26144;
    wire N__26143;
    wire N__26140;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26118;
    wire N__26113;
    wire N__26112;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26071;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26050;
    wire N__26047;
    wire N__26044;
    wire N__26043;
    wire N__26040;
    wire N__26039;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26027;
    wire N__26020;
    wire N__26019;
    wire N__26018;
    wire N__26013;
    wire N__26010;
    wire N__26005;
    wire N__26004;
    wire N__25999;
    wire N__25998;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25960;
    wire N__25957;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25939;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25912;
    wire N__25911;
    wire N__25908;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25885;
    wire N__25882;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25871;
    wire N__25870;
    wire N__25867;
    wire N__25864;
    wire N__25859;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25836;
    wire N__25835;
    wire N__25832;
    wire N__25827;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25792;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25763;
    wire N__25760;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25749;
    wire N__25746;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25726;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25692;
    wire N__25691;
    wire N__25688;
    wire N__25683;
    wire N__25678;
    wire N__25677;
    wire N__25676;
    wire N__25673;
    wire N__25672;
    wire N__25669;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25629;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25601;
    wire N__25596;
    wire N__25593;
    wire N__25588;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25578;
    wire N__25577;
    wire N__25574;
    wire N__25569;
    wire N__25564;
    wire N__25561;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25553;
    wire N__25552;
    wire N__25549;
    wire N__25546;
    wire N__25541;
    wire N__25534;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25519;
    wire N__25516;
    wire N__25511;
    wire N__25508;
    wire N__25501;
    wire N__25498;
    wire N__25497;
    wire N__25494;
    wire N__25493;
    wire N__25492;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25469;
    wire N__25466;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25452;
    wire N__25451;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25435;
    wire N__25432;
    wire N__25427;
    wire N__25424;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25381;
    wire N__25378;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25367;
    wire N__25366;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25351;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25332;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25315;
    wire N__25312;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25294;
    wire N__25293;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25251;
    wire N__25250;
    wire N__25249;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25200;
    wire N__25197;
    wire N__25196;
    wire N__25193;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25171;
    wire N__25162;
    wire N__25161;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25107;
    wire N__25106;
    wire N__25105;
    wire N__25104;
    wire N__25101;
    wire N__25096;
    wire N__25091;
    wire N__25084;
    wire N__25081;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25056;
    wire N__25053;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25039;
    wire N__25038;
    wire N__25033;
    wire N__25030;
    wire N__25025;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25008;
    wire N__25005;
    wire N__25004;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24983;
    wire N__24980;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24960;
    wire N__24957;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24944;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24932;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24920;
    wire N__24913;
    wire N__24910;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24898;
    wire N__24895;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24887;
    wire N__24886;
    wire N__24885;
    wire N__24880;
    wire N__24877;
    wire N__24872;
    wire N__24865;
    wire N__24862;
    wire N__24859;
    wire N__24856;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24840;
    wire N__24837;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24829;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24805;
    wire N__24802;
    wire N__24793;
    wire N__24790;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24757;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24740;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24699;
    wire N__24698;
    wire N__24697;
    wire N__24694;
    wire N__24687;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24640;
    wire N__24639;
    wire N__24636;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24618;
    wire N__24617;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24605;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24528;
    wire N__24525;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24505;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24489;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24447;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24435;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24420;
    wire N__24417;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24381;
    wire N__24376;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24364;
    wire N__24363;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24328;
    wire N__24327;
    wire N__24324;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24307;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24293;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24250;
    wire N__24247;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24235;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24223;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24212;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24184;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24154;
    wire N__24151;
    wire N__24150;
    wire N__24147;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24118;
    wire N__24115;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24085;
    wire N__24082;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24068;
    wire N__24067;
    wire N__24062;
    wire N__24057;
    wire N__24052;
    wire N__24049;
    wire N__24048;
    wire N__24047;
    wire N__24044;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24034;
    wire N__24031;
    wire N__24026;
    wire N__24019;
    wire N__24016;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24004;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23979;
    wire N__23976;
    wire N__23973;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23949;
    wire N__23948;
    wire N__23945;
    wire N__23940;
    wire N__23937;
    wire N__23932;
    wire N__23929;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23921;
    wire N__23920;
    wire N__23915;
    wire N__23912;
    wire N__23911;
    wire N__23908;
    wire N__23903;
    wire N__23900;
    wire N__23893;
    wire N__23892;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23868;
    wire N__23865;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23845;
    wire N__23844;
    wire N__23841;
    wire N__23838;
    wire N__23835;
    wire N__23832;
    wire N__23829;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23802;
    wire N__23801;
    wire N__23798;
    wire N__23793;
    wire N__23788;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23774;
    wire N__23773;
    wire N__23768;
    wire N__23763;
    wire N__23758;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23740;
    wire N__23739;
    wire N__23736;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23656;
    wire N__23653;
    wire N__23652;
    wire N__23651;
    wire N__23648;
    wire N__23643;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23619;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23604;
    wire N__23601;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23554;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23539;
    wire N__23536;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23512;
    wire N__23509;
    wire N__23500;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23492;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23472;
    wire N__23469;
    wire N__23468;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23456;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23436;
    wire N__23433;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23358;
    wire N__23355;
    wire N__23354;
    wire N__23353;
    wire N__23350;
    wire N__23347;
    wire N__23342;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23256;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23248;
    wire N__23245;
    wire N__23240;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23222;
    wire N__23215;
    wire N__23212;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23112;
    wire N__23111;
    wire N__23108;
    wire N__23103;
    wire N__23098;
    wire N__23095;
    wire N__23094;
    wire N__23093;
    wire N__23090;
    wire N__23085;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23033;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22997;
    wire N__22996;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22982;
    wire N__22975;
    wire N__22972;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22954;
    wire N__22951;
    wire N__22950;
    wire N__22947;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22936;
    wire N__22933;
    wire N__22928;
    wire N__22927;
    wire N__22926;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22911;
    wire N__22906;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22869;
    wire N__22866;
    wire N__22865;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22834;
    wire N__22831;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22823;
    wire N__22822;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22807;
    wire N__22800;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22778;
    wire N__22773;
    wire N__22770;
    wire N__22769;
    wire N__22768;
    wire N__22763;
    wire N__22758;
    wire N__22755;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22695;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22678;
    wire N__22675;
    wire N__22672;
    wire N__22671;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22663;
    wire N__22660;
    wire N__22655;
    wire N__22652;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22623;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22603;
    wire N__22598;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22573;
    wire N__22572;
    wire N__22571;
    wire N__22568;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22541;
    wire N__22534;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22468;
    wire N__22465;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22441;
    wire N__22438;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22375;
    wire N__22372;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22364;
    wire N__22363;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22347;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22308;
    wire N__22307;
    wire N__22304;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22282;
    wire N__22281;
    wire N__22278;
    wire N__22273;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22246;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22198;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22190;
    wire N__22189;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22161;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22146;
    wire N__22145;
    wire N__22142;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22078;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21955;
    wire N__21954;
    wire N__21951;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21935;
    wire N__21932;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21883;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21875;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21863;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21837;
    wire N__21836;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21810;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21735;
    wire N__21734;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21722;
    wire N__21715;
    wire N__21712;
    wire N__21711;
    wire N__21708;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21687;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21652;
    wire N__21649;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21617;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21605;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21581;
    wire N__21580;
    wire N__21579;
    wire N__21574;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21522;
    wire N__21521;
    wire N__21518;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21463;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21446;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21434;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21417;
    wire N__21416;
    wire N__21415;
    wire N__21414;
    wire N__21413;
    wire N__21412;
    wire N__21409;
    wire N__21408;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21381;
    wire N__21380;
    wire N__21379;
    wire N__21376;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21353;
    wire N__21346;
    wire N__21345;
    wire N__21340;
    wire N__21335;
    wire N__21332;
    wire N__21325;
    wire N__21322;
    wire N__21321;
    wire N__21320;
    wire N__21319;
    wire N__21318;
    wire N__21315;
    wire N__21314;
    wire N__21313;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21289;
    wire N__21288;
    wire N__21283;
    wire N__21280;
    wire N__21275;
    wire N__21270;
    wire N__21267;
    wire N__21262;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21250;
    wire N__21247;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21231;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21195;
    wire N__21192;
    wire N__21191;
    wire N__21190;
    wire N__21189;
    wire N__21188;
    wire N__21187;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21149;
    wire N__21148;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21123;
    wire N__21120;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21105;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21079;
    wire N__21078;
    wire N__21077;
    wire N__21076;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21045;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21030;
    wire N__21027;
    wire N__21016;
    wire N__21013;
    wire N__21012;
    wire N__21009;
    wire N__21008;
    wire N__21007;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20995;
    wire N__20992;
    wire N__20983;
    wire N__20980;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20931;
    wire N__20930;
    wire N__20927;
    wire N__20922;
    wire N__20917;
    wire N__20916;
    wire N__20915;
    wire N__20912;
    wire N__20911;
    wire N__20908;
    wire N__20903;
    wire N__20900;
    wire N__20899;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20882;
    wire N__20877;
    wire N__20874;
    wire N__20863;
    wire N__20860;
    wire N__20859;
    wire N__20854;
    wire N__20851;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20839;
    wire N__20836;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20824;
    wire N__20821;
    wire N__20820;
    wire N__20815;
    wire N__20812;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20798;
    wire N__20793;
    wire N__20790;
    wire N__20785;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20749;
    wire N__20748;
    wire N__20745;
    wire N__20744;
    wire N__20743;
    wire N__20740;
    wire N__20739;
    wire N__20736;
    wire N__20731;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20719;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20647;
    wire N__20644;
    wire N__20643;
    wire N__20642;
    wire N__20641;
    wire N__20640;
    wire N__20639;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20611;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20599;
    wire N__20596;
    wire N__20587;
    wire N__20586;
    wire N__20585;
    wire N__20584;
    wire N__20583;
    wire N__20582;
    wire N__20581;
    wire N__20580;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20572;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20540;
    wire N__20531;
    wire N__20530;
    wire N__20525;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20511;
    wire N__20510;
    wire N__20509;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20497;
    wire N__20490;
    wire N__20487;
    wire N__20476;
    wire N__20475;
    wire N__20472;
    wire N__20471;
    wire N__20470;
    wire N__20469;
    wire N__20468;
    wire N__20463;
    wire N__20460;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20427;
    wire N__20416;
    wire N__20415;
    wire N__20414;
    wire N__20413;
    wire N__20412;
    wire N__20411;
    wire N__20410;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20406;
    wire N__20405;
    wire N__20404;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20393;
    wire N__20392;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20380;
    wire N__20373;
    wire N__20368;
    wire N__20363;
    wire N__20356;
    wire N__20355;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20334;
    wire N__20329;
    wire N__20326;
    wire N__20325;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20310;
    wire N__20305;
    wire N__20300;
    wire N__20297;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20265;
    wire N__20264;
    wire N__20263;
    wire N__20260;
    wire N__20253;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20191;
    wire N__20188;
    wire N__20187;
    wire N__20186;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20164;
    wire N__20163;
    wire N__20160;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20124;
    wire N__20119;
    wire N__20116;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20089;
    wire N__20086;
    wire N__20085;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20071;
    wire N__20068;
    wire N__20063;
    wire N__20060;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20043;
    wire N__20042;
    wire N__20041;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20026;
    wire N__20017;
    wire N__20014;
    wire N__20013;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19984;
    wire N__19983;
    wire N__19980;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19958;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19924;
    wire N__19923;
    wire N__19922;
    wire N__19919;
    wire N__19914;
    wire N__19909;
    wire N__19906;
    wire N__19905;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19884;
    wire N__19881;
    wire N__19878;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19830;
    wire N__19827;
    wire N__19826;
    wire N__19825;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19811;
    wire N__19804;
    wire N__19801;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19793;
    wire N__19792;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19777;
    wire N__19772;
    wire N__19769;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19670;
    wire N__19669;
    wire N__19668;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19645;
    wire N__19642;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19630;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19615;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19603;
    wire N__19602;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19585;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19507;
    wire N__19504;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19371;
    wire N__19370;
    wire N__19369;
    wire N__19368;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19346;
    wire N__19343;
    wire N__19342;
    wire N__19341;
    wire N__19340;
    wire N__19337;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19312;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19300;
    wire N__19299;
    wire N__19298;
    wire N__19297;
    wire N__19296;
    wire N__19293;
    wire N__19292;
    wire N__19287;
    wire N__19284;
    wire N__19283;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19257;
    wire N__19252;
    wire N__19249;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19224;
    wire N__19223;
    wire N__19222;
    wire N__19221;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19213;
    wire N__19210;
    wire N__19209;
    wire N__19208;
    wire N__19207;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19181;
    wire N__19180;
    wire N__19179;
    wire N__19178;
    wire N__19177;
    wire N__19176;
    wire N__19175;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19167;
    wire N__19160;
    wire N__19153;
    wire N__19142;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19118;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19087;
    wire N__19084;
    wire N__19083;
    wire N__19082;
    wire N__19081;
    wire N__19080;
    wire N__19079;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19058;
    wire N__19057;
    wire N__19056;
    wire N__19051;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19035;
    wire N__19034;
    wire N__19033;
    wire N__19032;
    wire N__19031;
    wire N__19030;
    wire N__19029;
    wire N__19028;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19016;
    wire N__19013;
    wire N__19008;
    wire N__18997;
    wire N__18994;
    wire N__18979;
    wire N__18978;
    wire N__18977;
    wire N__18976;
    wire N__18973;
    wire N__18968;
    wire N__18967;
    wire N__18964;
    wire N__18959;
    wire N__18956;
    wire N__18955;
    wire N__18954;
    wire N__18951;
    wire N__18946;
    wire N__18943;
    wire N__18940;
    wire N__18935;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18874;
    wire N__18871;
    wire N__18870;
    wire N__18865;
    wire N__18862;
    wire N__18861;
    wire N__18858;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18832;
    wire N__18829;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18817;
    wire N__18814;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18806;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18796;
    wire N__18793;
    wire N__18792;
    wire N__18785;
    wire N__18782;
    wire N__18781;
    wire N__18780;
    wire N__18779;
    wire N__18776;
    wire N__18771;
    wire N__18768;
    wire N__18763;
    wire N__18754;
    wire N__18751;
    wire N__18750;
    wire N__18749;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18735;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18568;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18538;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18517;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18505;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18490;
    wire N__18487;
    wire N__18486;
    wire N__18483;
    wire N__18480;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18412;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18367;
    wire N__18364;
    wire N__18363;
    wire N__18362;
    wire N__18361;
    wire N__18358;
    wire N__18357;
    wire N__18356;
    wire N__18355;
    wire N__18354;
    wire N__18349;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18330;
    wire N__18329;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18314;
    wire N__18309;
    wire N__18306;
    wire N__18301;
    wire N__18292;
    wire N__18283;
    wire N__18282;
    wire N__18281;
    wire N__18280;
    wire N__18279;
    wire N__18278;
    wire N__18277;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18269;
    wire N__18268;
    wire N__18267;
    wire N__18266;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18248;
    wire N__18247;
    wire N__18246;
    wire N__18243;
    wire N__18238;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18220;
    wire N__18217;
    wire N__18210;
    wire N__18205;
    wire N__18190;
    wire N__18187;
    wire N__18184;
    wire N__18181;
    wire N__18180;
    wire N__18179;
    wire N__18178;
    wire N__18177;
    wire N__18176;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18152;
    wire N__18149;
    wire N__18144;
    wire N__18139;
    wire N__18138;
    wire N__18137;
    wire N__18136;
    wire N__18133;
    wire N__18132;
    wire N__18131;
    wire N__18130;
    wire N__18125;
    wire N__18120;
    wire N__18117;
    wire N__18116;
    wire N__18113;
    wire N__18112;
    wire N__18111;
    wire N__18110;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18098;
    wire N__18091;
    wire N__18086;
    wire N__18083;
    wire N__18070;
    wire N__18067;
    wire N__18066;
    wire N__18065;
    wire N__18062;
    wire N__18057;
    wire N__18056;
    wire N__18055;
    wire N__18050;
    wire N__18049;
    wire N__18048;
    wire N__18047;
    wire N__18046;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18030;
    wire N__18027;
    wire N__18016;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18004;
    wire N__18001;
    wire N__17998;
    wire N__17995;
    wire N__17994;
    wire N__17991;
    wire N__17988;
    wire N__17983;
    wire N__17982;
    wire N__17981;
    wire N__17978;
    wire N__17973;
    wire N__17968;
    wire N__17965;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17953;
    wire N__17952;
    wire N__17949;
    wire N__17948;
    wire N__17945;
    wire N__17940;
    wire N__17935;
    wire N__17934;
    wire N__17931;
    wire N__17928;
    wire N__17925;
    wire N__17922;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17890;
    wire N__17887;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17877;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17867;
    wire N__17866;
    wire N__17863;
    wire N__17860;
    wire N__17855;
    wire N__17852;
    wire N__17845;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17837;
    wire N__17836;
    wire N__17833;
    wire N__17830;
    wire N__17827;
    wire N__17824;
    wire N__17815;
    wire N__17812;
    wire N__17809;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17797;
    wire N__17794;
    wire N__17791;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17764;
    wire N__17761;
    wire N__17758;
    wire N__17755;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17743;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17733;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17725;
    wire N__17722;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17685;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17595;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17562;
    wire N__17561;
    wire N__17560;
    wire N__17559;
    wire N__17556;
    wire N__17547;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17535;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17509;
    wire N__17508;
    wire N__17507;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17499;
    wire N__17496;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17473;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17436;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17422;
    wire N__17421;
    wire N__17418;
    wire N__17413;
    wire N__17408;
    wire N__17401;
    wire N__17398;
    wire N__17397;
    wire N__17394;
    wire N__17391;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17360;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17341;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17319;
    wire N__17318;
    wire N__17317;
    wire N__17310;
    wire N__17307;
    wire N__17302;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17277;
    wire N__17274;
    wire N__17271;
    wire N__17266;
    wire N__17265;
    wire N__17260;
    wire N__17257;
    wire N__17256;
    wire N__17253;
    wire N__17250;
    wire N__17247;
    wire N__17242;
    wire N__17239;
    wire N__17238;
    wire N__17237;
    wire N__17236;
    wire N__17235;
    wire N__17234;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17191;
    wire N__17190;
    wire N__17187;
    wire N__17186;
    wire N__17185;
    wire N__17184;
    wire N__17183;
    wire N__17180;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17151;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17121;
    wire N__17120;
    wire N__17119;
    wire N__17118;
    wire N__17117;
    wire N__17116;
    wire N__17111;
    wire N__17104;
    wire N__17101;
    wire N__17100;
    wire N__17099;
    wire N__17098;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17086;
    wire N__17081;
    wire N__17076;
    wire N__17065;
    wire N__17062;
    wire N__17061;
    wire N__17060;
    wire N__17059;
    wire N__17058;
    wire N__17055;
    wire N__17052;
    wire N__17051;
    wire N__17050;
    wire N__17049;
    wire N__17046;
    wire N__17045;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17017;
    wire N__17002;
    wire N__17001;
    wire N__17000;
    wire N__16999;
    wire N__16998;
    wire N__16997;
    wire N__16996;
    wire N__16993;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16985;
    wire N__16984;
    wire N__16983;
    wire N__16980;
    wire N__16979;
    wire N__16978;
    wire N__16977;
    wire N__16974;
    wire N__16973;
    wire N__16972;
    wire N__16969;
    wire N__16968;
    wire N__16967;
    wire N__16962;
    wire N__16959;
    wire N__16950;
    wire N__16949;
    wire N__16946;
    wire N__16937;
    wire N__16932;
    wire N__16923;
    wire N__16920;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16894;
    wire N__16891;
    wire N__16890;
    wire N__16887;
    wire N__16884;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16858;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16846;
    wire N__16843;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16818;
    wire N__16813;
    wire N__16810;
    wire N__16809;
    wire N__16808;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16797;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16779;
    wire N__16770;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16741;
    wire N__16738;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16728;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16703;
    wire N__16700;
    wire N__16695;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16680;
    wire N__16679;
    wire N__16678;
    wire N__16677;
    wire N__16674;
    wire N__16673;
    wire N__16672;
    wire N__16671;
    wire N__16670;
    wire N__16669;
    wire N__16668;
    wire N__16667;
    wire N__16666;
    wire N__16665;
    wire N__16664;
    wire N__16663;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16631;
    wire N__16626;
    wire N__16621;
    wire N__16600;
    wire N__16599;
    wire N__16596;
    wire N__16591;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16581;
    wire N__16580;
    wire N__16579;
    wire N__16576;
    wire N__16571;
    wire N__16570;
    wire N__16567;
    wire N__16566;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16546;
    wire N__16541;
    wire N__16538;
    wire N__16533;
    wire N__16530;
    wire N__16519;
    wire N__16516;
    wire N__16515;
    wire N__16514;
    wire N__16513;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16489;
    wire N__16486;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16470;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16434;
    wire N__16433;
    wire N__16432;
    wire N__16431;
    wire N__16430;
    wire N__16427;
    wire N__16420;
    wire N__16417;
    wire N__16416;
    wire N__16415;
    wire N__16412;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16371;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16363;
    wire N__16360;
    wire N__16355;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16284;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16273;
    wire N__16272;
    wire N__16271;
    wire N__16264;
    wire N__16261;
    wire N__16256;
    wire N__16253;
    wire N__16246;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16227;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16171;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16156;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16126;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16111;
    wire N__16108;
    wire N__16107;
    wire N__16104;
    wire N__16103;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16091;
    wire N__16084;
    wire N__16081;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16035;
    wire N__16030;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16015;
    wire N__16012;
    wire N__16011;
    wire N__16008;
    wire N__16005;
    wire N__16002;
    wire N__15997;
    wire N__15994;
    wire N__15993;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15979;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15963;
    wire N__15960;
    wire N__15959;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15928;
    wire N__15925;
    wire N__15922;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15861;
    wire N__15858;
    wire N__15857;
    wire N__15854;
    wire N__15853;
    wire N__15850;
    wire N__15847;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15829;
    wire N__15826;
    wire N__15823;
    wire N__15822;
    wire N__15821;
    wire N__15818;
    wire N__15813;
    wire N__15810;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15783;
    wire N__15782;
    wire N__15781;
    wire N__15780;
    wire N__15777;
    wire N__15772;
    wire N__15767;
    wire N__15762;
    wire N__15757;
    wire N__15756;
    wire N__15753;
    wire N__15750;
    wire N__15749;
    wire N__15744;
    wire N__15741;
    wire N__15738;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15702;
    wire N__15701;
    wire N__15700;
    wire N__15697;
    wire N__15690;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15675;
    wire N__15670;
    wire N__15667;
    wire N__15666;
    wire N__15665;
    wire N__15664;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15639;
    wire N__15634;
    wire N__15633;
    wire N__15632;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15624;
    wire N__15619;
    wire N__15614;
    wire N__15611;
    wire N__15604;
    wire N__15603;
    wire N__15602;
    wire N__15599;
    wire N__15598;
    wire N__15595;
    wire N__15594;
    wire N__15591;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15576;
    wire N__15573;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15561;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15538;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15530;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15508;
    wire N__15505;
    wire N__15502;
    wire N__15499;
    wire N__15496;
    wire N__15493;
    wire N__15490;
    wire N__15487;
    wire N__15486;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15469;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15435;
    wire N__15432;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15405;
    wire N__15404;
    wire N__15403;
    wire N__15402;
    wire N__15393;
    wire N__15390;
    wire N__15385;
    wire N__15382;
    wire N__15379;
    wire N__15376;
    wire N__15373;
    wire N__15370;
    wire N__15367;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15357;
    wire N__15354;
    wire N__15351;
    wire N__15348;
    wire N__15343;
    wire N__15342;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15328;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15309;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15297;
    wire N__15292;
    wire N__15289;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15265;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15250;
    wire N__15249;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15235;
    wire N__15232;
    wire N__15231;
    wire N__15226;
    wire N__15223;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15211;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15193;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15181;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15137;
    wire N__15130;
    wire N__15127;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15115;
    wire N__15112;
    wire N__15111;
    wire N__15108;
    wire N__15105;
    wire N__15100;
    wire N__15097;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15085;
    wire N__15082;
    wire N__15081;
    wire N__15078;
    wire N__15075;
    wire N__15072;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15057;
    wire N__15054;
    wire N__15051;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15037;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15025;
    wire N__15022;
    wire N__15021;
    wire N__15018;
    wire N__15015;
    wire N__15012;
    wire N__15009;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14988;
    wire N__14985;
    wire N__14982;
    wire N__14977;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14967;
    wire N__14966;
    wire N__14965;
    wire N__14964;
    wire N__14963;
    wire N__14962;
    wire N__14951;
    wire N__14946;
    wire N__14941;
    wire N__14940;
    wire N__14939;
    wire N__14938;
    wire N__14935;
    wire N__14934;
    wire N__14933;
    wire N__14924;
    wire N__14919;
    wire N__14914;
    wire N__14913;
    wire N__14912;
    wire N__14911;
    wire N__14908;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14884;
    wire N__14883;
    wire N__14882;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14835;
    wire N__14832;
    wire N__14829;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14782;
    wire N__14779;
    wire N__14778;
    wire N__14775;
    wire N__14772;
    wire N__14767;
    wire N__14766;
    wire N__14765;
    wire N__14762;
    wire N__14761;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14731;
    wire N__14730;
    wire N__14729;
    wire N__14726;
    wire N__14725;
    wire N__14724;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14710;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14691;
    wire N__14690;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14678;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14661;
    wire N__14658;
    wire N__14655;
    wire N__14652;
    wire N__14647;
    wire N__14646;
    wire N__14643;
    wire N__14640;
    wire N__14639;
    wire N__14636;
    wire N__14635;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14527;
    wire N__14526;
    wire N__14525;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14511;
    wire N__14510;
    wire N__14509;
    wire N__14506;
    wire N__14505;
    wire N__14500;
    wire N__14497;
    wire N__14490;
    wire N__14487;
    wire N__14484;
    wire N__14481;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14427;
    wire N__14424;
    wire N__14421;
    wire N__14418;
    wire N__14415;
    wire N__14412;
    wire N__14407;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14397;
    wire N__14394;
    wire N__14393;
    wire N__14392;
    wire N__14391;
    wire N__14390;
    wire N__14389;
    wire N__14388;
    wire N__14387;
    wire N__14386;
    wire N__14385;
    wire N__14382;
    wire N__14379;
    wire N__14372;
    wire N__14369;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14339;
    wire N__14326;
    wire N__14323;
    wire N__14322;
    wire N__14319;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14303;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14262;
    wire N__14261;
    wire N__14260;
    wire N__14259;
    wire N__14258;
    wire N__14257;
    wire N__14256;
    wire N__14255;
    wire N__14254;
    wire N__14253;
    wire N__14252;
    wire N__14251;
    wire N__14250;
    wire N__14249;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14241;
    wire N__14240;
    wire N__14239;
    wire N__14238;
    wire N__14237;
    wire N__14236;
    wire N__14235;
    wire N__14234;
    wire N__14233;
    wire N__14232;
    wire N__14229;
    wire N__14226;
    wire N__14223;
    wire N__14220;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14181;
    wire N__14174;
    wire N__14169;
    wire N__14162;
    wire N__14153;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14128;
    wire N__14121;
    wire N__14114;
    wire N__14101;
    wire N__14098;
    wire N__14097;
    wire N__14096;
    wire N__14093;
    wire N__14088;
    wire N__14087;
    wire N__14086;
    wire N__14085;
    wire N__14084;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14068;
    wire N__14065;
    wire N__14056;
    wire N__14055;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14025;
    wire N__14024;
    wire N__14023;
    wire N__14022;
    wire N__14019;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__13999;
    wire N__13996;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13984;
    wire N__13983;
    wire N__13982;
    wire N__13981;
    wire N__13980;
    wire N__13979;
    wire N__13978;
    wire N__13977;
    wire N__13976;
    wire N__13973;
    wire N__13968;
    wire N__13963;
    wire N__13954;
    wire N__13951;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13926;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13902;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13878;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13861;
    wire N__13860;
    wire N__13857;
    wire N__13856;
    wire N__13855;
    wire N__13854;
    wire N__13853;
    wire N__13852;
    wire N__13851;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13831;
    wire N__13826;
    wire N__13819;
    wire N__13816;
    wire N__13807;
    wire N__13806;
    wire N__13805;
    wire N__13804;
    wire N__13803;
    wire N__13796;
    wire N__13795;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13777;
    wire N__13776;
    wire N__13773;
    wire N__13770;
    wire N__13765;
    wire N__13762;
    wire N__13761;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13725;
    wire N__13724;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13710;
    wire N__13703;
    wire N__13702;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13684;
    wire N__13681;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13662;
    wire N__13657;
    wire N__13656;
    wire N__13655;
    wire N__13654;
    wire N__13651;
    wire N__13646;
    wire N__13643;
    wire N__13642;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13627;
    wire N__13618;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13606;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13594;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13582;
    wire N__13581;
    wire N__13580;
    wire N__13579;
    wire N__13576;
    wire N__13571;
    wire N__13568;
    wire N__13561;
    wire N__13560;
    wire N__13557;
    wire N__13554;
    wire N__13549;
    wire N__13546;
    wire N__13543;
    wire N__13542;
    wire N__13541;
    wire N__13540;
    wire N__13539;
    wire N__13534;
    wire N__13529;
    wire N__13526;
    wire N__13519;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13492;
    wire N__13489;
    wire N__13486;
    wire N__13485;
    wire N__13482;
    wire N__13479;
    wire N__13478;
    wire N__13477;
    wire N__13476;
    wire N__13465;
    wire N__13462;
    wire N__13459;
    wire N__13456;
    wire N__13453;
    wire N__13450;
    wire N__13449;
    wire N__13448;
    wire N__13441;
    wire N__13440;
    wire N__13439;
    wire N__13436;
    wire N__13431;
    wire N__13428;
    wire N__13423;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13411;
    wire N__13410;
    wire N__13407;
    wire N__13404;
    wire N__13399;
    wire N__13398;
    wire N__13397;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13384;
    wire N__13375;
    wire N__13374;
    wire N__13373;
    wire N__13372;
    wire N__13369;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13351;
    wire N__13348;
    wire N__13345;
    wire N__13344;
    wire N__13341;
    wire N__13340;
    wire N__13339;
    wire N__13338;
    wire N__13335;
    wire N__13332;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13312;
    wire N__13309;
    wire N__13308;
    wire N__13307;
    wire N__13306;
    wire N__13305;
    wire N__13302;
    wire N__13299;
    wire N__13296;
    wire N__13291;
    wire N__13282;
    wire N__13281;
    wire N__13280;
    wire N__13279;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13265;
    wire N__13258;
    wire N__13255;
    wire N__13252;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13242;
    wire N__13241;
    wire N__13240;
    wire N__13239;
    wire N__13238;
    wire N__13233;
    wire N__13226;
    wire N__13225;
    wire N__13224;
    wire N__13223;
    wire N__13222;
    wire N__13219;
    wire N__13216;
    wire N__13213;
    wire N__13206;
    wire N__13203;
    wire N__13192;
    wire N__13189;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13138;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13123;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13108;
    wire N__13105;
    wire N__13102;
    wire N__13099;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13087;
    wire N__13084;
    wire N__13083;
    wire N__13080;
    wire N__13077;
    wire N__13074;
    wire N__13069;
    wire N__13066;
    wire N__13063;
    wire N__13060;
    wire N__13059;
    wire N__13058;
    wire N__13057;
    wire N__13056;
    wire N__13049;
    wire N__13048;
    wire N__13047;
    wire N__13046;
    wire N__13045;
    wire N__13042;
    wire N__13039;
    wire N__13036;
    wire N__13029;
    wire N__13026;
    wire N__13021;
    wire N__13012;
    wire N__13009;
    wire N__13006;
    wire N__13003;
    wire N__13000;
    wire N__12997;
    wire N__12994;
    wire N__12993;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12982;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12963;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12937;
    wire N__12934;
    wire N__12931;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12916;
    wire N__12913;
    wire N__12910;
    wire N__12907;
    wire N__12904;
    wire N__12901;
    wire N__12898;
    wire N__12895;
    wire N__12892;
    wire N__12889;
    wire N__12886;
    wire N__12885;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12865;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12853;
    wire N__12850;
    wire N__12849;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12832;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12819;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12802;
    wire N__12799;
    wire N__12796;
    wire N__12793;
    wire N__12790;
    wire N__12789;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12772;
    wire N__12769;
    wire N__12766;
    wire N__12763;
    wire N__12760;
    wire N__12757;
    wire N__12756;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12748;
    wire N__12745;
    wire N__12740;
    wire N__12737;
    wire N__12730;
    wire N__12727;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12673;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12643;
    wire N__12640;
    wire N__12637;
    wire N__12634;
    wire N__12631;
    wire N__12630;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12613;
    wire N__12612;
    wire N__12611;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12595;
    wire N__12594;
    wire N__12591;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12571;
    wire N__12570;
    wire N__12569;
    wire N__12566;
    wire N__12561;
    wire N__12556;
    wire N__12555;
    wire N__12554;
    wire N__12551;
    wire N__12546;
    wire N__12541;
    wire N__12538;
    wire N__12537;
    wire N__12536;
    wire N__12533;
    wire N__12528;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12511;
    wire N__12510;
    wire N__12509;
    wire N__12506;
    wire N__12501;
    wire N__12496;
    wire N__12493;
    wire N__12490;
    wire N__12487;
    wire N__12484;
    wire N__12481;
    wire N__12478;
    wire N__12475;
    wire N__12472;
    wire N__12469;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12457;
    wire N__12454;
    wire N__12451;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12439;
    wire N__12436;
    wire N__12433;
    wire N__12432;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12420;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12382;
    wire N__12379;
    wire N__12376;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12358;
    wire N__12355;
    wire N__12354;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12277;
    wire N__12276;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12243;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12139;
    wire N__12136;
    wire N__12133;
    wire N__12130;
    wire N__12127;
    wire N__12124;
    wire N__12121;
    wire N__12118;
    wire N__12115;
    wire N__12112;
    wire N__12109;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_21_0_;
    wire \c0.tx.n4414 ;
    wire \c0.tx.n4415 ;
    wire \c0.tx.n4416 ;
    wire \c0.tx.n4417 ;
    wire \c0.tx.n4418 ;
    wire \c0.tx.n4419 ;
    wire \c0.tx.n4420 ;
    wire \c0.tx.n4421 ;
    wire bfn_1_22_0_;
    wire n5037_cascade_;
    wire n3611;
    wire n4_adj_2008_cascade_;
    wire \c0.tx2.n5312_cascade_ ;
    wire \c0.n5815_cascade_ ;
    wire \c0.n5818 ;
    wire \c0.tx2.n5932_cascade_ ;
    wire \c0.n5917_cascade_ ;
    wire \c0.n5920_cascade_ ;
    wire \c0.n5662 ;
    wire \c0.tx2.r_Tx_Data_7 ;
    wire \c0.tx2.n5929 ;
    wire \c0.tx2.r_Tx_Data_6 ;
    wire \c0.tx2.r_Tx_Data_5 ;
    wire \c0.n5399_cascade_ ;
    wire \c0.n5857_cascade_ ;
    wire \c0.n5860 ;
    wire \c0.tx2.o_Tx_Serial_N_1798 ;
    wire n3_cascade_;
    wire \c0.data_in_frame_19_0 ;
    wire tx2_o;
    wire tx2_enable;
    wire \c0.n5402 ;
    wire \c0.data_in_frame_19_3 ;
    wire \c0.n5863 ;
    wire bfn_1_30_0_;
    wire \c0.rx.n4422 ;
    wire \c0.rx.n4423 ;
    wire \c0.rx.n4424 ;
    wire \c0.rx.n4425 ;
    wire \c0.rx.n4426 ;
    wire \c0.rx.n4427 ;
    wire \c0.rx.n4428 ;
    wire n2156_cascade_;
    wire n8;
    wire \c0.rx.n5298_cascade_ ;
    wire \c0.rx.n5536 ;
    wire \c0.rx.n5049 ;
    wire n5050;
    wire \c0.rx.n5923_cascade_ ;
    wire \c0.rx.n5926_cascade_ ;
    wire \c0.rx.n5537 ;
    wire n5490;
    wire \c0.rx.n3980_cascade_ ;
    wire \c0.rx.n5532 ;
    wire bfn_2_17_0_;
    wire \c0.n4378 ;
    wire \c0.tx_transmit_N_568_2 ;
    wire \c0.n4379 ;
    wire \c0.tx_transmit_N_568_3 ;
    wire \c0.n4380 ;
    wire \c0.n4381 ;
    wire \c0.byte_transmit_counter_5 ;
    wire \c0.n4382 ;
    wire \c0.byte_transmit_counter_6 ;
    wire \c0.n4383 ;
    wire \c0.byte_transmit_counter_7 ;
    wire \c0.n4384 ;
    wire \c0.n50 ;
    wire \c0.tx_active_prev ;
    wire \c0.n5540_cascade_ ;
    wire \c0.n5977_cascade_ ;
    wire n1760_cascade_;
    wire n1760;
    wire \c0.n1529_cascade_ ;
    wire \c0.n1801 ;
    wire \c0.tx.n315 ;
    wire n319;
    wire \c0.tx.n320 ;
    wire \c0.tx.n321 ;
    wire \c0.tx.r_Clock_Count_0 ;
    wire \c0.tx.n313 ;
    wire n316;
    wire n314;
    wire n317;
    wire r_Clock_Count_2;
    wire \c0.tx.r_Clock_Count_6 ;
    wire \c0.tx.r_Clock_Count_1 ;
    wire r_Clock_Count_5;
    wire r_Clock_Count_4;
    wire \c0.tx.n5_cascade_ ;
    wire r_Clock_Count_7;
    wire n3595_cascade_;
    wire \c0.tx.n5520 ;
    wire \c0.tx.r_Clock_Count_3 ;
    wire \c0.tx2.n5_cascade_ ;
    wire \c0.tx2.n3591 ;
    wire \c0.tx2.n3591_cascade_ ;
    wire r_SM_Main_2_N_1767_1_cascade_;
    wire \c0.tx2.r_Clock_Count_0 ;
    wire n2460;
    wire bfn_2_23_0_;
    wire \c0.tx2.r_Clock_Count_1 ;
    wire n2399;
    wire \c0.tx2.n4429 ;
    wire \c0.tx2.n4430 ;
    wire \c0.tx2.n4431 ;
    wire \c0.tx2.r_Clock_Count_4 ;
    wire n2382;
    wire \c0.tx2.n4432 ;
    wire \c0.tx2.r_Clock_Count_5 ;
    wire n2379;
    wire \c0.tx2.n4433 ;
    wire \c0.tx2.r_Clock_Count_6 ;
    wire n2376;
    wire \c0.tx2.n4434 ;
    wire \c0.tx2.n4435 ;
    wire \c0.tx2.n4436 ;
    wire r_Clock_Count_8_adj_2012;
    wire bfn_2_24_0_;
    wire n2369;
    wire \c0.tx2.r_Tx_Data_0 ;
    wire \c0.tx2.n5947 ;
    wire \c0.tx2.n5950 ;
    wire n1345;
    wire \c0.tx2.r_Tx_Data_4 ;
    wire \c0.tx2.r_Tx_Data_2 ;
    wire \c0.tx2.r_Tx_Data_3 ;
    wire \c0.n5665_cascade_ ;
    wire \c0.n5372_cascade_ ;
    wire \c0.n5659 ;
    wire \c0.n5938 ;
    wire \c0.n5971_cascade_ ;
    wire \c0.n5725_cascade_ ;
    wire \c0.n1058 ;
    wire \c0.n5728_cascade_ ;
    wire \c0.n5974 ;
    wire \c0.tx2.r_Tx_Data_1 ;
    wire \c0.tx2.n1592 ;
    wire \c0.n5803_cascade_ ;
    wire \c0.data_in_frame_18_1 ;
    wire \c0.n5369 ;
    wire \c0.n5869 ;
    wire \c0.n5959 ;
    wire \c0.n5962 ;
    wire \c0.data_in_frame_18_3 ;
    wire n5051;
    wire n5491;
    wire \c0.rx.n5535 ;
    wire \c0.rx.n2157 ;
    wire \c0.rx.n5538 ;
    wire \c0.rx.n5539 ;
    wire \c0.rx.n40 ;
    wire \c0.rx.r_SM_Main_2_N_1824_2_cascade_ ;
    wire n4474;
    wire n2156;
    wire n4474_cascade_;
    wire \c0.rx.n4_adj_1866_cascade_ ;
    wire \c0.rx.n4011 ;
    wire data_in_5_1;
    wire \c0.rx.r_Clock_Count_5 ;
    wire \c0.rx.r_Clock_Count_4 ;
    wire \c0.rx.n37 ;
    wire \c0.rx.r_Clock_Count_1 ;
    wire \c0.rx.n37_cascade_ ;
    wire \c0.rx.r_Clock_Count_3 ;
    wire r_SM_Main_2_N_1830_0;
    wire \c0.rx.r_Rx_Data_R ;
    wire n12_adj_1995_cascade_;
    wire n5316;
    wire n16_adj_1993;
    wire \c0.rx.n3573 ;
    wire \c0.rx.n3573_cascade_ ;
    wire \c0.n20_adj_1918_cascade_ ;
    wire \c0.n87 ;
    wire \c0.n87_cascade_ ;
    wire \c0.n16_adj_1909 ;
    wire \c0.tx_transmit_N_568_5 ;
    wire \c0.tx_transmit_N_568_6 ;
    wire \c0.tx_transmit_N_568_7 ;
    wire \c0.tx_transmit_N_568_4 ;
    wire \c0.n103 ;
    wire \c0.n109 ;
    wire \c0.n45 ;
    wire \c0.n109_cascade_ ;
    wire n4315_cascade_;
    wire n4316_cascade_;
    wire n7_adj_2002;
    wire n5066;
    wire tx_active;
    wire data_out_19_4;
    wire data_out_18_4;
    wire \c0.n17_cascade_ ;
    wire tx_data_4_N_keep_cascade_;
    wire n8_adj_2001;
    wire \c0.tx.r_SM_Main_2_N_1767_1_cascade_ ;
    wire n5041;
    wire \c0.tx_transmit ;
    wire \c0.tx.n12_cascade_ ;
    wire r_Clock_Count_8;
    wire n1307_cascade_;
    wire n3595;
    wire n4221;
    wire n2;
    wire n1307;
    wire n4_adj_2003_cascade_;
    wire n4155;
    wire n2372;
    wire \c0.tx2.r_Clock_Count_7 ;
    wire n2395;
    wire \c0.tx2.r_Clock_Count_2 ;
    wire r_SM_Main_0_adj_2011;
    wire r_SM_Main_2_N_1767_1;
    wire r_SM_Main_1_adj_2010;
    wire \c0.tx2.n2218_cascade_ ;
    wire \c0.tx2.n3577 ;
    wire \c0.n5953 ;
    wire \c0.n5956 ;
    wire n2392;
    wire r_SM_Main_2_adj_2009;
    wire n5037;
    wire \c0.tx2.r_Clock_Count_3 ;
    wire bfn_3_24_0_;
    wire \c0.n4400 ;
    wire \c0.n4401 ;
    wire \c0.n4402 ;
    wire \c0.n4403 ;
    wire \c0.byte_transmit_counter2_4 ;
    wire \c0.n5785_cascade_ ;
    wire \c0.n5426 ;
    wire \c0.n5788 ;
    wire \c0.n5968 ;
    wire \c0.n5363 ;
    wire \c0.data_in_frame_19_7 ;
    wire \c0.n5935 ;
    wire \c0.n5944 ;
    wire \c0.data_in_frame_19_6 ;
    wire \c0.n5456 ;
    wire data_in_18_3;
    wire \c0.n1893_cascade_ ;
    wire \c0.n20_adj_1921 ;
    wire \c0.n5459 ;
    wire \c0.n5737 ;
    wire \c0.data_in_frame_19_1 ;
    wire \c0.data_in_field_131 ;
    wire \c0.n2036_cascade_ ;
    wire \c0.n5273_cascade_ ;
    wire \c0.data_in_frame_18_7 ;
    wire \c0.n5671 ;
    wire rx_data_3;
    wire rx_data_5;
    wire r_Clock_Count_7_adj_2004;
    wire \c0.rx.r_Clock_Count_2 ;
    wire \c0.rx.n6 ;
    wire \c0.rx.n2213 ;
    wire \c0.rx.n2317 ;
    wire \c0.rx.r_Bit_Index_1 ;
    wire \c0.rx.r_Bit_Index_2 ;
    wire r_Clock_Count_0;
    wire r_Clock_Count_6;
    wire n8_adj_1996;
    wire tx_enable;
    wire bfn_4_16_0_;
    wire \c0.delay_counter_1 ;
    wire \c0.n4404 ;
    wire \c0.n4405 ;
    wire \c0.delay_counter_3 ;
    wire \c0.n4406 ;
    wire \c0.delay_counter_4 ;
    wire \c0.n4407 ;
    wire \c0.delay_counter_5 ;
    wire \c0.n4408 ;
    wire \c0.delay_counter_6 ;
    wire \c0.n4409 ;
    wire \c0.n4410 ;
    wire \c0.n4411 ;
    wire \c0.delay_counter_8 ;
    wire bfn_4_17_0_;
    wire \c0.n4412 ;
    wire \c0.n4413 ;
    wire \c0.delay_counter_10 ;
    wire n5077;
    wire n4_adj_1988;
    wire data_out_19_0;
    wire \c0.delay_counter_9 ;
    wire \c0.delay_counter_2 ;
    wire \c0.delay_counter_0 ;
    wire \c0.delay_counter_7 ;
    wire \c0.n18_adj_1908 ;
    wire n4_adj_2000;
    wire n5086_cascade_;
    wire n1525;
    wire n5156_cascade_;
    wire data_out_18_0;
    wire n5156;
    wire n5063;
    wire data_out_18_3;
    wire data_out_19_7;
    wire n7_adj_1998;
    wire n8_adj_1997;
    wire data_out_18_7;
    wire data_out_19_3;
    wire data_out_18_1;
    wire n4_adj_2007;
    wire r_Tx_Data_1;
    wire \c0.n9 ;
    wire \c0.n5501 ;
    wire \c0.n1173_cascade_ ;
    wire tx_data_0_N_keep_cascade_;
    wire r_Tx_Data_0;
    wire \c0.n5531 ;
    wire \c0.n15_cascade_ ;
    wire tx_data_1_N_keep;
    wire \c0.tx.r_SM_Main_2_N_1767_1 ;
    wire \c0.tx.n3507 ;
    wire \c0.tx.n3507_cascade_ ;
    wire n2307;
    wire n2200;
    wire n2307_cascade_;
    wire n805;
    wire \c0.tx2.r_Bit_Index_0 ;
    wire \c0.tx2.r_Bit_Index_1 ;
    wire \c0.tx2.r_Bit_Index_2 ;
    wire \c0.tx2.n2218 ;
    wire \c0.tx2.n2319 ;
    wire n5153;
    wire \c0.n3414_cascade_ ;
    wire \c0.n3414 ;
    wire \c0.FRAME_MATCHER_wait_for_transmission_N_909 ;
    wire \c0.r_SM_Main_2_N_1770_0 ;
    wire tx2_active;
    wire \c0.n195 ;
    wire \c0.n5845_cascade_ ;
    wire \c0.n2275 ;
    wire \c0.data_in_field_81 ;
    wire \c0.n1918_cascade_ ;
    wire \c0.n5192_cascade_ ;
    wire \c0.n30_adj_1897_cascade_ ;
    wire \c0.n36_cascade_ ;
    wire \c0.n5080_cascade_ ;
    wire \c0.n1990 ;
    wire \c0.n5192 ;
    wire \c0.n5080 ;
    wire \c0.n23_adj_1931 ;
    wire \c0.n21_adj_1928 ;
    wire \c0.n22_adj_1927_cascade_ ;
    wire \c0.n24_adj_1907 ;
    wire data_in_19_3;
    wire \c0.data_in_frame_18_0 ;
    wire \c0.data_in_frame_18_4 ;
    wire \c0.n22_adj_1881 ;
    wire \c0.n5266 ;
    wire \c0.data_in_field_101 ;
    wire \c0.n18_adj_1882_cascade_ ;
    wire \c0.n26_adj_1883 ;
    wire \c0.n5462 ;
    wire data_in_12_5;
    wire \c0.n5222_cascade_ ;
    wire \c0.n42 ;
    wire \c0.n33_cascade_ ;
    wire \c0.n2008_cascade_ ;
    wire \c0.n38_cascade_ ;
    wire \c0.data_in_frame_18_6 ;
    wire data_in_2_5;
    wire rx_data_6;
    wire \c0.rx.n2151_cascade_ ;
    wire n1709_cascade_;
    wire n4_adj_1990;
    wire rx_data_4;
    wire n4_adj_1992;
    wire data_out_11_0;
    wire data_out_18_2;
    wire data_out_19_2;
    wire \c0.n2249 ;
    wire \c0.n5522_cascade_ ;
    wire n4_adj_1991;
    wire data_out_18_5;
    wire n4_adj_1994;
    wire n5135;
    wire n5117;
    wire n5117_cascade_;
    wire n4316;
    wire data_out_19_5;
    wire tx_data_2_N_keep;
    wire data_out_11_3;
    wire data_out_11_2;
    wire \c0.n1805_cascade_ ;
    wire n135;
    wire \c0.n1805 ;
    wire n5173;
    wire data_out_11_7;
    wire data_out_10_7;
    wire n5079;
    wire data_out_19_1;
    wire \c0.n5519 ;
    wire \c0.n5980 ;
    wire r_Tx_Data_4;
    wire \c0.tx.n5713_cascade_ ;
    wire data_out_11_1;
    wire \c0.n9_adj_1880 ;
    wire \c0.n9_adj_1890 ;
    wire \c0.n5489 ;
    wire \c0.n991_cascade_ ;
    wire tx_data_5_N_keep_cascade_;
    wire r_Tx_Data_5;
    wire tx_data_3_N_keep;
    wire r_Tx_Data_3;
    wire r_Tx_Data_2;
    wire r_Bit_Index_1;
    wire r_Bit_Index_0;
    wire \c0.tx.n5719 ;
    wire r_Bit_Index_2;
    wire \c0.tx.n5716 ;
    wire \c0.tx.n5722 ;
    wire r_SM_Main_1;
    wire \c0.tx.o_Tx_Serial_N_1798_cascade_ ;
    wire r_SM_Main_0;
    wire r_SM_Main_2;
    wire \c0.tx.n3_cascade_ ;
    wire tx_o;
    wire \c0.n2018 ;
    wire \c0.data_in_frame_18_2 ;
    wire \c0.n5965 ;
    wire data_in_19_6;
    wire \c0.n22_adj_1901_cascade_ ;
    wire \c0.n23_adj_1932 ;
    wire \c0.n30_adj_1940_cascade_ ;
    wire \c0.n3563 ;
    wire \c0.n5280 ;
    wire \c0.n5277 ;
    wire \c0.n25_adj_1941 ;
    wire \c0.n5072 ;
    wire \c0.n26_adj_1915_cascade_ ;
    wire data_in_17_3;
    wire \c0.data_in_field_71 ;
    wire \c0.n26_cascade_ ;
    wire \c0.n27_adj_1919 ;
    wire \c0.n5250 ;
    wire \c0.n28_adj_1917_cascade_ ;
    wire \c0.n26_adj_1939 ;
    wire \c0.data_in_field_41 ;
    wire \c0.n14_cascade_ ;
    wire \c0.n15_adj_1894 ;
    wire \c0.n16_adj_1893_cascade_ ;
    wire \c0.n22_adj_1930 ;
    wire \c0.n2058 ;
    wire \c0.n5096_cascade_ ;
    wire \c0.n1785_cascade_ ;
    wire \c0.n22 ;
    wire data_in_13_5;
    wire \c0.n5150 ;
    wire \c0.data_in_field_109 ;
    wire \c0.n39 ;
    wire \c0.n45_adj_1885 ;
    wire \c0.n43 ;
    wire \c0.n30 ;
    wire \c0.n5275_cascade_ ;
    wire \c0.n24_adj_1929 ;
    wire \c0.n5182 ;
    wire \c0.n5147 ;
    wire \c0.n5182_cascade_ ;
    wire \c0.n40 ;
    wire \c0.data_in_field_119 ;
    wire \c0.n29 ;
    wire \c0.n20_adj_1906 ;
    wire data_in_4_3;
    wire data_in_16_6;
    wire \c0.n5731 ;
    wire \c0.n5264 ;
    wire \c0.n5264_cascade_ ;
    wire data_in_19_1;
    wire data_in_2_3;
    wire r_SM_Main_2_adj_2005;
    wire \c0.rx.r_SM_Main_1 ;
    wire \c0.rx.n5058 ;
    wire \c0.rx.r_Bit_Index_0 ;
    wire r_SM_Main_0_adj_2006;
    wire \c0.rx.n5058_cascade_ ;
    wire \c0.rx.r_SM_Main_2_N_1824_2 ;
    wire n4;
    wire n1714_cascade_;
    wire rx_data_1;
    wire data_in_0_7;
    wire n4_adj_1986;
    wire n1709;
    wire data_0;
    wire bfn_6_17_0_;
    wire data_1;
    wire \c0.n4385 ;
    wire data_2;
    wire \c0.n4386 ;
    wire data_3;
    wire \c0.n4387 ;
    wire \c0.n4388 ;
    wire data_5;
    wire \c0.n4389 ;
    wire data_6;
    wire \c0.n4390 ;
    wire data_7;
    wire \c0.n4391 ;
    wire \c0.n4392 ;
    wire bfn_6_18_0_;
    wire data_9;
    wire \c0.n4393 ;
    wire \c0.n4394 ;
    wire data_11;
    wire \c0.n4395 ;
    wire data_12;
    wire \c0.n4396 ;
    wire data_13;
    wire \c0.n4397 ;
    wire \c0.n4398 ;
    wire \c0.n4399 ;
    wire data_15;
    wire data_4;
    wire data_14;
    wire data_out_11_4;
    wire data_out_10_4;
    wire \c0.n9_adj_1887_cascade_ ;
    wire \c0.n15_adj_1889 ;
    wire data_8;
    wire \c0.n17_adj_1961 ;
    wire \c0.n1236_cascade_ ;
    wire \c0.n2247 ;
    wire \c0.n1227 ;
    wire \c0.n5511_cascade_ ;
    wire tx_data_7_N_keep_cascade_;
    wire r_Tx_Data_7;
    wire n1442;
    wire r_Tx_Data_6;
    wire data_out_10_0;
    wire n1748;
    wire n21_adj_1999;
    wire data_10;
    wire n4315;
    wire data_out_10_2;
    wire \c0.n5411 ;
    wire \c0.n5830 ;
    wire \c0.n5941 ;
    wire \c0.data_in_frame_19_2 ;
    wire \c0.data_in_frame_18_5 ;
    wire \c0.data_in_frame_19_5 ;
    wire data_in_14_5;
    wire \c0.n5809 ;
    wire \c0.n5241 ;
    wire \c0.tx2_transmit_N_1031_cascade_ ;
    wire \c0.n38_adj_1934 ;
    wire \c0.n14_adj_1900 ;
    wire data_in_15_0;
    wire \c0.n5210 ;
    wire \c0.tx2_transmit_N_1031 ;
    wire \c0.n1785 ;
    wire \c0.n11 ;
    wire \c0.n24_adj_1924 ;
    wire \c0.n5259_cascade_ ;
    wire \c0.n21_adj_1933 ;
    wire \c0.n16 ;
    wire \c0.n1893 ;
    wire \c0.n2008 ;
    wire \c0.n5225 ;
    wire \c0.n5198_cascade_ ;
    wire \c0.n6103 ;
    wire \c0.n28 ;
    wire \c0.n5198 ;
    wire \c0.n1918 ;
    wire \c0.n18_adj_1910 ;
    wire \c0.n17_adj_1912_cascade_ ;
    wire \c0.n12_adj_1911 ;
    wire \c0.n19_adj_1920 ;
    wire \c0.n28_adj_1902 ;
    wire \c0.n32 ;
    wire \c0.n29_adj_1905_cascade_ ;
    wire \c0.n31_adj_1904 ;
    wire \c0.n5278 ;
    wire \c0.data_in_field_134 ;
    wire \c0.n12_cascade_ ;
    wire \c0.n1880 ;
    wire \c0.n2036 ;
    wire \c0.n20_adj_1892 ;
    wire \c0.n2033 ;
    wire \c0.n10_adj_1963_cascade_ ;
    wire \c0.n5114 ;
    wire \c0.n5114_cascade_ ;
    wire \c0.n30_adj_1903 ;
    wire \c0.n5743 ;
    wire \c0.data_in_field_87 ;
    wire \c0.data_in_field_57 ;
    wire \c0.data_in_field_7 ;
    wire \c0.n5162_cascade_ ;
    wire data_in_18_1;
    wire \c0.n1825_cascade_ ;
    wire \c0.data_in_field_133 ;
    wire \c0.data_in_field_73 ;
    wire \c0.data_in_field_35 ;
    wire \c0.n18 ;
    wire \c0.data_in_field_137 ;
    wire \c0.n6_adj_1877 ;
    wire \c0.data_in_field_31 ;
    wire \c0.n28_adj_1886 ;
    wire \c0.n5222 ;
    wire \c0.n34 ;
    wire data_in_15_5;
    wire \c0.n1686_cascade_ ;
    wire \c0.data_in_field_25 ;
    wire data_in_19_7;
    wire r_Rx_Data;
    wire n1714;
    wire n3342;
    wire rx_data_7;
    wire data_in_17_1;
    wire data_out_19_6;
    wire data_out_18_6;
    wire data_out_11_5;
    wire n5176;
    wire \c0.n1590 ;
    wire data_out_11_6;
    wire \c0.byte_transmit_counter_1 ;
    wire data_out_10_6;
    wire \c0.byte_transmit_counter_0 ;
    wire \c0.n3567 ;
    wire \c0.byte_transmit_counter_3 ;
    wire \c0.n5523_cascade_ ;
    wire \c0.byte_transmit_counter_2 ;
    wire \c0.n1236 ;
    wire \c0.n5515 ;
    wire \c0.n5513_cascade_ ;
    wire \c0.byte_transmit_counter_4 ;
    wire tx_data_6_N_keep;
    wire data_out_10_5;
    wire data_out_10_1;
    wire data_out_10_3;
    wire n5132;
    wire \c0.n5839_cascade_ ;
    wire \c0.n5833_cascade_ ;
    wire \c0.n5417_cascade_ ;
    wire \c0.n5414 ;
    wire \c0.n5827 ;
    wire \c0.n5683_cascade_ ;
    wire \c0.n5695 ;
    wire \c0.n5480_cascade_ ;
    wire \c0.n5483 ;
    wire \c0.n5677_cascade_ ;
    wire \c0.n5680 ;
    wire data_in_18_5;
    wire \c0.n24_adj_1895 ;
    wire rx_data_0;
    wire data_in_19_0;
    wire \c0.n5429 ;
    wire \c0.n5791 ;
    wire \c0.n5432 ;
    wire \c0.data_in_field_30 ;
    wire \c0.data_in_field_13 ;
    wire \c0.n5393 ;
    wire data_in_14_7;
    wire \c0.n10_adj_1898 ;
    wire \c0.data_in_field_69 ;
    wire \c0.n5159 ;
    wire \c0.data_in_field_99 ;
    wire \c0.n5159_cascade_ ;
    wire \c0.data_in_field_105 ;
    wire \c0.n2095_cascade_ ;
    wire \c0.n1821 ;
    wire \c0.n34_adj_1896 ;
    wire \c0.data_in_field_11 ;
    wire \c0.n5821_cascade_ ;
    wire \c0.n5423 ;
    wire \c0.data_in_field_27 ;
    wire \c0.n2080 ;
    wire \c0.n2080_cascade_ ;
    wire \c0.n5243 ;
    wire \c0.n16_adj_1922 ;
    wire \c0.n25_adj_1926 ;
    wire \c0.n1978 ;
    wire \c0.n5261 ;
    wire \c0.n5689_cascade_ ;
    wire \c0.n5366 ;
    wire \c0.n14_adj_1967 ;
    wire \c0.n5276 ;
    wire \c0.n5201 ;
    wire \c0.n5276_cascade_ ;
    wire \c0.n37 ;
    wire \c0.data_in_field_36 ;
    wire \c0.data_in_field_22 ;
    wire \c0.n2005_cascade_ ;
    wire \c0.n10_adj_1873_cascade_ ;
    wire \c0.n1825 ;
    wire \c0.data_in_field_55 ;
    wire \c0.n13_adj_1951 ;
    wire \c0.data_in_field_23 ;
    wire \c0.n6107 ;
    wire \c0.n18_adj_1891 ;
    wire \c0.n5249 ;
    wire rx_data_2;
    wire \c0.n5255 ;
    wire data_in_1_3;
    wire \c0.n28_adj_1954 ;
    wire \c0.n26_adj_1955 ;
    wire \c0.n25_adj_1957_cascade_ ;
    wire \c0.n4465 ;
    wire \c0.data_in_field_17 ;
    wire data_in_1_4;
    wire data_in_11_7;
    wire data_in_10_7;
    wire data_in_2_7;
    wire \c0.n27_adj_1956 ;
    wire \c0.n26_adj_1958 ;
    wire \c0.data_in_field_135 ;
    wire \c0.data_in_field_113 ;
    wire \c0.n1772 ;
    wire \c0.n5144 ;
    wire \c0.n5144_cascade_ ;
    wire \c0.n31 ;
    wire data_in_8_5;
    wire data_in_8_7;
    wire \c0.n5447_cascade_ ;
    wire \c0.n5755_cascade_ ;
    wire \c0.n5758 ;
    wire \c0.data_in_field_54 ;
    wire \c0.data_in_field_10 ;
    wire \c0.n5438 ;
    wire \c0.data_in_field_82 ;
    wire \c0.n5767_cascade_ ;
    wire \c0.n5444 ;
    wire \c0.n5761 ;
    wire \c0.n13 ;
    wire \c0.data_in_field_117 ;
    wire \c0.n2074_cascade_ ;
    wire \c0.n10_adj_1888 ;
    wire \c0.data_in_field_95 ;
    wire \c0.n1851 ;
    wire \c0.data_in_field_96 ;
    wire \c0.n5099 ;
    wire \c0.n5162 ;
    wire \c0.n5213 ;
    wire \c0.n5099_cascade_ ;
    wire \c0.n19 ;
    wire \c0.data_in_field_104 ;
    wire data_in_0_6;
    wire data_in_12_0;
    wire \c0.data_in_field_89 ;
    wire \c0.data_in_field_120 ;
    wire \c0.n23_adj_1925 ;
    wire \c0.data_in_field_83 ;
    wire \c0.n5797 ;
    wire \c0.data_in_field_19 ;
    wire \c0.n23 ;
    wire data_in_3_3;
    wire \c0.n25_adj_1960 ;
    wire \c0.data_in_field_67 ;
    wire \c0.n5093 ;
    wire \c0.data_in_field_21 ;
    wire \c0.n5881 ;
    wire data_in_15_6;
    wire \c0.data_in_field_29 ;
    wire \c0.n2046 ;
    wire \c0.data_in_field_85 ;
    wire \c0.n2046_cascade_ ;
    wire \c0.n5108 ;
    wire data_in_7_1;
    wire data_in_6_1;
    wire \c0.data_in_field_141 ;
    wire data_in_1_6;
    wire data_in_9_7;
    wire data_in_6_7;
    wire data_in_3_1;
    wire data_in_7_5;
    wire data_in_18_6;
    wire data_in_17_6;
    wire data_in_1_5;
    wire data_in_7_7;
    wire \c0.data_in_field_121 ;
    wire data_in_3_7;
    wire data_in_17_5;
    wire data_in_16_5;
    wire data_in_19_2;
    wire \c0.n5779 ;
    wire data_in_13_0;
    wire data_in_14_0;
    wire \c0.n1929 ;
    wire \c0.data_in_field_112 ;
    wire \c0.n1929_cascade_ ;
    wire \c0.n10_adj_1870_cascade_ ;
    wire \c0.n5204 ;
    wire \c0.data_in_field_28 ;
    wire \c0.data_in_field_20 ;
    wire \c0.data_in_field_12 ;
    wire \c0.n5851_cascade_ ;
    wire \c0.n5408 ;
    wire \c0.n5267 ;
    wire \c0.n5905 ;
    wire \c0.n2074 ;
    wire data_in_19_5;
    wire \c0.n22_adj_1914 ;
    wire \c0.data_in_field_139 ;
    wire \c0.n1947_cascade_ ;
    wire \c0.n10 ;
    wire \c0.data_in_field_51 ;
    wire \c0.n1922 ;
    wire \c0.data_in_field_75 ;
    wire \c0.n5474 ;
    wire \c0.n26_adj_1884 ;
    wire \c0.data_in_field_98 ;
    wire data_in_12_7;
    wire \c0.data_in_field_103 ;
    wire \c0.data_in_field_61 ;
    wire \c0.n5875_cascade_ ;
    wire \c0.data_in_field_37 ;
    wire \c0.n5396 ;
    wire \c0.data_in_field_53 ;
    wire \c0.data_in_field_88 ;
    wire \c0.data_in_field_124 ;
    wire \c0.n1944 ;
    wire \c0.n1944_cascade_ ;
    wire \c0.n20_cascade_ ;
    wire \c0.data_in_field_43 ;
    wire \c0.n24 ;
    wire data_in_4_7;
    wire \c0.data_in_field_39 ;
    wire \c0.data_in_field_5 ;
    wire \c0.data_in_field_79 ;
    wire \c0.data_in_field_77 ;
    wire \c0.n10_adj_1871_cascade_ ;
    wire \c0.n5234 ;
    wire \c0.n1975 ;
    wire \c0.data_in_field_38 ;
    wire data_in_12_1;
    wire \c0.n2062 ;
    wire \c0.n1830 ;
    wire \c0.n5141 ;
    wire \c0.data_in_field_106 ;
    wire data_in_13_7;
    wire \c0.data_in_field_111 ;
    wire \c0.data_in_field_143 ;
    wire data_in_16_7;
    wire data_in_18_7;
    wire data_in_17_7;
    wire \c0.data_in_field_49 ;
    wire \c0.n2092_cascade_ ;
    wire \c0.n2043 ;
    wire \c0.n5246 ;
    wire data_in_0_2;
    wire \c0.data_in_field_9 ;
    wire \c0.n5749 ;
    wire \c0.data_in_field_1 ;
    wire \c0.n5453 ;
    wire \c0.data_in_field_59 ;
    wire data_in_6_6;
    wire data_in_13_4;
    wire data_in_2_4;
    wire \c0.data_in_field_115 ;
    wire data_in_9_1;
    wire data_in_7_6;
    wire data_in_10_4;
    wire data_in_10_3;
    wire data_in_9_3;
    wire \c0.n26_adj_1878 ;
    wire data_in_0_4;
    wire \c0.data_in_field_68 ;
    wire \c0.n5105 ;
    wire \c0.n5111 ;
    wire \c0.n35 ;
    wire data_in_16_3;
    wire data_in_18_4;
    wire data_in_17_4;
    wire \c0.data_in_field_63 ;
    wire \c0.data_in_field_62 ;
    wire \c0.n1795_cascade_ ;
    wire \c0.n6097 ;
    wire data_in_6_3;
    wire data_in_5_3;
    wire \c0.data_in_field_142 ;
    wire \c0.n1795 ;
    wire \c0.n11_adj_1913 ;
    wire data_in_11_4;
    wire \c0.data_in_field_92 ;
    wire data_in_11_5;
    wire \c0.data_in_field_93 ;
    wire \c0.n5707 ;
    wire \c0.n1838 ;
    wire data_in_5_0;
    wire \c0.n6_adj_1876_cascade_ ;
    wire \c0.data_in_field_132 ;
    wire \c0.n5129 ;
    wire \c0.n6_adj_1874 ;
    wire data_in_0_0;
    wire \c0.data_in_field_0 ;
    wire \c0.data_in_field_90 ;
    wire \c0.n22_adj_1935 ;
    wire data_in_5_6;
    wire \c0.data_in_field_2 ;
    wire \c0.data_in_field_108 ;
    wire \c0.n5102 ;
    wire data_in_5_7;
    wire \c0.data_in_field_47 ;
    wire data_in_15_7;
    wire \c0.data_in_field_127 ;
    wire data_in_16_0;
    wire data_in_1_7;
    wire data_in_10_5;
    wire data_in_9_5;
    wire data_in_0_5;
    wire data_in_1_2;
    wire data_in_6_5;
    wire data_in_4_6;
    wire data_in_6_0;
    wire \c0.data_in_field_60 ;
    wire \c0.n6_adj_1875 ;
    wire data_in_3_5;
    wire data_in_3_4;
    wire data_in_2_6;
    wire data_in_3_6;
    wire \c0.n28_adj_1953_cascade_ ;
    wire \c0.n22_adj_1952 ;
    wire \c0.n30_adj_1959 ;
    wire data_in_4_5;
    wire data_in_8_0;
    wire \c0.data_in_field_58 ;
    wire \c0.n5773_cascade_ ;
    wire \c0.data_in_field_34 ;
    wire \c0.n5441 ;
    wire \c0.n5477 ;
    wire data_in_16_4;
    wire data_in_15_4;
    wire data_in_8_6;
    wire data_in_11_1;
    wire data_in_10_1;
    wire data_in_11_0;
    wire \c0.data_in_field_14 ;
    wire \c0.n5911 ;
    wire \c0.data_in_field_6 ;
    wire \c0.data_in_field_138 ;
    wire \c0.data_in_field_130 ;
    wire \c0.n5123 ;
    wire \c0.n5123_cascade_ ;
    wire \c0.n5231 ;
    wire data_in_13_2;
    wire data_in_12_2;
    wire \c0.data_in_field_64 ;
    wire \c0.n5179 ;
    wire \c0.data_in_field_46 ;
    wire \c0.data_in_field_4 ;
    wire \c0.n1767_cascade_ ;
    wire \c0.n1899 ;
    wire \c0.n5126 ;
    wire \c0.data_in_field_140 ;
    wire \c0.n5126_cascade_ ;
    wire \c0.data_in_field_125 ;
    wire \c0.n20_adj_1899 ;
    wire data_in_14_6;
    wire \c0.n10_adj_1872 ;
    wire data_in_12_4;
    wire \c0.data_in_field_100 ;
    wire \c0.data_in_field_40 ;
    wire \c0.data_in_field_128 ;
    wire \c0.data_in_field_16 ;
    wire \c0.data_in_field_72 ;
    wire \c0.n5188 ;
    wire \c0.n5138_cascade_ ;
    wire \c0.n15_adj_1968 ;
    wire data_in_3_2;
    wire \c0.data_in_field_26 ;
    wire data_in_4_1;
    wire \c0.data_in_field_33 ;
    wire data_in_2_2;
    wire \c0.data_in_field_18 ;
    wire \c0.n6 ;
    wire data_in_4_0;
    wire \c0.data_in_field_32 ;
    wire data_in_13_6;
    wire n5332;
    wire n5331_cascade_;
    wire LED_c;
    wire \c0.data_in_field_97 ;
    wire \c0.n1972 ;
    wire data_in_9_4;
    wire \c0.data_in_field_76 ;
    wire data_in_0_1;
    wire data_in_5_5;
    wire \c0.data_in_field_45 ;
    wire data_in_9_0;
    wire data_in_2_1;
    wire data_in_1_1;
    wire \c0.data_in_field_48 ;
    wire \c0.n5701 ;
    wire data_in_4_4;
    wire data_in_6_4;
    wire data_in_7_2;
    wire data_in_10_6;
    wire data_in_9_6;
    wire data_in_10_0;
    wire \c0.data_in_field_80 ;
    wire data_in_8_2;
    wire data_in_14_2;
    wire \c0.data_in_field_114 ;
    wire data_in_4_2;
    wire \c0.data_in_field_66 ;
    wire \c0.data_in_field_84 ;
    wire \c0.n1969 ;
    wire \c0.n25 ;
    wire data_in_5_2;
    wire \c0.data_in_field_42 ;
    wire \c0.data_in_field_107 ;
    wire \c0.data_in_field_15 ;
    wire \c0.n20_adj_1916 ;
    wire data_in_8_1;
    wire \c0.data_in_field_65 ;
    wire data_in_16_1;
    wire data_in_15_1;
    wire data_in_14_4;
    wire \c0.data_in_field_116 ;
    wire \c0.n1815 ;
    wire \c0.n1815_cascade_ ;
    wire \c0.data_in_field_52 ;
    wire \c0.n27 ;
    wire data_in_14_1;
    wire data_in_13_1;
    wire data_in_7_0;
    wire \c0.data_in_field_56 ;
    wire \c0.data_in_field_129 ;
    wire \c0.n15_adj_1923 ;
    wire data_in_6_2;
    wire \c0.data_in_field_50 ;
    wire \c0.data_in_field_8 ;
    wire data_in_5_4;
    wire \c0.data_in_field_44 ;
    wire \c0.n1962 ;
    wire data_in_3_0;
    wire \c0.data_in_field_24 ;
    wire data_in_2_0;
    wire data_in_1_0;
    wire data_in_15_3;
    wire \c0.data_in_field_123 ;
    wire data_in_12_6;
    wire data_in_11_6;
    wire data_in_18_2;
    wire \c0.data_in_field_74 ;
    wire \c0.data_in_field_136 ;
    wire data_in_15_2;
    wire \c0.data_in_field_122 ;
    wire data_in_14_3;
    wire data_in_13_3;
    wire data_in_12_3;
    wire data_in_11_3;
    wire \c0.data_in_field_91 ;
    wire data_in_0_3;
    wire \c0.data_in_field_3 ;
    wire data_in_11_2;
    wire data_in_10_2;
    wire data_in_9_2;
    wire data_in_8_3;
    wire data_in_7_3;
    wire data_in_18_0;
    wire data_in_17_0;
    wire \c0.data_in_field_118 ;
    wire \c0.data_in_field_126 ;
    wire \c0.byte_transmit_counter2_0 ;
    wire \c0.data_in_field_86 ;
    wire \c0.data_in_field_94 ;
    wire \c0.data_in_field_70 ;
    wire \c0.n5899_cascade_ ;
    wire \c0.data_in_field_78 ;
    wire \c0.n5893 ;
    wire \c0.data_in_field_102 ;
    wire \c0.byte_transmit_counter2_1 ;
    wire \c0.data_in_field_110 ;
    wire \c0.n5384 ;
    wire \c0.n5387_cascade_ ;
    wire \c0.byte_transmit_counter2_2 ;
    wire \c0.n5378 ;
    wire \c0.n5381 ;
    wire \c0.n5887_cascade_ ;
    wire \c0.byte_transmit_counter2_3 ;
    wire \c0.n5890 ;
    wire \c0.n5219 ;
    wire \c0.n5138 ;
    wire \c0.n1896 ;
    wire data_in_8_4;
    wire data_in_7_4;
    wire rx_data_ready;
    wire data_in_17_2;
    wire data_in_16_2;
    wire n26;
    wire bfn_15_25_0_;
    wire n25;
    wire n4437;
    wire n24;
    wire n4438;
    wire n23;
    wire n4439;
    wire n22;
    wire n4440;
    wire n21;
    wire n4441;
    wire n20;
    wire n4442;
    wire n19;
    wire n4443;
    wire n4444;
    wire n18;
    wire bfn_15_26_0_;
    wire n17;
    wire n4445;
    wire n16;
    wire n4446;
    wire n15;
    wire n4447;
    wire n14;
    wire n4448;
    wire n13;
    wire n4449;
    wire n12;
    wire n4450;
    wire n11;
    wire n4451;
    wire n4452;
    wire n10;
    wire bfn_15_27_0_;
    wire n9;
    wire n4453;
    wire n8_adj_1989;
    wire n4454;
    wire n7;
    wire n4455;
    wire n6;
    wire n4456;
    wire blink_counter_21;
    wire n4457;
    wire blink_counter_22;
    wire n4458;
    wire blink_counter_23;
    wire n4459;
    wire n4460;
    wire blink_counter_24;
    wire bfn_15_28_0_;
    wire n4461;
    wire blink_counter_25;
    wire data_in_19_4;
    wire \c0.FRAME_MATCHER_wait_for_transmission ;
    wire \c0.n1686 ;
    wire \c0.data_in_frame_19_4 ;
    wire CLK_c;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__37526),
            .DIN(N__37525),
            .DOUT(N__37524),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__37526),
            .PADOUT(N__37525),
            .PADIN(N__37524),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29815),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__37517),
            .DIN(N__37516),
            .DOUT(N__37515),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__37517),
            .PADOUT(N__37516),
            .PADIN(N__37515),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__37508),
            .DIN(N__37507),
            .DOUT(N__37506),
            .PACKAGEPIN(PIN_2));
    defparam rx_input_preio.PIN_TYPE=6'b000000;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__37508),
            .PADOUT(N__37507),
            .PADIN(N__37506),
            .CLOCKENABLE(VCCG0),
            .DIN0(\c0.rx.r_Rx_Data_R ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__35351),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx2_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx2_output_iopad.PULLUP=1'b1;
    IO_PAD tx2_output_iopad (
            .OE(N__37499),
            .DIN(N__37498),
            .DOUT(N__37497),
            .PACKAGEPIN(PIN_3));
    defparam tx2_output_preio.PIN_TYPE=6'b101001;
    defparam tx2_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx2_output_preio (
            .PADOEN(N__37499),
            .PADOUT(N__37498),
            .PADIN(N__37497),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12276),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__12256));
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__37490),
            .DIN(N__37489),
            .DOUT(N__37488),
            .PACKAGEPIN(PIN_1));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__37490),
            .PADOUT(N__37489),
            .PADIN(N__37488),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__16890),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__14842));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__37481),
            .DIN(N__37480),
            .DOUT(N__37479),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__37481),
            .PADOUT(N__37480),
            .PADIN(N__37479),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__9468 (
            .O(N__37462),
            .I(N__37456));
    InMux I__9467 (
            .O(N__37461),
            .I(N__37456));
    LocalMux I__9466 (
            .O(N__37456),
            .I(N__37453));
    Span4Mux_v I__9465 (
            .O(N__37453),
            .I(N__37449));
    InMux I__9464 (
            .O(N__37452),
            .I(N__37446));
    Odrv4 I__9463 (
            .O(N__37449),
            .I(blink_counter_21));
    LocalMux I__9462 (
            .O(N__37446),
            .I(blink_counter_21));
    InMux I__9461 (
            .O(N__37441),
            .I(n4457));
    InMux I__9460 (
            .O(N__37438),
            .I(N__37432));
    InMux I__9459 (
            .O(N__37437),
            .I(N__37432));
    LocalMux I__9458 (
            .O(N__37432),
            .I(N__37429));
    Span4Mux_v I__9457 (
            .O(N__37429),
            .I(N__37425));
    InMux I__9456 (
            .O(N__37428),
            .I(N__37422));
    Odrv4 I__9455 (
            .O(N__37425),
            .I(blink_counter_22));
    LocalMux I__9454 (
            .O(N__37422),
            .I(blink_counter_22));
    InMux I__9453 (
            .O(N__37417),
            .I(n4458));
    CascadeMux I__9452 (
            .O(N__37414),
            .I(N__37410));
    InMux I__9451 (
            .O(N__37413),
            .I(N__37405));
    InMux I__9450 (
            .O(N__37410),
            .I(N__37405));
    LocalMux I__9449 (
            .O(N__37405),
            .I(N__37402));
    Span4Mux_h I__9448 (
            .O(N__37402),
            .I(N__37398));
    InMux I__9447 (
            .O(N__37401),
            .I(N__37395));
    Odrv4 I__9446 (
            .O(N__37398),
            .I(blink_counter_23));
    LocalMux I__9445 (
            .O(N__37395),
            .I(blink_counter_23));
    InMux I__9444 (
            .O(N__37390),
            .I(n4459));
    CascadeMux I__9443 (
            .O(N__37387),
            .I(N__37384));
    InMux I__9442 (
            .O(N__37384),
            .I(N__37378));
    InMux I__9441 (
            .O(N__37383),
            .I(N__37378));
    LocalMux I__9440 (
            .O(N__37378),
            .I(N__37375));
    Span4Mux_v I__9439 (
            .O(N__37375),
            .I(N__37371));
    InMux I__9438 (
            .O(N__37374),
            .I(N__37368));
    Odrv4 I__9437 (
            .O(N__37371),
            .I(blink_counter_24));
    LocalMux I__9436 (
            .O(N__37368),
            .I(blink_counter_24));
    InMux I__9435 (
            .O(N__37363),
            .I(bfn_15_28_0_));
    InMux I__9434 (
            .O(N__37360),
            .I(n4461));
    InMux I__9433 (
            .O(N__37357),
            .I(N__37354));
    LocalMux I__9432 (
            .O(N__37354),
            .I(N__37351));
    Span4Mux_v I__9431 (
            .O(N__37351),
            .I(N__37347));
    InMux I__9430 (
            .O(N__37350),
            .I(N__37344));
    Odrv4 I__9429 (
            .O(N__37347),
            .I(blink_counter_25));
    LocalMux I__9428 (
            .O(N__37344),
            .I(blink_counter_25));
    InMux I__9427 (
            .O(N__37339),
            .I(N__37335));
    CascadeMux I__9426 (
            .O(N__37338),
            .I(N__37331));
    LocalMux I__9425 (
            .O(N__37335),
            .I(N__37328));
    InMux I__9424 (
            .O(N__37334),
            .I(N__37325));
    InMux I__9423 (
            .O(N__37331),
            .I(N__37322));
    Span12Mux_s7_v I__9422 (
            .O(N__37328),
            .I(N__37319));
    LocalMux I__9421 (
            .O(N__37325),
            .I(N__37316));
    LocalMux I__9420 (
            .O(N__37322),
            .I(N__37312));
    Span12Mux_h I__9419 (
            .O(N__37319),
            .I(N__37309));
    Span4Mux_h I__9418 (
            .O(N__37316),
            .I(N__37306));
    InMux I__9417 (
            .O(N__37315),
            .I(N__37303));
    Span12Mux_v I__9416 (
            .O(N__37312),
            .I(N__37300));
    Odrv12 I__9415 (
            .O(N__37309),
            .I(data_in_19_4));
    Odrv4 I__9414 (
            .O(N__37306),
            .I(data_in_19_4));
    LocalMux I__9413 (
            .O(N__37303),
            .I(data_in_19_4));
    Odrv12 I__9412 (
            .O(N__37300),
            .I(data_in_19_4));
    CascadeMux I__9411 (
            .O(N__37291),
            .I(N__37286));
    CascadeMux I__9410 (
            .O(N__37290),
            .I(N__37282));
    CascadeMux I__9409 (
            .O(N__37289),
            .I(N__37262));
    InMux I__9408 (
            .O(N__37286),
            .I(N__37258));
    InMux I__9407 (
            .O(N__37285),
            .I(N__37251));
    InMux I__9406 (
            .O(N__37282),
            .I(N__37251));
    InMux I__9405 (
            .O(N__37281),
            .I(N__37251));
    InMux I__9404 (
            .O(N__37280),
            .I(N__37243));
    InMux I__9403 (
            .O(N__37279),
            .I(N__37243));
    InMux I__9402 (
            .O(N__37278),
            .I(N__37243));
    InMux I__9401 (
            .O(N__37277),
            .I(N__37232));
    InMux I__9400 (
            .O(N__37276),
            .I(N__37232));
    InMux I__9399 (
            .O(N__37275),
            .I(N__37232));
    InMux I__9398 (
            .O(N__37274),
            .I(N__37232));
    InMux I__9397 (
            .O(N__37273),
            .I(N__37232));
    CascadeMux I__9396 (
            .O(N__37272),
            .I(N__37223));
    CascadeMux I__9395 (
            .O(N__37271),
            .I(N__37219));
    CascadeMux I__9394 (
            .O(N__37270),
            .I(N__37215));
    CascadeMux I__9393 (
            .O(N__37269),
            .I(N__37209));
    CascadeMux I__9392 (
            .O(N__37268),
            .I(N__37204));
    CascadeMux I__9391 (
            .O(N__37267),
            .I(N__37196));
    CascadeMux I__9390 (
            .O(N__37266),
            .I(N__37191));
    InMux I__9389 (
            .O(N__37265),
            .I(N__37181));
    InMux I__9388 (
            .O(N__37262),
            .I(N__37176));
    InMux I__9387 (
            .O(N__37261),
            .I(N__37176));
    LocalMux I__9386 (
            .O(N__37258),
            .I(N__37171));
    LocalMux I__9385 (
            .O(N__37251),
            .I(N__37171));
    CascadeMux I__9384 (
            .O(N__37250),
            .I(N__37168));
    LocalMux I__9383 (
            .O(N__37243),
            .I(N__37158));
    LocalMux I__9382 (
            .O(N__37232),
            .I(N__37155));
    CascadeMux I__9381 (
            .O(N__37231),
            .I(N__37139));
    CascadeMux I__9380 (
            .O(N__37230),
            .I(N__37136));
    CascadeMux I__9379 (
            .O(N__37229),
            .I(N__37133));
    CascadeMux I__9378 (
            .O(N__37228),
            .I(N__37129));
    CascadeMux I__9377 (
            .O(N__37227),
            .I(N__37120));
    CascadeMux I__9376 (
            .O(N__37226),
            .I(N__37117));
    InMux I__9375 (
            .O(N__37223),
            .I(N__37111));
    InMux I__9374 (
            .O(N__37222),
            .I(N__37111));
    InMux I__9373 (
            .O(N__37219),
            .I(N__37106));
    InMux I__9372 (
            .O(N__37218),
            .I(N__37106));
    InMux I__9371 (
            .O(N__37215),
            .I(N__37099));
    InMux I__9370 (
            .O(N__37214),
            .I(N__37099));
    InMux I__9369 (
            .O(N__37213),
            .I(N__37099));
    InMux I__9368 (
            .O(N__37212),
            .I(N__37090));
    InMux I__9367 (
            .O(N__37209),
            .I(N__37090));
    InMux I__9366 (
            .O(N__37208),
            .I(N__37090));
    InMux I__9365 (
            .O(N__37207),
            .I(N__37090));
    InMux I__9364 (
            .O(N__37204),
            .I(N__37083));
    CascadeMux I__9363 (
            .O(N__37203),
            .I(N__37080));
    InMux I__9362 (
            .O(N__37202),
            .I(N__37074));
    InMux I__9361 (
            .O(N__37201),
            .I(N__37074));
    CascadeMux I__9360 (
            .O(N__37200),
            .I(N__37071));
    InMux I__9359 (
            .O(N__37199),
            .I(N__37061));
    InMux I__9358 (
            .O(N__37196),
            .I(N__37061));
    InMux I__9357 (
            .O(N__37195),
            .I(N__37061));
    CascadeMux I__9356 (
            .O(N__37194),
            .I(N__37055));
    InMux I__9355 (
            .O(N__37191),
            .I(N__37050));
    InMux I__9354 (
            .O(N__37190),
            .I(N__37045));
    InMux I__9353 (
            .O(N__37189),
            .I(N__37045));
    InMux I__9352 (
            .O(N__37188),
            .I(N__37042));
    InMux I__9351 (
            .O(N__37187),
            .I(N__37033));
    InMux I__9350 (
            .O(N__37186),
            .I(N__37033));
    InMux I__9349 (
            .O(N__37185),
            .I(N__37033));
    InMux I__9348 (
            .O(N__37184),
            .I(N__37033));
    LocalMux I__9347 (
            .O(N__37181),
            .I(N__37026));
    LocalMux I__9346 (
            .O(N__37176),
            .I(N__37026));
    Span4Mux_h I__9345 (
            .O(N__37171),
            .I(N__37026));
    InMux I__9344 (
            .O(N__37168),
            .I(N__37021));
    InMux I__9343 (
            .O(N__37167),
            .I(N__37021));
    InMux I__9342 (
            .O(N__37166),
            .I(N__37010));
    InMux I__9341 (
            .O(N__37165),
            .I(N__37010));
    InMux I__9340 (
            .O(N__37164),
            .I(N__37010));
    InMux I__9339 (
            .O(N__37163),
            .I(N__37010));
    InMux I__9338 (
            .O(N__37162),
            .I(N__37010));
    CascadeMux I__9337 (
            .O(N__37161),
            .I(N__36993));
    Span4Mux_v I__9336 (
            .O(N__37158),
            .I(N__36984));
    Span4Mux_v I__9335 (
            .O(N__37155),
            .I(N__36984));
    InMux I__9334 (
            .O(N__37154),
            .I(N__36977));
    InMux I__9333 (
            .O(N__37153),
            .I(N__36977));
    InMux I__9332 (
            .O(N__37152),
            .I(N__36977));
    InMux I__9331 (
            .O(N__37151),
            .I(N__36966));
    InMux I__9330 (
            .O(N__37150),
            .I(N__36966));
    InMux I__9329 (
            .O(N__37149),
            .I(N__36966));
    InMux I__9328 (
            .O(N__37148),
            .I(N__36966));
    InMux I__9327 (
            .O(N__37147),
            .I(N__36966));
    InMux I__9326 (
            .O(N__37146),
            .I(N__36957));
    InMux I__9325 (
            .O(N__37145),
            .I(N__36957));
    InMux I__9324 (
            .O(N__37144),
            .I(N__36957));
    InMux I__9323 (
            .O(N__37143),
            .I(N__36957));
    InMux I__9322 (
            .O(N__37142),
            .I(N__36945));
    InMux I__9321 (
            .O(N__37139),
            .I(N__36945));
    InMux I__9320 (
            .O(N__37136),
            .I(N__36938));
    InMux I__9319 (
            .O(N__37133),
            .I(N__36938));
    InMux I__9318 (
            .O(N__37132),
            .I(N__36938));
    InMux I__9317 (
            .O(N__37129),
            .I(N__36934));
    InMux I__9316 (
            .O(N__37128),
            .I(N__36927));
    InMux I__9315 (
            .O(N__37127),
            .I(N__36927));
    InMux I__9314 (
            .O(N__37126),
            .I(N__36927));
    InMux I__9313 (
            .O(N__37125),
            .I(N__36922));
    InMux I__9312 (
            .O(N__37124),
            .I(N__36922));
    InMux I__9311 (
            .O(N__37123),
            .I(N__36913));
    InMux I__9310 (
            .O(N__37120),
            .I(N__36913));
    InMux I__9309 (
            .O(N__37117),
            .I(N__36913));
    InMux I__9308 (
            .O(N__37116),
            .I(N__36913));
    LocalMux I__9307 (
            .O(N__37111),
            .I(N__36910));
    LocalMux I__9306 (
            .O(N__37106),
            .I(N__36907));
    LocalMux I__9305 (
            .O(N__37099),
            .I(N__36902));
    LocalMux I__9304 (
            .O(N__37090),
            .I(N__36902));
    InMux I__9303 (
            .O(N__37089),
            .I(N__36895));
    InMux I__9302 (
            .O(N__37088),
            .I(N__36895));
    InMux I__9301 (
            .O(N__37087),
            .I(N__36895));
    CascadeMux I__9300 (
            .O(N__37086),
            .I(N__36890));
    LocalMux I__9299 (
            .O(N__37083),
            .I(N__36885));
    InMux I__9298 (
            .O(N__37080),
            .I(N__36882));
    CascadeMux I__9297 (
            .O(N__37079),
            .I(N__36877));
    LocalMux I__9296 (
            .O(N__37074),
            .I(N__36874));
    InMux I__9295 (
            .O(N__37071),
            .I(N__36865));
    InMux I__9294 (
            .O(N__37070),
            .I(N__36865));
    InMux I__9293 (
            .O(N__37069),
            .I(N__36865));
    InMux I__9292 (
            .O(N__37068),
            .I(N__36865));
    LocalMux I__9291 (
            .O(N__37061),
            .I(N__36862));
    InMux I__9290 (
            .O(N__37060),
            .I(N__36857));
    InMux I__9289 (
            .O(N__37059),
            .I(N__36857));
    InMux I__9288 (
            .O(N__37058),
            .I(N__36854));
    InMux I__9287 (
            .O(N__37055),
            .I(N__36849));
    InMux I__9286 (
            .O(N__37054),
            .I(N__36849));
    InMux I__9285 (
            .O(N__37053),
            .I(N__36842));
    LocalMux I__9284 (
            .O(N__37050),
            .I(N__36837));
    LocalMux I__9283 (
            .O(N__37045),
            .I(N__36837));
    LocalMux I__9282 (
            .O(N__37042),
            .I(N__36826));
    LocalMux I__9281 (
            .O(N__37033),
            .I(N__36826));
    Span4Mux_h I__9280 (
            .O(N__37026),
            .I(N__36826));
    LocalMux I__9279 (
            .O(N__37021),
            .I(N__36826));
    LocalMux I__9278 (
            .O(N__37010),
            .I(N__36826));
    InMux I__9277 (
            .O(N__37009),
            .I(N__36823));
    InMux I__9276 (
            .O(N__37008),
            .I(N__36816));
    InMux I__9275 (
            .O(N__37007),
            .I(N__36816));
    InMux I__9274 (
            .O(N__37006),
            .I(N__36816));
    CascadeMux I__9273 (
            .O(N__37005),
            .I(N__36811));
    CascadeMux I__9272 (
            .O(N__37004),
            .I(N__36808));
    CascadeMux I__9271 (
            .O(N__37003),
            .I(N__36799));
    CascadeMux I__9270 (
            .O(N__37002),
            .I(N__36795));
    CascadeMux I__9269 (
            .O(N__37001),
            .I(N__36792));
    CascadeMux I__9268 (
            .O(N__37000),
            .I(N__36788));
    CascadeMux I__9267 (
            .O(N__36999),
            .I(N__36782));
    InMux I__9266 (
            .O(N__36998),
            .I(N__36775));
    InMux I__9265 (
            .O(N__36997),
            .I(N__36775));
    InMux I__9264 (
            .O(N__36996),
            .I(N__36775));
    InMux I__9263 (
            .O(N__36993),
            .I(N__36766));
    InMux I__9262 (
            .O(N__36992),
            .I(N__36766));
    InMux I__9261 (
            .O(N__36991),
            .I(N__36766));
    InMux I__9260 (
            .O(N__36990),
            .I(N__36766));
    InMux I__9259 (
            .O(N__36989),
            .I(N__36763));
    Span4Mux_v I__9258 (
            .O(N__36984),
            .I(N__36760));
    LocalMux I__9257 (
            .O(N__36977),
            .I(N__36757));
    LocalMux I__9256 (
            .O(N__36966),
            .I(N__36752));
    LocalMux I__9255 (
            .O(N__36957),
            .I(N__36752));
    InMux I__9254 (
            .O(N__36956),
            .I(N__36745));
    InMux I__9253 (
            .O(N__36955),
            .I(N__36745));
    InMux I__9252 (
            .O(N__36954),
            .I(N__36745));
    InMux I__9251 (
            .O(N__36953),
            .I(N__36742));
    InMux I__9250 (
            .O(N__36952),
            .I(N__36739));
    InMux I__9249 (
            .O(N__36951),
            .I(N__36734));
    InMux I__9248 (
            .O(N__36950),
            .I(N__36734));
    LocalMux I__9247 (
            .O(N__36945),
            .I(N__36729));
    LocalMux I__9246 (
            .O(N__36938),
            .I(N__36729));
    InMux I__9245 (
            .O(N__36937),
            .I(N__36726));
    LocalMux I__9244 (
            .O(N__36934),
            .I(N__36723));
    LocalMux I__9243 (
            .O(N__36927),
            .I(N__36716));
    LocalMux I__9242 (
            .O(N__36922),
            .I(N__36716));
    LocalMux I__9241 (
            .O(N__36913),
            .I(N__36716));
    Span4Mux_v I__9240 (
            .O(N__36910),
            .I(N__36711));
    Span4Mux_h I__9239 (
            .O(N__36907),
            .I(N__36711));
    Span4Mux_h I__9238 (
            .O(N__36902),
            .I(N__36706));
    LocalMux I__9237 (
            .O(N__36895),
            .I(N__36706));
    InMux I__9236 (
            .O(N__36894),
            .I(N__36699));
    InMux I__9235 (
            .O(N__36893),
            .I(N__36699));
    InMux I__9234 (
            .O(N__36890),
            .I(N__36692));
    InMux I__9233 (
            .O(N__36889),
            .I(N__36692));
    InMux I__9232 (
            .O(N__36888),
            .I(N__36692));
    Span4Mux_s3_h I__9231 (
            .O(N__36885),
            .I(N__36686));
    LocalMux I__9230 (
            .O(N__36882),
            .I(N__36686));
    InMux I__9229 (
            .O(N__36881),
            .I(N__36681));
    InMux I__9228 (
            .O(N__36880),
            .I(N__36681));
    InMux I__9227 (
            .O(N__36877),
            .I(N__36678));
    Span4Mux_h I__9226 (
            .O(N__36874),
            .I(N__36673));
    LocalMux I__9225 (
            .O(N__36865),
            .I(N__36673));
    Span4Mux_h I__9224 (
            .O(N__36862),
            .I(N__36666));
    LocalMux I__9223 (
            .O(N__36857),
            .I(N__36666));
    LocalMux I__9222 (
            .O(N__36854),
            .I(N__36666));
    LocalMux I__9221 (
            .O(N__36849),
            .I(N__36663));
    InMux I__9220 (
            .O(N__36848),
            .I(N__36654));
    InMux I__9219 (
            .O(N__36847),
            .I(N__36654));
    InMux I__9218 (
            .O(N__36846),
            .I(N__36654));
    InMux I__9217 (
            .O(N__36845),
            .I(N__36654));
    LocalMux I__9216 (
            .O(N__36842),
            .I(N__36651));
    Span4Mux_h I__9215 (
            .O(N__36837),
            .I(N__36640));
    Span4Mux_v I__9214 (
            .O(N__36826),
            .I(N__36640));
    LocalMux I__9213 (
            .O(N__36823),
            .I(N__36640));
    LocalMux I__9212 (
            .O(N__36816),
            .I(N__36640));
    InMux I__9211 (
            .O(N__36815),
            .I(N__36630));
    InMux I__9210 (
            .O(N__36814),
            .I(N__36630));
    InMux I__9209 (
            .O(N__36811),
            .I(N__36627));
    InMux I__9208 (
            .O(N__36808),
            .I(N__36622));
    InMux I__9207 (
            .O(N__36807),
            .I(N__36622));
    InMux I__9206 (
            .O(N__36806),
            .I(N__36615));
    InMux I__9205 (
            .O(N__36805),
            .I(N__36615));
    InMux I__9204 (
            .O(N__36804),
            .I(N__36615));
    InMux I__9203 (
            .O(N__36803),
            .I(N__36612));
    InMux I__9202 (
            .O(N__36802),
            .I(N__36609));
    InMux I__9201 (
            .O(N__36799),
            .I(N__36599));
    InMux I__9200 (
            .O(N__36798),
            .I(N__36599));
    InMux I__9199 (
            .O(N__36795),
            .I(N__36592));
    InMux I__9198 (
            .O(N__36792),
            .I(N__36592));
    InMux I__9197 (
            .O(N__36791),
            .I(N__36592));
    InMux I__9196 (
            .O(N__36788),
            .I(N__36587));
    InMux I__9195 (
            .O(N__36787),
            .I(N__36587));
    InMux I__9194 (
            .O(N__36786),
            .I(N__36584));
    InMux I__9193 (
            .O(N__36785),
            .I(N__36579));
    InMux I__9192 (
            .O(N__36782),
            .I(N__36579));
    LocalMux I__9191 (
            .O(N__36775),
            .I(N__36574));
    LocalMux I__9190 (
            .O(N__36766),
            .I(N__36574));
    LocalMux I__9189 (
            .O(N__36763),
            .I(N__36567));
    Span4Mux_h I__9188 (
            .O(N__36760),
            .I(N__36567));
    Span4Mux_v I__9187 (
            .O(N__36757),
            .I(N__36567));
    Span4Mux_s3_v I__9186 (
            .O(N__36752),
            .I(N__36562));
    LocalMux I__9185 (
            .O(N__36745),
            .I(N__36562));
    LocalMux I__9184 (
            .O(N__36742),
            .I(N__36557));
    LocalMux I__9183 (
            .O(N__36739),
            .I(N__36557));
    LocalMux I__9182 (
            .O(N__36734),
            .I(N__36542));
    Span4Mux_s3_v I__9181 (
            .O(N__36729),
            .I(N__36542));
    LocalMux I__9180 (
            .O(N__36726),
            .I(N__36542));
    Span4Mux_h I__9179 (
            .O(N__36723),
            .I(N__36542));
    Span4Mux_h I__9178 (
            .O(N__36716),
            .I(N__36542));
    Span4Mux_h I__9177 (
            .O(N__36711),
            .I(N__36542));
    Span4Mux_h I__9176 (
            .O(N__36706),
            .I(N__36542));
    InMux I__9175 (
            .O(N__36705),
            .I(N__36537));
    InMux I__9174 (
            .O(N__36704),
            .I(N__36537));
    LocalMux I__9173 (
            .O(N__36699),
            .I(N__36532));
    LocalMux I__9172 (
            .O(N__36692),
            .I(N__36532));
    InMux I__9171 (
            .O(N__36691),
            .I(N__36529));
    Span4Mux_v I__9170 (
            .O(N__36686),
            .I(N__36524));
    LocalMux I__9169 (
            .O(N__36681),
            .I(N__36524));
    LocalMux I__9168 (
            .O(N__36678),
            .I(N__36513));
    Span4Mux_v I__9167 (
            .O(N__36673),
            .I(N__36513));
    Span4Mux_v I__9166 (
            .O(N__36666),
            .I(N__36513));
    Span4Mux_v I__9165 (
            .O(N__36663),
            .I(N__36513));
    LocalMux I__9164 (
            .O(N__36654),
            .I(N__36513));
    Span4Mux_h I__9163 (
            .O(N__36651),
            .I(N__36510));
    CascadeMux I__9162 (
            .O(N__36650),
            .I(N__36505));
    CascadeMux I__9161 (
            .O(N__36649),
            .I(N__36502));
    Span4Mux_v I__9160 (
            .O(N__36640),
            .I(N__36497));
    InMux I__9159 (
            .O(N__36639),
            .I(N__36491));
    InMux I__9158 (
            .O(N__36638),
            .I(N__36486));
    InMux I__9157 (
            .O(N__36637),
            .I(N__36486));
    CascadeMux I__9156 (
            .O(N__36636),
            .I(N__36483));
    CascadeMux I__9155 (
            .O(N__36635),
            .I(N__36479));
    LocalMux I__9154 (
            .O(N__36630),
            .I(N__36466));
    LocalMux I__9153 (
            .O(N__36627),
            .I(N__36466));
    LocalMux I__9152 (
            .O(N__36622),
            .I(N__36466));
    LocalMux I__9151 (
            .O(N__36615),
            .I(N__36466));
    LocalMux I__9150 (
            .O(N__36612),
            .I(N__36466));
    LocalMux I__9149 (
            .O(N__36609),
            .I(N__36466));
    InMux I__9148 (
            .O(N__36608),
            .I(N__36455));
    InMux I__9147 (
            .O(N__36607),
            .I(N__36455));
    InMux I__9146 (
            .O(N__36606),
            .I(N__36455));
    InMux I__9145 (
            .O(N__36605),
            .I(N__36455));
    InMux I__9144 (
            .O(N__36604),
            .I(N__36455));
    LocalMux I__9143 (
            .O(N__36599),
            .I(N__36446));
    LocalMux I__9142 (
            .O(N__36592),
            .I(N__36446));
    LocalMux I__9141 (
            .O(N__36587),
            .I(N__36446));
    LocalMux I__9140 (
            .O(N__36584),
            .I(N__36446));
    LocalMux I__9139 (
            .O(N__36579),
            .I(N__36441));
    Span4Mux_v I__9138 (
            .O(N__36574),
            .I(N__36441));
    Span4Mux_h I__9137 (
            .O(N__36567),
            .I(N__36438));
    Span4Mux_v I__9136 (
            .O(N__36562),
            .I(N__36430));
    Span4Mux_h I__9135 (
            .O(N__36557),
            .I(N__36430));
    Span4Mux_v I__9134 (
            .O(N__36542),
            .I(N__36430));
    LocalMux I__9133 (
            .O(N__36537),
            .I(N__36425));
    Span4Mux_v I__9132 (
            .O(N__36532),
            .I(N__36425));
    LocalMux I__9131 (
            .O(N__36529),
            .I(N__36416));
    Span4Mux_h I__9130 (
            .O(N__36524),
            .I(N__36416));
    Span4Mux_h I__9129 (
            .O(N__36513),
            .I(N__36416));
    Span4Mux_v I__9128 (
            .O(N__36510),
            .I(N__36416));
    InMux I__9127 (
            .O(N__36509),
            .I(N__36413));
    InMux I__9126 (
            .O(N__36508),
            .I(N__36402));
    InMux I__9125 (
            .O(N__36505),
            .I(N__36402));
    InMux I__9124 (
            .O(N__36502),
            .I(N__36402));
    InMux I__9123 (
            .O(N__36501),
            .I(N__36402));
    InMux I__9122 (
            .O(N__36500),
            .I(N__36402));
    Span4Mux_h I__9121 (
            .O(N__36497),
            .I(N__36399));
    InMux I__9120 (
            .O(N__36496),
            .I(N__36392));
    InMux I__9119 (
            .O(N__36495),
            .I(N__36392));
    InMux I__9118 (
            .O(N__36494),
            .I(N__36392));
    LocalMux I__9117 (
            .O(N__36491),
            .I(N__36387));
    LocalMux I__9116 (
            .O(N__36486),
            .I(N__36387));
    InMux I__9115 (
            .O(N__36483),
            .I(N__36380));
    InMux I__9114 (
            .O(N__36482),
            .I(N__36380));
    InMux I__9113 (
            .O(N__36479),
            .I(N__36380));
    Span12Mux_h I__9112 (
            .O(N__36466),
            .I(N__36377));
    LocalMux I__9111 (
            .O(N__36455),
            .I(N__36368));
    Span4Mux_v I__9110 (
            .O(N__36446),
            .I(N__36368));
    Span4Mux_v I__9109 (
            .O(N__36441),
            .I(N__36368));
    Span4Mux_v I__9108 (
            .O(N__36438),
            .I(N__36368));
    InMux I__9107 (
            .O(N__36437),
            .I(N__36365));
    Span4Mux_h I__9106 (
            .O(N__36430),
            .I(N__36362));
    Span4Mux_h I__9105 (
            .O(N__36425),
            .I(N__36357));
    Span4Mux_v I__9104 (
            .O(N__36416),
            .I(N__36357));
    LocalMux I__9103 (
            .O(N__36413),
            .I(N__36350));
    LocalMux I__9102 (
            .O(N__36402),
            .I(N__36350));
    Span4Mux_h I__9101 (
            .O(N__36399),
            .I(N__36350));
    LocalMux I__9100 (
            .O(N__36392),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv12 I__9099 (
            .O(N__36387),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    LocalMux I__9098 (
            .O(N__36380),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv12 I__9097 (
            .O(N__36377),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__9096 (
            .O(N__36368),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    LocalMux I__9095 (
            .O(N__36365),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__9094 (
            .O(N__36362),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__9093 (
            .O(N__36357),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__9092 (
            .O(N__36350),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    CascadeMux I__9091 (
            .O(N__36331),
            .I(N__36324));
    CascadeMux I__9090 (
            .O(N__36330),
            .I(N__36316));
    InMux I__9089 (
            .O(N__36329),
            .I(N__36302));
    InMux I__9088 (
            .O(N__36328),
            .I(N__36302));
    InMux I__9087 (
            .O(N__36327),
            .I(N__36302));
    InMux I__9086 (
            .O(N__36324),
            .I(N__36299));
    InMux I__9085 (
            .O(N__36323),
            .I(N__36294));
    InMux I__9084 (
            .O(N__36322),
            .I(N__36294));
    InMux I__9083 (
            .O(N__36321),
            .I(N__36282));
    InMux I__9082 (
            .O(N__36320),
            .I(N__36282));
    InMux I__9081 (
            .O(N__36319),
            .I(N__36282));
    InMux I__9080 (
            .O(N__36316),
            .I(N__36277));
    InMux I__9079 (
            .O(N__36315),
            .I(N__36277));
    InMux I__9078 (
            .O(N__36314),
            .I(N__36274));
    CascadeMux I__9077 (
            .O(N__36313),
            .I(N__36267));
    InMux I__9076 (
            .O(N__36312),
            .I(N__36258));
    InMux I__9075 (
            .O(N__36311),
            .I(N__36244));
    InMux I__9074 (
            .O(N__36310),
            .I(N__36244));
    InMux I__9073 (
            .O(N__36309),
            .I(N__36244));
    LocalMux I__9072 (
            .O(N__36302),
            .I(N__36241));
    LocalMux I__9071 (
            .O(N__36299),
            .I(N__36236));
    LocalMux I__9070 (
            .O(N__36294),
            .I(N__36236));
    CascadeMux I__9069 (
            .O(N__36293),
            .I(N__36232));
    InMux I__9068 (
            .O(N__36292),
            .I(N__36219));
    CascadeMux I__9067 (
            .O(N__36291),
            .I(N__36212));
    CascadeMux I__9066 (
            .O(N__36290),
            .I(N__36209));
    InMux I__9065 (
            .O(N__36289),
            .I(N__36190));
    LocalMux I__9064 (
            .O(N__36282),
            .I(N__36183));
    LocalMux I__9063 (
            .O(N__36277),
            .I(N__36183));
    LocalMux I__9062 (
            .O(N__36274),
            .I(N__36183));
    InMux I__9061 (
            .O(N__36273),
            .I(N__36176));
    InMux I__9060 (
            .O(N__36272),
            .I(N__36176));
    InMux I__9059 (
            .O(N__36271),
            .I(N__36176));
    CascadeMux I__9058 (
            .O(N__36270),
            .I(N__36164));
    InMux I__9057 (
            .O(N__36267),
            .I(N__36154));
    InMux I__9056 (
            .O(N__36266),
            .I(N__36154));
    InMux I__9055 (
            .O(N__36265),
            .I(N__36147));
    InMux I__9054 (
            .O(N__36264),
            .I(N__36147));
    InMux I__9053 (
            .O(N__36263),
            .I(N__36147));
    CascadeMux I__9052 (
            .O(N__36262),
            .I(N__36143));
    CascadeMux I__9051 (
            .O(N__36261),
            .I(N__36140));
    LocalMux I__9050 (
            .O(N__36258),
            .I(N__36137));
    InMux I__9049 (
            .O(N__36257),
            .I(N__36130));
    InMux I__9048 (
            .O(N__36256),
            .I(N__36130));
    InMux I__9047 (
            .O(N__36255),
            .I(N__36130));
    InMux I__9046 (
            .O(N__36254),
            .I(N__36123));
    InMux I__9045 (
            .O(N__36253),
            .I(N__36123));
    InMux I__9044 (
            .O(N__36252),
            .I(N__36123));
    InMux I__9043 (
            .O(N__36251),
            .I(N__36120));
    LocalMux I__9042 (
            .O(N__36244),
            .I(N__36113));
    Span4Mux_v I__9041 (
            .O(N__36241),
            .I(N__36113));
    Span4Mux_v I__9040 (
            .O(N__36236),
            .I(N__36113));
    InMux I__9039 (
            .O(N__36235),
            .I(N__36102));
    InMux I__9038 (
            .O(N__36232),
            .I(N__36102));
    InMux I__9037 (
            .O(N__36231),
            .I(N__36102));
    InMux I__9036 (
            .O(N__36230),
            .I(N__36102));
    InMux I__9035 (
            .O(N__36229),
            .I(N__36102));
    InMux I__9034 (
            .O(N__36228),
            .I(N__36096));
    InMux I__9033 (
            .O(N__36227),
            .I(N__36096));
    InMux I__9032 (
            .O(N__36226),
            .I(N__36091));
    InMux I__9031 (
            .O(N__36225),
            .I(N__36091));
    CascadeMux I__9030 (
            .O(N__36224),
            .I(N__36088));
    InMux I__9029 (
            .O(N__36223),
            .I(N__36076));
    InMux I__9028 (
            .O(N__36222),
            .I(N__36076));
    LocalMux I__9027 (
            .O(N__36219),
            .I(N__36073));
    InMux I__9026 (
            .O(N__36218),
            .I(N__36064));
    InMux I__9025 (
            .O(N__36217),
            .I(N__36064));
    InMux I__9024 (
            .O(N__36216),
            .I(N__36064));
    InMux I__9023 (
            .O(N__36215),
            .I(N__36064));
    InMux I__9022 (
            .O(N__36212),
            .I(N__36050));
    InMux I__9021 (
            .O(N__36209),
            .I(N__36050));
    InMux I__9020 (
            .O(N__36208),
            .I(N__36050));
    InMux I__9019 (
            .O(N__36207),
            .I(N__36045));
    InMux I__9018 (
            .O(N__36206),
            .I(N__36045));
    InMux I__9017 (
            .O(N__36205),
            .I(N__36042));
    CascadeMux I__9016 (
            .O(N__36204),
            .I(N__36027));
    InMux I__9015 (
            .O(N__36203),
            .I(N__36019));
    InMux I__9014 (
            .O(N__36202),
            .I(N__36019));
    InMux I__9013 (
            .O(N__36201),
            .I(N__36014));
    CascadeMux I__9012 (
            .O(N__36200),
            .I(N__36007));
    InMux I__9011 (
            .O(N__36199),
            .I(N__36000));
    InMux I__9010 (
            .O(N__36198),
            .I(N__36000));
    InMux I__9009 (
            .O(N__36197),
            .I(N__35997));
    CascadeMux I__9008 (
            .O(N__36196),
            .I(N__35993));
    InMux I__9007 (
            .O(N__36195),
            .I(N__35981));
    InMux I__9006 (
            .O(N__36194),
            .I(N__35981));
    CascadeMux I__9005 (
            .O(N__36193),
            .I(N__35978));
    LocalMux I__9004 (
            .O(N__36190),
            .I(N__35975));
    Span4Mux_v I__9003 (
            .O(N__36183),
            .I(N__35970));
    LocalMux I__9002 (
            .O(N__36176),
            .I(N__35970));
    InMux I__9001 (
            .O(N__36175),
            .I(N__35967));
    InMux I__9000 (
            .O(N__36174),
            .I(N__35961));
    InMux I__8999 (
            .O(N__36173),
            .I(N__35956));
    InMux I__8998 (
            .O(N__36172),
            .I(N__35956));
    InMux I__8997 (
            .O(N__36171),
            .I(N__35951));
    InMux I__8996 (
            .O(N__36170),
            .I(N__35951));
    InMux I__8995 (
            .O(N__36169),
            .I(N__35944));
    InMux I__8994 (
            .O(N__36168),
            .I(N__35944));
    InMux I__8993 (
            .O(N__36167),
            .I(N__35944));
    InMux I__8992 (
            .O(N__36164),
            .I(N__35939));
    InMux I__8991 (
            .O(N__36163),
            .I(N__35939));
    InMux I__8990 (
            .O(N__36162),
            .I(N__35930));
    InMux I__8989 (
            .O(N__36161),
            .I(N__35930));
    InMux I__8988 (
            .O(N__36160),
            .I(N__35930));
    InMux I__8987 (
            .O(N__36159),
            .I(N__35930));
    LocalMux I__8986 (
            .O(N__36154),
            .I(N__35925));
    LocalMux I__8985 (
            .O(N__36147),
            .I(N__35925));
    InMux I__8984 (
            .O(N__36146),
            .I(N__35922));
    InMux I__8983 (
            .O(N__36143),
            .I(N__35917));
    InMux I__8982 (
            .O(N__36140),
            .I(N__35917));
    Span4Mux_s1_v I__8981 (
            .O(N__36137),
            .I(N__35904));
    LocalMux I__8980 (
            .O(N__36130),
            .I(N__35904));
    LocalMux I__8979 (
            .O(N__36123),
            .I(N__35904));
    LocalMux I__8978 (
            .O(N__36120),
            .I(N__35904));
    Span4Mux_h I__8977 (
            .O(N__36113),
            .I(N__35904));
    LocalMux I__8976 (
            .O(N__36102),
            .I(N__35904));
    InMux I__8975 (
            .O(N__36101),
            .I(N__35901));
    LocalMux I__8974 (
            .O(N__36096),
            .I(N__35896));
    LocalMux I__8973 (
            .O(N__36091),
            .I(N__35896));
    InMux I__8972 (
            .O(N__36088),
            .I(N__35887));
    InMux I__8971 (
            .O(N__36087),
            .I(N__35887));
    InMux I__8970 (
            .O(N__36086),
            .I(N__35887));
    InMux I__8969 (
            .O(N__36085),
            .I(N__35887));
    InMux I__8968 (
            .O(N__36084),
            .I(N__35878));
    InMux I__8967 (
            .O(N__36083),
            .I(N__35878));
    InMux I__8966 (
            .O(N__36082),
            .I(N__35878));
    InMux I__8965 (
            .O(N__36081),
            .I(N__35878));
    LocalMux I__8964 (
            .O(N__36076),
            .I(N__35875));
    Span4Mux_h I__8963 (
            .O(N__36073),
            .I(N__35870));
    LocalMux I__8962 (
            .O(N__36064),
            .I(N__35870));
    InMux I__8961 (
            .O(N__36063),
            .I(N__35865));
    InMux I__8960 (
            .O(N__36062),
            .I(N__35865));
    InMux I__8959 (
            .O(N__36061),
            .I(N__35846));
    InMux I__8958 (
            .O(N__36060),
            .I(N__35846));
    InMux I__8957 (
            .O(N__36059),
            .I(N__35846));
    InMux I__8956 (
            .O(N__36058),
            .I(N__35846));
    InMux I__8955 (
            .O(N__36057),
            .I(N__35846));
    LocalMux I__8954 (
            .O(N__36050),
            .I(N__35839));
    LocalMux I__8953 (
            .O(N__36045),
            .I(N__35839));
    LocalMux I__8952 (
            .O(N__36042),
            .I(N__35839));
    InMux I__8951 (
            .O(N__36041),
            .I(N__35832));
    InMux I__8950 (
            .O(N__36040),
            .I(N__35832));
    InMux I__8949 (
            .O(N__36039),
            .I(N__35825));
    InMux I__8948 (
            .O(N__36038),
            .I(N__35825));
    InMux I__8947 (
            .O(N__36037),
            .I(N__35825));
    InMux I__8946 (
            .O(N__36036),
            .I(N__35818));
    InMux I__8945 (
            .O(N__36035),
            .I(N__35818));
    InMux I__8944 (
            .O(N__36034),
            .I(N__35818));
    InMux I__8943 (
            .O(N__36033),
            .I(N__35809));
    InMux I__8942 (
            .O(N__36032),
            .I(N__35809));
    InMux I__8941 (
            .O(N__36031),
            .I(N__35809));
    InMux I__8940 (
            .O(N__36030),
            .I(N__35809));
    InMux I__8939 (
            .O(N__36027),
            .I(N__35800));
    InMux I__8938 (
            .O(N__36026),
            .I(N__35800));
    InMux I__8937 (
            .O(N__36025),
            .I(N__35800));
    InMux I__8936 (
            .O(N__36024),
            .I(N__35800));
    LocalMux I__8935 (
            .O(N__36019),
            .I(N__35797));
    InMux I__8934 (
            .O(N__36018),
            .I(N__35792));
    InMux I__8933 (
            .O(N__36017),
            .I(N__35792));
    LocalMux I__8932 (
            .O(N__36014),
            .I(N__35789));
    InMux I__8931 (
            .O(N__36013),
            .I(N__35786));
    InMux I__8930 (
            .O(N__36012),
            .I(N__35781));
    InMux I__8929 (
            .O(N__36011),
            .I(N__35781));
    InMux I__8928 (
            .O(N__36010),
            .I(N__35772));
    InMux I__8927 (
            .O(N__36007),
            .I(N__35772));
    InMux I__8926 (
            .O(N__36006),
            .I(N__35772));
    InMux I__8925 (
            .O(N__36005),
            .I(N__35772));
    LocalMux I__8924 (
            .O(N__36000),
            .I(N__35769));
    LocalMux I__8923 (
            .O(N__35997),
            .I(N__35765));
    InMux I__8922 (
            .O(N__35996),
            .I(N__35762));
    InMux I__8921 (
            .O(N__35993),
            .I(N__35755));
    InMux I__8920 (
            .O(N__35992),
            .I(N__35755));
    InMux I__8919 (
            .O(N__35991),
            .I(N__35755));
    InMux I__8918 (
            .O(N__35990),
            .I(N__35744));
    InMux I__8917 (
            .O(N__35989),
            .I(N__35744));
    InMux I__8916 (
            .O(N__35988),
            .I(N__35744));
    InMux I__8915 (
            .O(N__35987),
            .I(N__35744));
    InMux I__8914 (
            .O(N__35986),
            .I(N__35744));
    LocalMux I__8913 (
            .O(N__35981),
            .I(N__35741));
    InMux I__8912 (
            .O(N__35978),
            .I(N__35738));
    Span4Mux_v I__8911 (
            .O(N__35975),
            .I(N__35735));
    Span4Mux_h I__8910 (
            .O(N__35970),
            .I(N__35730));
    LocalMux I__8909 (
            .O(N__35967),
            .I(N__35730));
    InMux I__8908 (
            .O(N__35966),
            .I(N__35727));
    InMux I__8907 (
            .O(N__35965),
            .I(N__35722));
    InMux I__8906 (
            .O(N__35964),
            .I(N__35722));
    LocalMux I__8905 (
            .O(N__35961),
            .I(N__35717));
    LocalMux I__8904 (
            .O(N__35956),
            .I(N__35717));
    LocalMux I__8903 (
            .O(N__35951),
            .I(N__35706));
    LocalMux I__8902 (
            .O(N__35944),
            .I(N__35706));
    LocalMux I__8901 (
            .O(N__35939),
            .I(N__35706));
    LocalMux I__8900 (
            .O(N__35930),
            .I(N__35706));
    Span4Mux_v I__8899 (
            .O(N__35925),
            .I(N__35706));
    LocalMux I__8898 (
            .O(N__35922),
            .I(N__35701));
    LocalMux I__8897 (
            .O(N__35917),
            .I(N__35701));
    Span4Mux_v I__8896 (
            .O(N__35904),
            .I(N__35698));
    LocalMux I__8895 (
            .O(N__35901),
            .I(N__35683));
    Span4Mux_h I__8894 (
            .O(N__35896),
            .I(N__35683));
    LocalMux I__8893 (
            .O(N__35887),
            .I(N__35683));
    LocalMux I__8892 (
            .O(N__35878),
            .I(N__35683));
    Span4Mux_v I__8891 (
            .O(N__35875),
            .I(N__35683));
    Span4Mux_h I__8890 (
            .O(N__35870),
            .I(N__35683));
    LocalMux I__8889 (
            .O(N__35865),
            .I(N__35683));
    InMux I__8888 (
            .O(N__35864),
            .I(N__35680));
    InMux I__8887 (
            .O(N__35863),
            .I(N__35677));
    InMux I__8886 (
            .O(N__35862),
            .I(N__35674));
    InMux I__8885 (
            .O(N__35861),
            .I(N__35663));
    InMux I__8884 (
            .O(N__35860),
            .I(N__35663));
    InMux I__8883 (
            .O(N__35859),
            .I(N__35663));
    InMux I__8882 (
            .O(N__35858),
            .I(N__35663));
    InMux I__8881 (
            .O(N__35857),
            .I(N__35663));
    LocalMux I__8880 (
            .O(N__35846),
            .I(N__35660));
    Span4Mux_v I__8879 (
            .O(N__35839),
            .I(N__35657));
    InMux I__8878 (
            .O(N__35838),
            .I(N__35654));
    CascadeMux I__8877 (
            .O(N__35837),
            .I(N__35636));
    LocalMux I__8876 (
            .O(N__35832),
            .I(N__35633));
    LocalMux I__8875 (
            .O(N__35825),
            .I(N__35628));
    LocalMux I__8874 (
            .O(N__35818),
            .I(N__35628));
    LocalMux I__8873 (
            .O(N__35809),
            .I(N__35625));
    LocalMux I__8872 (
            .O(N__35800),
            .I(N__35620));
    Span4Mux_v I__8871 (
            .O(N__35797),
            .I(N__35620));
    LocalMux I__8870 (
            .O(N__35792),
            .I(N__35615));
    Span4Mux_v I__8869 (
            .O(N__35789),
            .I(N__35615));
    LocalMux I__8868 (
            .O(N__35786),
            .I(N__35606));
    LocalMux I__8867 (
            .O(N__35781),
            .I(N__35606));
    LocalMux I__8866 (
            .O(N__35772),
            .I(N__35606));
    Span4Mux_v I__8865 (
            .O(N__35769),
            .I(N__35606));
    InMux I__8864 (
            .O(N__35768),
            .I(N__35603));
    Span4Mux_v I__8863 (
            .O(N__35765),
            .I(N__35600));
    LocalMux I__8862 (
            .O(N__35762),
            .I(N__35595));
    LocalMux I__8861 (
            .O(N__35755),
            .I(N__35595));
    LocalMux I__8860 (
            .O(N__35744),
            .I(N__35590));
    Span4Mux_v I__8859 (
            .O(N__35741),
            .I(N__35590));
    LocalMux I__8858 (
            .O(N__35738),
            .I(N__35583));
    Span4Mux_s0_h I__8857 (
            .O(N__35735),
            .I(N__35583));
    Span4Mux_v I__8856 (
            .O(N__35730),
            .I(N__35583));
    LocalMux I__8855 (
            .O(N__35727),
            .I(N__35574));
    LocalMux I__8854 (
            .O(N__35722),
            .I(N__35574));
    Span4Mux_v I__8853 (
            .O(N__35717),
            .I(N__35574));
    Span4Mux_v I__8852 (
            .O(N__35706),
            .I(N__35574));
    Span4Mux_v I__8851 (
            .O(N__35701),
            .I(N__35571));
    Span4Mux_s1_v I__8850 (
            .O(N__35698),
            .I(N__35566));
    Span4Mux_v I__8849 (
            .O(N__35683),
            .I(N__35566));
    LocalMux I__8848 (
            .O(N__35680),
            .I(N__35559));
    LocalMux I__8847 (
            .O(N__35677),
            .I(N__35559));
    LocalMux I__8846 (
            .O(N__35674),
            .I(N__35559));
    LocalMux I__8845 (
            .O(N__35663),
            .I(N__35556));
    Span4Mux_h I__8844 (
            .O(N__35660),
            .I(N__35549));
    Span4Mux_h I__8843 (
            .O(N__35657),
            .I(N__35549));
    LocalMux I__8842 (
            .O(N__35654),
            .I(N__35549));
    InMux I__8841 (
            .O(N__35653),
            .I(N__35546));
    InMux I__8840 (
            .O(N__35652),
            .I(N__35543));
    InMux I__8839 (
            .O(N__35651),
            .I(N__35536));
    InMux I__8838 (
            .O(N__35650),
            .I(N__35536));
    InMux I__8837 (
            .O(N__35649),
            .I(N__35536));
    InMux I__8836 (
            .O(N__35648),
            .I(N__35529));
    InMux I__8835 (
            .O(N__35647),
            .I(N__35529));
    InMux I__8834 (
            .O(N__35646),
            .I(N__35529));
    InMux I__8833 (
            .O(N__35645),
            .I(N__35524));
    InMux I__8832 (
            .O(N__35644),
            .I(N__35524));
    InMux I__8831 (
            .O(N__35643),
            .I(N__35517));
    InMux I__8830 (
            .O(N__35642),
            .I(N__35517));
    InMux I__8829 (
            .O(N__35641),
            .I(N__35517));
    InMux I__8828 (
            .O(N__35640),
            .I(N__35512));
    InMux I__8827 (
            .O(N__35639),
            .I(N__35512));
    InMux I__8826 (
            .O(N__35636),
            .I(N__35509));
    Span4Mux_h I__8825 (
            .O(N__35633),
            .I(N__35506));
    Span4Mux_h I__8824 (
            .O(N__35628),
            .I(N__35503));
    Span4Mux_v I__8823 (
            .O(N__35625),
            .I(N__35494));
    Span4Mux_h I__8822 (
            .O(N__35620),
            .I(N__35494));
    Span4Mux_v I__8821 (
            .O(N__35615),
            .I(N__35494));
    Span4Mux_v I__8820 (
            .O(N__35606),
            .I(N__35494));
    LocalMux I__8819 (
            .O(N__35603),
            .I(N__35481));
    Span4Mux_s1_v I__8818 (
            .O(N__35600),
            .I(N__35481));
    Span4Mux_v I__8817 (
            .O(N__35595),
            .I(N__35481));
    Span4Mux_v I__8816 (
            .O(N__35590),
            .I(N__35481));
    Span4Mux_h I__8815 (
            .O(N__35583),
            .I(N__35481));
    Span4Mux_h I__8814 (
            .O(N__35574),
            .I(N__35481));
    Span4Mux_s1_v I__8813 (
            .O(N__35571),
            .I(N__35476));
    Span4Mux_h I__8812 (
            .O(N__35566),
            .I(N__35476));
    Span12Mux_h I__8811 (
            .O(N__35559),
            .I(N__35469));
    Span12Mux_v I__8810 (
            .O(N__35556),
            .I(N__35469));
    Sp12to4 I__8809 (
            .O(N__35549),
            .I(N__35469));
    LocalMux I__8808 (
            .O(N__35546),
            .I(\c0.n1686 ));
    LocalMux I__8807 (
            .O(N__35543),
            .I(\c0.n1686 ));
    LocalMux I__8806 (
            .O(N__35536),
            .I(\c0.n1686 ));
    LocalMux I__8805 (
            .O(N__35529),
            .I(\c0.n1686 ));
    LocalMux I__8804 (
            .O(N__35524),
            .I(\c0.n1686 ));
    LocalMux I__8803 (
            .O(N__35517),
            .I(\c0.n1686 ));
    LocalMux I__8802 (
            .O(N__35512),
            .I(\c0.n1686 ));
    LocalMux I__8801 (
            .O(N__35509),
            .I(\c0.n1686 ));
    Odrv4 I__8800 (
            .O(N__35506),
            .I(\c0.n1686 ));
    Odrv4 I__8799 (
            .O(N__35503),
            .I(\c0.n1686 ));
    Odrv4 I__8798 (
            .O(N__35494),
            .I(\c0.n1686 ));
    Odrv4 I__8797 (
            .O(N__35481),
            .I(\c0.n1686 ));
    Odrv4 I__8796 (
            .O(N__35476),
            .I(\c0.n1686 ));
    Odrv12 I__8795 (
            .O(N__35469),
            .I(\c0.n1686 ));
    CascadeMux I__8794 (
            .O(N__35440),
            .I(N__35437));
    InMux I__8793 (
            .O(N__35437),
            .I(N__35434));
    LocalMux I__8792 (
            .O(N__35434),
            .I(N__35431));
    Span4Mux_s3_h I__8791 (
            .O(N__35431),
            .I(N__35428));
    Span4Mux_h I__8790 (
            .O(N__35428),
            .I(N__35425));
    Span4Mux_h I__8789 (
            .O(N__35425),
            .I(N__35421));
    InMux I__8788 (
            .O(N__35424),
            .I(N__35418));
    Span4Mux_h I__8787 (
            .O(N__35421),
            .I(N__35415));
    LocalMux I__8786 (
            .O(N__35418),
            .I(\c0.data_in_frame_19_4 ));
    Odrv4 I__8785 (
            .O(N__35415),
            .I(\c0.data_in_frame_19_4 ));
    ClkMux I__8784 (
            .O(N__35410),
            .I(N__34984));
    ClkMux I__8783 (
            .O(N__35409),
            .I(N__34984));
    ClkMux I__8782 (
            .O(N__35408),
            .I(N__34984));
    ClkMux I__8781 (
            .O(N__35407),
            .I(N__34984));
    ClkMux I__8780 (
            .O(N__35406),
            .I(N__34984));
    ClkMux I__8779 (
            .O(N__35405),
            .I(N__34984));
    ClkMux I__8778 (
            .O(N__35404),
            .I(N__34984));
    ClkMux I__8777 (
            .O(N__35403),
            .I(N__34984));
    ClkMux I__8776 (
            .O(N__35402),
            .I(N__34984));
    ClkMux I__8775 (
            .O(N__35401),
            .I(N__34984));
    ClkMux I__8774 (
            .O(N__35400),
            .I(N__34984));
    ClkMux I__8773 (
            .O(N__35399),
            .I(N__34984));
    ClkMux I__8772 (
            .O(N__35398),
            .I(N__34984));
    ClkMux I__8771 (
            .O(N__35397),
            .I(N__34984));
    ClkMux I__8770 (
            .O(N__35396),
            .I(N__34984));
    ClkMux I__8769 (
            .O(N__35395),
            .I(N__34984));
    ClkMux I__8768 (
            .O(N__35394),
            .I(N__34984));
    ClkMux I__8767 (
            .O(N__35393),
            .I(N__34984));
    ClkMux I__8766 (
            .O(N__35392),
            .I(N__34984));
    ClkMux I__8765 (
            .O(N__35391),
            .I(N__34984));
    ClkMux I__8764 (
            .O(N__35390),
            .I(N__34984));
    ClkMux I__8763 (
            .O(N__35389),
            .I(N__34984));
    ClkMux I__8762 (
            .O(N__35388),
            .I(N__34984));
    ClkMux I__8761 (
            .O(N__35387),
            .I(N__34984));
    ClkMux I__8760 (
            .O(N__35386),
            .I(N__34984));
    ClkMux I__8759 (
            .O(N__35385),
            .I(N__34984));
    ClkMux I__8758 (
            .O(N__35384),
            .I(N__34984));
    ClkMux I__8757 (
            .O(N__35383),
            .I(N__34984));
    ClkMux I__8756 (
            .O(N__35382),
            .I(N__34984));
    ClkMux I__8755 (
            .O(N__35381),
            .I(N__34984));
    ClkMux I__8754 (
            .O(N__35380),
            .I(N__34984));
    ClkMux I__8753 (
            .O(N__35379),
            .I(N__34984));
    ClkMux I__8752 (
            .O(N__35378),
            .I(N__34984));
    ClkMux I__8751 (
            .O(N__35377),
            .I(N__34984));
    ClkMux I__8750 (
            .O(N__35376),
            .I(N__34984));
    ClkMux I__8749 (
            .O(N__35375),
            .I(N__34984));
    ClkMux I__8748 (
            .O(N__35374),
            .I(N__34984));
    ClkMux I__8747 (
            .O(N__35373),
            .I(N__34984));
    ClkMux I__8746 (
            .O(N__35372),
            .I(N__34984));
    ClkMux I__8745 (
            .O(N__35371),
            .I(N__34984));
    ClkMux I__8744 (
            .O(N__35370),
            .I(N__34984));
    ClkMux I__8743 (
            .O(N__35369),
            .I(N__34984));
    ClkMux I__8742 (
            .O(N__35368),
            .I(N__34984));
    ClkMux I__8741 (
            .O(N__35367),
            .I(N__34984));
    ClkMux I__8740 (
            .O(N__35366),
            .I(N__34984));
    ClkMux I__8739 (
            .O(N__35365),
            .I(N__34984));
    ClkMux I__8738 (
            .O(N__35364),
            .I(N__34984));
    ClkMux I__8737 (
            .O(N__35363),
            .I(N__34984));
    ClkMux I__8736 (
            .O(N__35362),
            .I(N__34984));
    ClkMux I__8735 (
            .O(N__35361),
            .I(N__34984));
    ClkMux I__8734 (
            .O(N__35360),
            .I(N__34984));
    ClkMux I__8733 (
            .O(N__35359),
            .I(N__34984));
    ClkMux I__8732 (
            .O(N__35358),
            .I(N__34984));
    ClkMux I__8731 (
            .O(N__35357),
            .I(N__34984));
    ClkMux I__8730 (
            .O(N__35356),
            .I(N__34984));
    ClkMux I__8729 (
            .O(N__35355),
            .I(N__34984));
    ClkMux I__8728 (
            .O(N__35354),
            .I(N__34984));
    ClkMux I__8727 (
            .O(N__35353),
            .I(N__34984));
    ClkMux I__8726 (
            .O(N__35352),
            .I(N__34984));
    ClkMux I__8725 (
            .O(N__35351),
            .I(N__34984));
    ClkMux I__8724 (
            .O(N__35350),
            .I(N__34984));
    ClkMux I__8723 (
            .O(N__35349),
            .I(N__34984));
    ClkMux I__8722 (
            .O(N__35348),
            .I(N__34984));
    ClkMux I__8721 (
            .O(N__35347),
            .I(N__34984));
    ClkMux I__8720 (
            .O(N__35346),
            .I(N__34984));
    ClkMux I__8719 (
            .O(N__35345),
            .I(N__34984));
    ClkMux I__8718 (
            .O(N__35344),
            .I(N__34984));
    ClkMux I__8717 (
            .O(N__35343),
            .I(N__34984));
    ClkMux I__8716 (
            .O(N__35342),
            .I(N__34984));
    ClkMux I__8715 (
            .O(N__35341),
            .I(N__34984));
    ClkMux I__8714 (
            .O(N__35340),
            .I(N__34984));
    ClkMux I__8713 (
            .O(N__35339),
            .I(N__34984));
    ClkMux I__8712 (
            .O(N__35338),
            .I(N__34984));
    ClkMux I__8711 (
            .O(N__35337),
            .I(N__34984));
    ClkMux I__8710 (
            .O(N__35336),
            .I(N__34984));
    ClkMux I__8709 (
            .O(N__35335),
            .I(N__34984));
    ClkMux I__8708 (
            .O(N__35334),
            .I(N__34984));
    ClkMux I__8707 (
            .O(N__35333),
            .I(N__34984));
    ClkMux I__8706 (
            .O(N__35332),
            .I(N__34984));
    ClkMux I__8705 (
            .O(N__35331),
            .I(N__34984));
    ClkMux I__8704 (
            .O(N__35330),
            .I(N__34984));
    ClkMux I__8703 (
            .O(N__35329),
            .I(N__34984));
    ClkMux I__8702 (
            .O(N__35328),
            .I(N__34984));
    ClkMux I__8701 (
            .O(N__35327),
            .I(N__34984));
    ClkMux I__8700 (
            .O(N__35326),
            .I(N__34984));
    ClkMux I__8699 (
            .O(N__35325),
            .I(N__34984));
    ClkMux I__8698 (
            .O(N__35324),
            .I(N__34984));
    ClkMux I__8697 (
            .O(N__35323),
            .I(N__34984));
    ClkMux I__8696 (
            .O(N__35322),
            .I(N__34984));
    ClkMux I__8695 (
            .O(N__35321),
            .I(N__34984));
    ClkMux I__8694 (
            .O(N__35320),
            .I(N__34984));
    ClkMux I__8693 (
            .O(N__35319),
            .I(N__34984));
    ClkMux I__8692 (
            .O(N__35318),
            .I(N__34984));
    ClkMux I__8691 (
            .O(N__35317),
            .I(N__34984));
    ClkMux I__8690 (
            .O(N__35316),
            .I(N__34984));
    ClkMux I__8689 (
            .O(N__35315),
            .I(N__34984));
    ClkMux I__8688 (
            .O(N__35314),
            .I(N__34984));
    ClkMux I__8687 (
            .O(N__35313),
            .I(N__34984));
    ClkMux I__8686 (
            .O(N__35312),
            .I(N__34984));
    ClkMux I__8685 (
            .O(N__35311),
            .I(N__34984));
    ClkMux I__8684 (
            .O(N__35310),
            .I(N__34984));
    ClkMux I__8683 (
            .O(N__35309),
            .I(N__34984));
    ClkMux I__8682 (
            .O(N__35308),
            .I(N__34984));
    ClkMux I__8681 (
            .O(N__35307),
            .I(N__34984));
    ClkMux I__8680 (
            .O(N__35306),
            .I(N__34984));
    ClkMux I__8679 (
            .O(N__35305),
            .I(N__34984));
    ClkMux I__8678 (
            .O(N__35304),
            .I(N__34984));
    ClkMux I__8677 (
            .O(N__35303),
            .I(N__34984));
    ClkMux I__8676 (
            .O(N__35302),
            .I(N__34984));
    ClkMux I__8675 (
            .O(N__35301),
            .I(N__34984));
    ClkMux I__8674 (
            .O(N__35300),
            .I(N__34984));
    ClkMux I__8673 (
            .O(N__35299),
            .I(N__34984));
    ClkMux I__8672 (
            .O(N__35298),
            .I(N__34984));
    ClkMux I__8671 (
            .O(N__35297),
            .I(N__34984));
    ClkMux I__8670 (
            .O(N__35296),
            .I(N__34984));
    ClkMux I__8669 (
            .O(N__35295),
            .I(N__34984));
    ClkMux I__8668 (
            .O(N__35294),
            .I(N__34984));
    ClkMux I__8667 (
            .O(N__35293),
            .I(N__34984));
    ClkMux I__8666 (
            .O(N__35292),
            .I(N__34984));
    ClkMux I__8665 (
            .O(N__35291),
            .I(N__34984));
    ClkMux I__8664 (
            .O(N__35290),
            .I(N__34984));
    ClkMux I__8663 (
            .O(N__35289),
            .I(N__34984));
    ClkMux I__8662 (
            .O(N__35288),
            .I(N__34984));
    ClkMux I__8661 (
            .O(N__35287),
            .I(N__34984));
    ClkMux I__8660 (
            .O(N__35286),
            .I(N__34984));
    ClkMux I__8659 (
            .O(N__35285),
            .I(N__34984));
    ClkMux I__8658 (
            .O(N__35284),
            .I(N__34984));
    ClkMux I__8657 (
            .O(N__35283),
            .I(N__34984));
    ClkMux I__8656 (
            .O(N__35282),
            .I(N__34984));
    ClkMux I__8655 (
            .O(N__35281),
            .I(N__34984));
    ClkMux I__8654 (
            .O(N__35280),
            .I(N__34984));
    ClkMux I__8653 (
            .O(N__35279),
            .I(N__34984));
    ClkMux I__8652 (
            .O(N__35278),
            .I(N__34984));
    ClkMux I__8651 (
            .O(N__35277),
            .I(N__34984));
    ClkMux I__8650 (
            .O(N__35276),
            .I(N__34984));
    ClkMux I__8649 (
            .O(N__35275),
            .I(N__34984));
    ClkMux I__8648 (
            .O(N__35274),
            .I(N__34984));
    ClkMux I__8647 (
            .O(N__35273),
            .I(N__34984));
    ClkMux I__8646 (
            .O(N__35272),
            .I(N__34984));
    ClkMux I__8645 (
            .O(N__35271),
            .I(N__34984));
    ClkMux I__8644 (
            .O(N__35270),
            .I(N__34984));
    ClkMux I__8643 (
            .O(N__35269),
            .I(N__34984));
    GlobalMux I__8642 (
            .O(N__34984),
            .I(N__34981));
    gio2CtrlBuf I__8641 (
            .O(N__34981),
            .I(CLK_c));
    InMux I__8640 (
            .O(N__34978),
            .I(N__34975));
    LocalMux I__8639 (
            .O(N__34975),
            .I(n13));
    InMux I__8638 (
            .O(N__34972),
            .I(n4449));
    InMux I__8637 (
            .O(N__34969),
            .I(N__34966));
    LocalMux I__8636 (
            .O(N__34966),
            .I(n12));
    InMux I__8635 (
            .O(N__34963),
            .I(n4450));
    InMux I__8634 (
            .O(N__34960),
            .I(N__34957));
    LocalMux I__8633 (
            .O(N__34957),
            .I(n11));
    InMux I__8632 (
            .O(N__34954),
            .I(n4451));
    InMux I__8631 (
            .O(N__34951),
            .I(N__34948));
    LocalMux I__8630 (
            .O(N__34948),
            .I(n10));
    InMux I__8629 (
            .O(N__34945),
            .I(bfn_15_27_0_));
    InMux I__8628 (
            .O(N__34942),
            .I(N__34939));
    LocalMux I__8627 (
            .O(N__34939),
            .I(n9));
    InMux I__8626 (
            .O(N__34936),
            .I(n4453));
    InMux I__8625 (
            .O(N__34933),
            .I(N__34930));
    LocalMux I__8624 (
            .O(N__34930),
            .I(n8_adj_1989));
    InMux I__8623 (
            .O(N__34927),
            .I(n4454));
    InMux I__8622 (
            .O(N__34924),
            .I(N__34921));
    LocalMux I__8621 (
            .O(N__34921),
            .I(n7));
    InMux I__8620 (
            .O(N__34918),
            .I(n4455));
    InMux I__8619 (
            .O(N__34915),
            .I(N__34912));
    LocalMux I__8618 (
            .O(N__34912),
            .I(n6));
    InMux I__8617 (
            .O(N__34909),
            .I(n4456));
    InMux I__8616 (
            .O(N__34906),
            .I(N__34903));
    LocalMux I__8615 (
            .O(N__34903),
            .I(n21));
    InMux I__8614 (
            .O(N__34900),
            .I(n4441));
    InMux I__8613 (
            .O(N__34897),
            .I(N__34894));
    LocalMux I__8612 (
            .O(N__34894),
            .I(n20));
    InMux I__8611 (
            .O(N__34891),
            .I(n4442));
    InMux I__8610 (
            .O(N__34888),
            .I(N__34885));
    LocalMux I__8609 (
            .O(N__34885),
            .I(n19));
    InMux I__8608 (
            .O(N__34882),
            .I(n4443));
    InMux I__8607 (
            .O(N__34879),
            .I(N__34876));
    LocalMux I__8606 (
            .O(N__34876),
            .I(n18));
    InMux I__8605 (
            .O(N__34873),
            .I(bfn_15_26_0_));
    InMux I__8604 (
            .O(N__34870),
            .I(N__34867));
    LocalMux I__8603 (
            .O(N__34867),
            .I(n17));
    InMux I__8602 (
            .O(N__34864),
            .I(n4445));
    InMux I__8601 (
            .O(N__34861),
            .I(N__34858));
    LocalMux I__8600 (
            .O(N__34858),
            .I(n16));
    InMux I__8599 (
            .O(N__34855),
            .I(n4446));
    InMux I__8598 (
            .O(N__34852),
            .I(N__34849));
    LocalMux I__8597 (
            .O(N__34849),
            .I(n15));
    InMux I__8596 (
            .O(N__34846),
            .I(n4447));
    InMux I__8595 (
            .O(N__34843),
            .I(N__34840));
    LocalMux I__8594 (
            .O(N__34840),
            .I(n14));
    InMux I__8593 (
            .O(N__34837),
            .I(n4448));
    CascadeMux I__8592 (
            .O(N__34834),
            .I(\c0.n5887_cascade_ ));
    InMux I__8591 (
            .O(N__34831),
            .I(N__34822));
    InMux I__8590 (
            .O(N__34830),
            .I(N__34822));
    InMux I__8589 (
            .O(N__34829),
            .I(N__34817));
    InMux I__8588 (
            .O(N__34828),
            .I(N__34814));
    CascadeMux I__8587 (
            .O(N__34827),
            .I(N__34808));
    LocalMux I__8586 (
            .O(N__34822),
            .I(N__34801));
    InMux I__8585 (
            .O(N__34821),
            .I(N__34797));
    InMux I__8584 (
            .O(N__34820),
            .I(N__34794));
    LocalMux I__8583 (
            .O(N__34817),
            .I(N__34789));
    LocalMux I__8582 (
            .O(N__34814),
            .I(N__34789));
    InMux I__8581 (
            .O(N__34813),
            .I(N__34786));
    InMux I__8580 (
            .O(N__34812),
            .I(N__34783));
    InMux I__8579 (
            .O(N__34811),
            .I(N__34778));
    InMux I__8578 (
            .O(N__34808),
            .I(N__34778));
    InMux I__8577 (
            .O(N__34807),
            .I(N__34775));
    InMux I__8576 (
            .O(N__34806),
            .I(N__34772));
    InMux I__8575 (
            .O(N__34805),
            .I(N__34769));
    InMux I__8574 (
            .O(N__34804),
            .I(N__34766));
    Span4Mux_v I__8573 (
            .O(N__34801),
            .I(N__34763));
    CascadeMux I__8572 (
            .O(N__34800),
            .I(N__34758));
    LocalMux I__8571 (
            .O(N__34797),
            .I(N__34755));
    LocalMux I__8570 (
            .O(N__34794),
            .I(N__34748));
    Span4Mux_h I__8569 (
            .O(N__34789),
            .I(N__34748));
    LocalMux I__8568 (
            .O(N__34786),
            .I(N__34748));
    LocalMux I__8567 (
            .O(N__34783),
            .I(N__34744));
    LocalMux I__8566 (
            .O(N__34778),
            .I(N__34735));
    LocalMux I__8565 (
            .O(N__34775),
            .I(N__34735));
    LocalMux I__8564 (
            .O(N__34772),
            .I(N__34735));
    LocalMux I__8563 (
            .O(N__34769),
            .I(N__34735));
    LocalMux I__8562 (
            .O(N__34766),
            .I(N__34730));
    Span4Mux_h I__8561 (
            .O(N__34763),
            .I(N__34730));
    InMux I__8560 (
            .O(N__34762),
            .I(N__34727));
    InMux I__8559 (
            .O(N__34761),
            .I(N__34722));
    InMux I__8558 (
            .O(N__34758),
            .I(N__34722));
    Span4Mux_s3_h I__8557 (
            .O(N__34755),
            .I(N__34717));
    Span4Mux_h I__8556 (
            .O(N__34748),
            .I(N__34717));
    InMux I__8555 (
            .O(N__34747),
            .I(N__34714));
    Span4Mux_h I__8554 (
            .O(N__34744),
            .I(N__34707));
    Span4Mux_v I__8553 (
            .O(N__34735),
            .I(N__34707));
    Span4Mux_h I__8552 (
            .O(N__34730),
            .I(N__34707));
    LocalMux I__8551 (
            .O(N__34727),
            .I(\c0.byte_transmit_counter2_3 ));
    LocalMux I__8550 (
            .O(N__34722),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__8549 (
            .O(N__34717),
            .I(\c0.byte_transmit_counter2_3 ));
    LocalMux I__8548 (
            .O(N__34714),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__8547 (
            .O(N__34707),
            .I(\c0.byte_transmit_counter2_3 ));
    InMux I__8546 (
            .O(N__34696),
            .I(N__34693));
    LocalMux I__8545 (
            .O(N__34693),
            .I(N__34690));
    Span12Mux_h I__8544 (
            .O(N__34690),
            .I(N__34687));
    Odrv12 I__8543 (
            .O(N__34687),
            .I(\c0.n5890 ));
    InMux I__8542 (
            .O(N__34684),
            .I(N__34681));
    LocalMux I__8541 (
            .O(N__34681),
            .I(N__34677));
    InMux I__8540 (
            .O(N__34680),
            .I(N__34674));
    Span4Mux_h I__8539 (
            .O(N__34677),
            .I(N__34671));
    LocalMux I__8538 (
            .O(N__34674),
            .I(N__34668));
    Span4Mux_h I__8537 (
            .O(N__34671),
            .I(N__34664));
    Span4Mux_h I__8536 (
            .O(N__34668),
            .I(N__34661));
    InMux I__8535 (
            .O(N__34667),
            .I(N__34658));
    Odrv4 I__8534 (
            .O(N__34664),
            .I(\c0.n5219 ));
    Odrv4 I__8533 (
            .O(N__34661),
            .I(\c0.n5219 ));
    LocalMux I__8532 (
            .O(N__34658),
            .I(\c0.n5219 ));
    InMux I__8531 (
            .O(N__34651),
            .I(N__34648));
    LocalMux I__8530 (
            .O(N__34648),
            .I(N__34644));
    InMux I__8529 (
            .O(N__34647),
            .I(N__34641));
    Odrv4 I__8528 (
            .O(N__34644),
            .I(\c0.n5138 ));
    LocalMux I__8527 (
            .O(N__34641),
            .I(\c0.n5138 ));
    CascadeMux I__8526 (
            .O(N__34636),
            .I(N__34633));
    InMux I__8525 (
            .O(N__34633),
            .I(N__34630));
    LocalMux I__8524 (
            .O(N__34630),
            .I(N__34627));
    Span4Mux_h I__8523 (
            .O(N__34627),
            .I(N__34624));
    Span4Mux_h I__8522 (
            .O(N__34624),
            .I(N__34621));
    Odrv4 I__8521 (
            .O(N__34621),
            .I(\c0.n1896 ));
    InMux I__8520 (
            .O(N__34618),
            .I(N__34614));
    CascadeMux I__8519 (
            .O(N__34617),
            .I(N__34610));
    LocalMux I__8518 (
            .O(N__34614),
            .I(N__34607));
    InMux I__8517 (
            .O(N__34613),
            .I(N__34604));
    InMux I__8516 (
            .O(N__34610),
            .I(N__34601));
    Span4Mux_h I__8515 (
            .O(N__34607),
            .I(N__34598));
    LocalMux I__8514 (
            .O(N__34604),
            .I(data_in_8_4));
    LocalMux I__8513 (
            .O(N__34601),
            .I(data_in_8_4));
    Odrv4 I__8512 (
            .O(N__34598),
            .I(data_in_8_4));
    CascadeMux I__8511 (
            .O(N__34591),
            .I(N__34588));
    InMux I__8510 (
            .O(N__34588),
            .I(N__34584));
    InMux I__8509 (
            .O(N__34587),
            .I(N__34581));
    LocalMux I__8508 (
            .O(N__34584),
            .I(N__34576));
    LocalMux I__8507 (
            .O(N__34581),
            .I(N__34576));
    Span4Mux_v I__8506 (
            .O(N__34576),
            .I(N__34573));
    Span4Mux_h I__8505 (
            .O(N__34573),
            .I(N__34569));
    InMux I__8504 (
            .O(N__34572),
            .I(N__34566));
    Odrv4 I__8503 (
            .O(N__34569),
            .I(data_in_7_4));
    LocalMux I__8502 (
            .O(N__34566),
            .I(data_in_7_4));
    CascadeMux I__8501 (
            .O(N__34561),
            .I(N__34554));
    InMux I__8500 (
            .O(N__34560),
            .I(N__34514));
    InMux I__8499 (
            .O(N__34559),
            .I(N__34514));
    InMux I__8498 (
            .O(N__34558),
            .I(N__34514));
    InMux I__8497 (
            .O(N__34557),
            .I(N__34514));
    InMux I__8496 (
            .O(N__34554),
            .I(N__34509));
    InMux I__8495 (
            .O(N__34553),
            .I(N__34509));
    InMux I__8494 (
            .O(N__34552),
            .I(N__34506));
    CascadeMux I__8493 (
            .O(N__34551),
            .I(N__34502));
    InMux I__8492 (
            .O(N__34550),
            .I(N__34487));
    InMux I__8491 (
            .O(N__34549),
            .I(N__34482));
    InMux I__8490 (
            .O(N__34548),
            .I(N__34482));
    CascadeMux I__8489 (
            .O(N__34547),
            .I(N__34479));
    CascadeMux I__8488 (
            .O(N__34546),
            .I(N__34475));
    InMux I__8487 (
            .O(N__34545),
            .I(N__34468));
    InMux I__8486 (
            .O(N__34544),
            .I(N__34468));
    InMux I__8485 (
            .O(N__34543),
            .I(N__34461));
    InMux I__8484 (
            .O(N__34542),
            .I(N__34455));
    InMux I__8483 (
            .O(N__34541),
            .I(N__34452));
    InMux I__8482 (
            .O(N__34540),
            .I(N__34441));
    InMux I__8481 (
            .O(N__34539),
            .I(N__34441));
    InMux I__8480 (
            .O(N__34538),
            .I(N__34438));
    CascadeMux I__8479 (
            .O(N__34537),
            .I(N__34435));
    CascadeMux I__8478 (
            .O(N__34536),
            .I(N__34432));
    CascadeMux I__8477 (
            .O(N__34535),
            .I(N__34418));
    CascadeMux I__8476 (
            .O(N__34534),
            .I(N__34409));
    InMux I__8475 (
            .O(N__34533),
            .I(N__34403));
    InMux I__8474 (
            .O(N__34532),
            .I(N__34398));
    InMux I__8473 (
            .O(N__34531),
            .I(N__34398));
    InMux I__8472 (
            .O(N__34530),
            .I(N__34391));
    InMux I__8471 (
            .O(N__34529),
            .I(N__34391));
    InMux I__8470 (
            .O(N__34528),
            .I(N__34391));
    InMux I__8469 (
            .O(N__34527),
            .I(N__34386));
    InMux I__8468 (
            .O(N__34526),
            .I(N__34386));
    InMux I__8467 (
            .O(N__34525),
            .I(N__34383));
    InMux I__8466 (
            .O(N__34524),
            .I(N__34380));
    InMux I__8465 (
            .O(N__34523),
            .I(N__34375));
    LocalMux I__8464 (
            .O(N__34514),
            .I(N__34368));
    LocalMux I__8463 (
            .O(N__34509),
            .I(N__34368));
    LocalMux I__8462 (
            .O(N__34506),
            .I(N__34368));
    CascadeMux I__8461 (
            .O(N__34505),
            .I(N__34364));
    InMux I__8460 (
            .O(N__34502),
            .I(N__34354));
    InMux I__8459 (
            .O(N__34501),
            .I(N__34354));
    InMux I__8458 (
            .O(N__34500),
            .I(N__34354));
    InMux I__8457 (
            .O(N__34499),
            .I(N__34349));
    InMux I__8456 (
            .O(N__34498),
            .I(N__34349));
    InMux I__8455 (
            .O(N__34497),
            .I(N__34342));
    InMux I__8454 (
            .O(N__34496),
            .I(N__34342));
    InMux I__8453 (
            .O(N__34495),
            .I(N__34342));
    InMux I__8452 (
            .O(N__34494),
            .I(N__34337));
    InMux I__8451 (
            .O(N__34493),
            .I(N__34337));
    InMux I__8450 (
            .O(N__34492),
            .I(N__34334));
    InMux I__8449 (
            .O(N__34491),
            .I(N__34329));
    InMux I__8448 (
            .O(N__34490),
            .I(N__34329));
    LocalMux I__8447 (
            .O(N__34487),
            .I(N__34324));
    LocalMux I__8446 (
            .O(N__34482),
            .I(N__34324));
    InMux I__8445 (
            .O(N__34479),
            .I(N__34321));
    InMux I__8444 (
            .O(N__34478),
            .I(N__34310));
    InMux I__8443 (
            .O(N__34475),
            .I(N__34310));
    InMux I__8442 (
            .O(N__34474),
            .I(N__34310));
    InMux I__8441 (
            .O(N__34473),
            .I(N__34310));
    LocalMux I__8440 (
            .O(N__34468),
            .I(N__34307));
    InMux I__8439 (
            .O(N__34467),
            .I(N__34302));
    InMux I__8438 (
            .O(N__34466),
            .I(N__34302));
    InMux I__8437 (
            .O(N__34465),
            .I(N__34297));
    InMux I__8436 (
            .O(N__34464),
            .I(N__34297));
    LocalMux I__8435 (
            .O(N__34461),
            .I(N__34291));
    InMux I__8434 (
            .O(N__34460),
            .I(N__34288));
    InMux I__8433 (
            .O(N__34459),
            .I(N__34273));
    InMux I__8432 (
            .O(N__34458),
            .I(N__34273));
    LocalMux I__8431 (
            .O(N__34455),
            .I(N__34268));
    LocalMux I__8430 (
            .O(N__34452),
            .I(N__34268));
    InMux I__8429 (
            .O(N__34451),
            .I(N__34263));
    InMux I__8428 (
            .O(N__34450),
            .I(N__34263));
    InMux I__8427 (
            .O(N__34449),
            .I(N__34260));
    InMux I__8426 (
            .O(N__34448),
            .I(N__34257));
    InMux I__8425 (
            .O(N__34447),
            .I(N__34252));
    InMux I__8424 (
            .O(N__34446),
            .I(N__34252));
    LocalMux I__8423 (
            .O(N__34441),
            .I(N__34247));
    LocalMux I__8422 (
            .O(N__34438),
            .I(N__34247));
    InMux I__8421 (
            .O(N__34435),
            .I(N__34232));
    InMux I__8420 (
            .O(N__34432),
            .I(N__34232));
    InMux I__8419 (
            .O(N__34431),
            .I(N__34232));
    InMux I__8418 (
            .O(N__34430),
            .I(N__34232));
    InMux I__8417 (
            .O(N__34429),
            .I(N__34232));
    InMux I__8416 (
            .O(N__34428),
            .I(N__34232));
    InMux I__8415 (
            .O(N__34427),
            .I(N__34232));
    InMux I__8414 (
            .O(N__34426),
            .I(N__34221));
    InMux I__8413 (
            .O(N__34425),
            .I(N__34221));
    InMux I__8412 (
            .O(N__34424),
            .I(N__34221));
    InMux I__8411 (
            .O(N__34423),
            .I(N__34221));
    InMux I__8410 (
            .O(N__34422),
            .I(N__34221));
    InMux I__8409 (
            .O(N__34421),
            .I(N__34212));
    InMux I__8408 (
            .O(N__34418),
            .I(N__34203));
    InMux I__8407 (
            .O(N__34417),
            .I(N__34203));
    InMux I__8406 (
            .O(N__34416),
            .I(N__34203));
    InMux I__8405 (
            .O(N__34415),
            .I(N__34203));
    InMux I__8404 (
            .O(N__34414),
            .I(N__34196));
    InMux I__8403 (
            .O(N__34413),
            .I(N__34196));
    InMux I__8402 (
            .O(N__34412),
            .I(N__34196));
    InMux I__8401 (
            .O(N__34409),
            .I(N__34189));
    InMux I__8400 (
            .O(N__34408),
            .I(N__34189));
    InMux I__8399 (
            .O(N__34407),
            .I(N__34189));
    InMux I__8398 (
            .O(N__34406),
            .I(N__34186));
    LocalMux I__8397 (
            .O(N__34403),
            .I(N__34181));
    LocalMux I__8396 (
            .O(N__34398),
            .I(N__34181));
    LocalMux I__8395 (
            .O(N__34391),
            .I(N__34172));
    LocalMux I__8394 (
            .O(N__34386),
            .I(N__34172));
    LocalMux I__8393 (
            .O(N__34383),
            .I(N__34172));
    LocalMux I__8392 (
            .O(N__34380),
            .I(N__34172));
    CascadeMux I__8391 (
            .O(N__34379),
            .I(N__34169));
    InMux I__8390 (
            .O(N__34378),
            .I(N__34163));
    LocalMux I__8389 (
            .O(N__34375),
            .I(N__34158));
    Span4Mux_v I__8388 (
            .O(N__34368),
            .I(N__34158));
    InMux I__8387 (
            .O(N__34367),
            .I(N__34153));
    InMux I__8386 (
            .O(N__34364),
            .I(N__34153));
    CascadeMux I__8385 (
            .O(N__34363),
            .I(N__34148));
    InMux I__8384 (
            .O(N__34362),
            .I(N__34142));
    InMux I__8383 (
            .O(N__34361),
            .I(N__34142));
    LocalMux I__8382 (
            .O(N__34354),
            .I(N__34135));
    LocalMux I__8381 (
            .O(N__34349),
            .I(N__34132));
    LocalMux I__8380 (
            .O(N__34342),
            .I(N__34127));
    LocalMux I__8379 (
            .O(N__34337),
            .I(N__34127));
    LocalMux I__8378 (
            .O(N__34334),
            .I(N__34118));
    LocalMux I__8377 (
            .O(N__34329),
            .I(N__34118));
    Span4Mux_h I__8376 (
            .O(N__34324),
            .I(N__34118));
    LocalMux I__8375 (
            .O(N__34321),
            .I(N__34118));
    InMux I__8374 (
            .O(N__34320),
            .I(N__34115));
    InMux I__8373 (
            .O(N__34319),
            .I(N__34112));
    LocalMux I__8372 (
            .O(N__34310),
            .I(N__34103));
    Span4Mux_v I__8371 (
            .O(N__34307),
            .I(N__34103));
    LocalMux I__8370 (
            .O(N__34302),
            .I(N__34103));
    LocalMux I__8369 (
            .O(N__34297),
            .I(N__34103));
    CascadeMux I__8368 (
            .O(N__34296),
            .I(N__34100));
    InMux I__8367 (
            .O(N__34295),
            .I(N__34095));
    InMux I__8366 (
            .O(N__34294),
            .I(N__34095));
    Span4Mux_h I__8365 (
            .O(N__34291),
            .I(N__34090));
    LocalMux I__8364 (
            .O(N__34288),
            .I(N__34090));
    InMux I__8363 (
            .O(N__34287),
            .I(N__34083));
    InMux I__8362 (
            .O(N__34286),
            .I(N__34083));
    InMux I__8361 (
            .O(N__34285),
            .I(N__34083));
    CascadeMux I__8360 (
            .O(N__34284),
            .I(N__34078));
    InMux I__8359 (
            .O(N__34283),
            .I(N__34068));
    InMux I__8358 (
            .O(N__34282),
            .I(N__34068));
    InMux I__8357 (
            .O(N__34281),
            .I(N__34061));
    InMux I__8356 (
            .O(N__34280),
            .I(N__34061));
    InMux I__8355 (
            .O(N__34279),
            .I(N__34061));
    InMux I__8354 (
            .O(N__34278),
            .I(N__34058));
    LocalMux I__8353 (
            .O(N__34273),
            .I(N__34051));
    Span4Mux_v I__8352 (
            .O(N__34268),
            .I(N__34051));
    LocalMux I__8351 (
            .O(N__34263),
            .I(N__34051));
    LocalMux I__8350 (
            .O(N__34260),
            .I(N__34038));
    LocalMux I__8349 (
            .O(N__34257),
            .I(N__34038));
    LocalMux I__8348 (
            .O(N__34252),
            .I(N__34038));
    Span4Mux_v I__8347 (
            .O(N__34247),
            .I(N__34038));
    LocalMux I__8346 (
            .O(N__34232),
            .I(N__34038));
    LocalMux I__8345 (
            .O(N__34221),
            .I(N__34038));
    InMux I__8344 (
            .O(N__34220),
            .I(N__34032));
    InMux I__8343 (
            .O(N__34219),
            .I(N__34026));
    InMux I__8342 (
            .O(N__34218),
            .I(N__34023));
    InMux I__8341 (
            .O(N__34217),
            .I(N__34016));
    InMux I__8340 (
            .O(N__34216),
            .I(N__34016));
    InMux I__8339 (
            .O(N__34215),
            .I(N__34016));
    LocalMux I__8338 (
            .O(N__34212),
            .I(N__34000));
    LocalMux I__8337 (
            .O(N__34203),
            .I(N__34000));
    LocalMux I__8336 (
            .O(N__34196),
            .I(N__34000));
    LocalMux I__8335 (
            .O(N__34189),
            .I(N__34000));
    LocalMux I__8334 (
            .O(N__34186),
            .I(N__33993));
    Span4Mux_h I__8333 (
            .O(N__34181),
            .I(N__33993));
    Span4Mux_v I__8332 (
            .O(N__34172),
            .I(N__33993));
    InMux I__8331 (
            .O(N__34169),
            .I(N__33988));
    InMux I__8330 (
            .O(N__34168),
            .I(N__33988));
    InMux I__8329 (
            .O(N__34167),
            .I(N__33983));
    InMux I__8328 (
            .O(N__34166),
            .I(N__33983));
    LocalMux I__8327 (
            .O(N__34163),
            .I(N__33976));
    Span4Mux_h I__8326 (
            .O(N__34158),
            .I(N__33976));
    LocalMux I__8325 (
            .O(N__34153),
            .I(N__33976));
    InMux I__8324 (
            .O(N__34152),
            .I(N__33973));
    InMux I__8323 (
            .O(N__34151),
            .I(N__33970));
    InMux I__8322 (
            .O(N__34148),
            .I(N__33967));
    InMux I__8321 (
            .O(N__34147),
            .I(N__33964));
    LocalMux I__8320 (
            .O(N__34142),
            .I(N__33961));
    InMux I__8319 (
            .O(N__34141),
            .I(N__33954));
    InMux I__8318 (
            .O(N__34140),
            .I(N__33954));
    InMux I__8317 (
            .O(N__34139),
            .I(N__33954));
    InMux I__8316 (
            .O(N__34138),
            .I(N__33951));
    Span4Mux_v I__8315 (
            .O(N__34135),
            .I(N__33948));
    IoSpan4Mux I__8314 (
            .O(N__34132),
            .I(N__33941));
    Span4Mux_v I__8313 (
            .O(N__34127),
            .I(N__33941));
    Span4Mux_v I__8312 (
            .O(N__34118),
            .I(N__33941));
    LocalMux I__8311 (
            .O(N__34115),
            .I(N__33934));
    LocalMux I__8310 (
            .O(N__34112),
            .I(N__33934));
    Span4Mux_v I__8309 (
            .O(N__34103),
            .I(N__33934));
    InMux I__8308 (
            .O(N__34100),
            .I(N__33931));
    LocalMux I__8307 (
            .O(N__34095),
            .I(N__33926));
    Span4Mux_v I__8306 (
            .O(N__34090),
            .I(N__33926));
    LocalMux I__8305 (
            .O(N__34083),
            .I(N__33923));
    InMux I__8304 (
            .O(N__34082),
            .I(N__33907));
    InMux I__8303 (
            .O(N__34081),
            .I(N__33907));
    InMux I__8302 (
            .O(N__34078),
            .I(N__33907));
    InMux I__8301 (
            .O(N__34077),
            .I(N__33907));
    InMux I__8300 (
            .O(N__34076),
            .I(N__33907));
    InMux I__8299 (
            .O(N__34075),
            .I(N__33904));
    InMux I__8298 (
            .O(N__34074),
            .I(N__33901));
    InMux I__8297 (
            .O(N__34073),
            .I(N__33898));
    LocalMux I__8296 (
            .O(N__34068),
            .I(N__33895));
    LocalMux I__8295 (
            .O(N__34061),
            .I(N__33886));
    LocalMux I__8294 (
            .O(N__34058),
            .I(N__33886));
    Span4Mux_h I__8293 (
            .O(N__34051),
            .I(N__33886));
    Span4Mux_v I__8292 (
            .O(N__34038),
            .I(N__33886));
    InMux I__8291 (
            .O(N__34037),
            .I(N__33865));
    InMux I__8290 (
            .O(N__34036),
            .I(N__33865));
    InMux I__8289 (
            .O(N__34035),
            .I(N__33865));
    LocalMux I__8288 (
            .O(N__34032),
            .I(N__33862));
    InMux I__8287 (
            .O(N__34031),
            .I(N__33855));
    InMux I__8286 (
            .O(N__34030),
            .I(N__33855));
    InMux I__8285 (
            .O(N__34029),
            .I(N__33855));
    LocalMux I__8284 (
            .O(N__34026),
            .I(N__33852));
    LocalMux I__8283 (
            .O(N__34023),
            .I(N__33847));
    LocalMux I__8282 (
            .O(N__34016),
            .I(N__33847));
    InMux I__8281 (
            .O(N__34015),
            .I(N__33842));
    InMux I__8280 (
            .O(N__34014),
            .I(N__33842));
    InMux I__8279 (
            .O(N__34013),
            .I(N__33837));
    InMux I__8278 (
            .O(N__34012),
            .I(N__33837));
    InMux I__8277 (
            .O(N__34011),
            .I(N__33830));
    InMux I__8276 (
            .O(N__34010),
            .I(N__33830));
    InMux I__8275 (
            .O(N__34009),
            .I(N__33830));
    Span4Mux_v I__8274 (
            .O(N__34000),
            .I(N__33827));
    Span4Mux_v I__8273 (
            .O(N__33993),
            .I(N__33824));
    LocalMux I__8272 (
            .O(N__33988),
            .I(N__33817));
    LocalMux I__8271 (
            .O(N__33983),
            .I(N__33817));
    Span4Mux_v I__8270 (
            .O(N__33976),
            .I(N__33817));
    LocalMux I__8269 (
            .O(N__33973),
            .I(N__33812));
    LocalMux I__8268 (
            .O(N__33970),
            .I(N__33812));
    LocalMux I__8267 (
            .O(N__33967),
            .I(N__33805));
    LocalMux I__8266 (
            .O(N__33964),
            .I(N__33805));
    Span4Mux_v I__8265 (
            .O(N__33961),
            .I(N__33805));
    LocalMux I__8264 (
            .O(N__33954),
            .I(N__33794));
    LocalMux I__8263 (
            .O(N__33951),
            .I(N__33794));
    Span4Mux_h I__8262 (
            .O(N__33948),
            .I(N__33794));
    Span4Mux_s0_v I__8261 (
            .O(N__33941),
            .I(N__33794));
    Span4Mux_v I__8260 (
            .O(N__33934),
            .I(N__33794));
    LocalMux I__8259 (
            .O(N__33931),
            .I(N__33787));
    Span4Mux_h I__8258 (
            .O(N__33926),
            .I(N__33787));
    Span4Mux_v I__8257 (
            .O(N__33923),
            .I(N__33787));
    InMux I__8256 (
            .O(N__33922),
            .I(N__33784));
    InMux I__8255 (
            .O(N__33921),
            .I(N__33775));
    InMux I__8254 (
            .O(N__33920),
            .I(N__33775));
    InMux I__8253 (
            .O(N__33919),
            .I(N__33775));
    InMux I__8252 (
            .O(N__33918),
            .I(N__33775));
    LocalMux I__8251 (
            .O(N__33907),
            .I(N__33764));
    LocalMux I__8250 (
            .O(N__33904),
            .I(N__33764));
    LocalMux I__8249 (
            .O(N__33901),
            .I(N__33764));
    LocalMux I__8248 (
            .O(N__33898),
            .I(N__33764));
    Sp12to4 I__8247 (
            .O(N__33895),
            .I(N__33764));
    Span4Mux_v I__8246 (
            .O(N__33886),
            .I(N__33761));
    InMux I__8245 (
            .O(N__33885),
            .I(N__33758));
    InMux I__8244 (
            .O(N__33884),
            .I(N__33753));
    InMux I__8243 (
            .O(N__33883),
            .I(N__33753));
    InMux I__8242 (
            .O(N__33882),
            .I(N__33746));
    InMux I__8241 (
            .O(N__33881),
            .I(N__33746));
    InMux I__8240 (
            .O(N__33880),
            .I(N__33746));
    InMux I__8239 (
            .O(N__33879),
            .I(N__33739));
    InMux I__8238 (
            .O(N__33878),
            .I(N__33739));
    InMux I__8237 (
            .O(N__33877),
            .I(N__33739));
    InMux I__8236 (
            .O(N__33876),
            .I(N__33734));
    InMux I__8235 (
            .O(N__33875),
            .I(N__33734));
    InMux I__8234 (
            .O(N__33874),
            .I(N__33727));
    InMux I__8233 (
            .O(N__33873),
            .I(N__33727));
    InMux I__8232 (
            .O(N__33872),
            .I(N__33727));
    LocalMux I__8231 (
            .O(N__33865),
            .I(N__33724));
    Span4Mux_h I__8230 (
            .O(N__33862),
            .I(N__33721));
    LocalMux I__8229 (
            .O(N__33855),
            .I(N__33714));
    Span4Mux_v I__8228 (
            .O(N__33852),
            .I(N__33714));
    Span4Mux_v I__8227 (
            .O(N__33847),
            .I(N__33714));
    LocalMux I__8226 (
            .O(N__33842),
            .I(N__33701));
    LocalMux I__8225 (
            .O(N__33837),
            .I(N__33701));
    LocalMux I__8224 (
            .O(N__33830),
            .I(N__33701));
    Span4Mux_h I__8223 (
            .O(N__33827),
            .I(N__33701));
    Span4Mux_h I__8222 (
            .O(N__33824),
            .I(N__33701));
    Span4Mux_v I__8221 (
            .O(N__33817),
            .I(N__33701));
    Span4Mux_v I__8220 (
            .O(N__33812),
            .I(N__33692));
    Span4Mux_v I__8219 (
            .O(N__33805),
            .I(N__33692));
    Span4Mux_h I__8218 (
            .O(N__33794),
            .I(N__33692));
    Span4Mux_v I__8217 (
            .O(N__33787),
            .I(N__33692));
    LocalMux I__8216 (
            .O(N__33784),
            .I(N__33683));
    LocalMux I__8215 (
            .O(N__33775),
            .I(N__33683));
    Span12Mux_v I__8214 (
            .O(N__33764),
            .I(N__33683));
    Sp12to4 I__8213 (
            .O(N__33761),
            .I(N__33683));
    LocalMux I__8212 (
            .O(N__33758),
            .I(rx_data_ready));
    LocalMux I__8211 (
            .O(N__33753),
            .I(rx_data_ready));
    LocalMux I__8210 (
            .O(N__33746),
            .I(rx_data_ready));
    LocalMux I__8209 (
            .O(N__33739),
            .I(rx_data_ready));
    LocalMux I__8208 (
            .O(N__33734),
            .I(rx_data_ready));
    LocalMux I__8207 (
            .O(N__33727),
            .I(rx_data_ready));
    Odrv4 I__8206 (
            .O(N__33724),
            .I(rx_data_ready));
    Odrv4 I__8205 (
            .O(N__33721),
            .I(rx_data_ready));
    Odrv4 I__8204 (
            .O(N__33714),
            .I(rx_data_ready));
    Odrv4 I__8203 (
            .O(N__33701),
            .I(rx_data_ready));
    Odrv4 I__8202 (
            .O(N__33692),
            .I(rx_data_ready));
    Odrv12 I__8201 (
            .O(N__33683),
            .I(rx_data_ready));
    InMux I__8200 (
            .O(N__33658),
            .I(N__33655));
    LocalMux I__8199 (
            .O(N__33655),
            .I(N__33652));
    Span4Mux_h I__8198 (
            .O(N__33652),
            .I(N__33647));
    InMux I__8197 (
            .O(N__33651),
            .I(N__33644));
    InMux I__8196 (
            .O(N__33650),
            .I(N__33641));
    Odrv4 I__8195 (
            .O(N__33647),
            .I(data_in_17_2));
    LocalMux I__8194 (
            .O(N__33644),
            .I(data_in_17_2));
    LocalMux I__8193 (
            .O(N__33641),
            .I(data_in_17_2));
    CascadeMux I__8192 (
            .O(N__33634),
            .I(N__33631));
    InMux I__8191 (
            .O(N__33631),
            .I(N__33627));
    InMux I__8190 (
            .O(N__33630),
            .I(N__33624));
    LocalMux I__8189 (
            .O(N__33627),
            .I(N__33619));
    LocalMux I__8188 (
            .O(N__33624),
            .I(N__33619));
    Span4Mux_v I__8187 (
            .O(N__33619),
            .I(N__33616));
    Span4Mux_h I__8186 (
            .O(N__33616),
            .I(N__33612));
    InMux I__8185 (
            .O(N__33615),
            .I(N__33609));
    Odrv4 I__8184 (
            .O(N__33612),
            .I(data_in_16_2));
    LocalMux I__8183 (
            .O(N__33609),
            .I(data_in_16_2));
    InMux I__8182 (
            .O(N__33604),
            .I(N__33601));
    LocalMux I__8181 (
            .O(N__33601),
            .I(n26));
    InMux I__8180 (
            .O(N__33598),
            .I(bfn_15_25_0_));
    InMux I__8179 (
            .O(N__33595),
            .I(N__33592));
    LocalMux I__8178 (
            .O(N__33592),
            .I(n25));
    InMux I__8177 (
            .O(N__33589),
            .I(n4437));
    InMux I__8176 (
            .O(N__33586),
            .I(N__33583));
    LocalMux I__8175 (
            .O(N__33583),
            .I(n24));
    InMux I__8174 (
            .O(N__33580),
            .I(n4438));
    InMux I__8173 (
            .O(N__33577),
            .I(N__33574));
    LocalMux I__8172 (
            .O(N__33574),
            .I(n23));
    InMux I__8171 (
            .O(N__33571),
            .I(n4439));
    InMux I__8170 (
            .O(N__33568),
            .I(N__33565));
    LocalMux I__8169 (
            .O(N__33565),
            .I(n22));
    InMux I__8168 (
            .O(N__33562),
            .I(n4440));
    CascadeMux I__8167 (
            .O(N__33559),
            .I(N__33555));
    InMux I__8166 (
            .O(N__33558),
            .I(N__33552));
    InMux I__8165 (
            .O(N__33555),
            .I(N__33548));
    LocalMux I__8164 (
            .O(N__33552),
            .I(N__33545));
    InMux I__8163 (
            .O(N__33551),
            .I(N__33542));
    LocalMux I__8162 (
            .O(N__33548),
            .I(data_in_9_2));
    Odrv12 I__8161 (
            .O(N__33545),
            .I(data_in_9_2));
    LocalMux I__8160 (
            .O(N__33542),
            .I(data_in_9_2));
    CascadeMux I__8159 (
            .O(N__33535),
            .I(N__33532));
    InMux I__8158 (
            .O(N__33532),
            .I(N__33528));
    InMux I__8157 (
            .O(N__33531),
            .I(N__33525));
    LocalMux I__8156 (
            .O(N__33528),
            .I(N__33522));
    LocalMux I__8155 (
            .O(N__33525),
            .I(N__33519));
    Span4Mux_h I__8154 (
            .O(N__33522),
            .I(N__33513));
    Span4Mux_h I__8153 (
            .O(N__33519),
            .I(N__33513));
    InMux I__8152 (
            .O(N__33518),
            .I(N__33510));
    Odrv4 I__8151 (
            .O(N__33513),
            .I(data_in_8_3));
    LocalMux I__8150 (
            .O(N__33510),
            .I(data_in_8_3));
    InMux I__8149 (
            .O(N__33505),
            .I(N__33502));
    LocalMux I__8148 (
            .O(N__33502),
            .I(N__33498));
    InMux I__8147 (
            .O(N__33501),
            .I(N__33495));
    Span4Mux_s1_v I__8146 (
            .O(N__33498),
            .I(N__33490));
    LocalMux I__8145 (
            .O(N__33495),
            .I(N__33490));
    Span4Mux_h I__8144 (
            .O(N__33490),
            .I(N__33486));
    InMux I__8143 (
            .O(N__33489),
            .I(N__33483));
    Odrv4 I__8142 (
            .O(N__33486),
            .I(data_in_7_3));
    LocalMux I__8141 (
            .O(N__33483),
            .I(data_in_7_3));
    InMux I__8140 (
            .O(N__33478),
            .I(N__33473));
    InMux I__8139 (
            .O(N__33477),
            .I(N__33470));
    CascadeMux I__8138 (
            .O(N__33476),
            .I(N__33467));
    LocalMux I__8137 (
            .O(N__33473),
            .I(N__33464));
    LocalMux I__8136 (
            .O(N__33470),
            .I(N__33461));
    InMux I__8135 (
            .O(N__33467),
            .I(N__33458));
    Span4Mux_h I__8134 (
            .O(N__33464),
            .I(N__33455));
    Span4Mux_h I__8133 (
            .O(N__33461),
            .I(N__33449));
    LocalMux I__8132 (
            .O(N__33458),
            .I(N__33449));
    Span4Mux_h I__8131 (
            .O(N__33455),
            .I(N__33446));
    InMux I__8130 (
            .O(N__33454),
            .I(N__33443));
    Span4Mux_v I__8129 (
            .O(N__33449),
            .I(N__33440));
    Odrv4 I__8128 (
            .O(N__33446),
            .I(data_in_18_0));
    LocalMux I__8127 (
            .O(N__33443),
            .I(data_in_18_0));
    Odrv4 I__8126 (
            .O(N__33440),
            .I(data_in_18_0));
    CascadeMux I__8125 (
            .O(N__33433),
            .I(N__33429));
    InMux I__8124 (
            .O(N__33432),
            .I(N__33426));
    InMux I__8123 (
            .O(N__33429),
            .I(N__33423));
    LocalMux I__8122 (
            .O(N__33426),
            .I(N__33420));
    LocalMux I__8121 (
            .O(N__33423),
            .I(N__33416));
    Span4Mux_v I__8120 (
            .O(N__33420),
            .I(N__33413));
    InMux I__8119 (
            .O(N__33419),
            .I(N__33410));
    Odrv4 I__8118 (
            .O(N__33416),
            .I(data_in_17_0));
    Odrv4 I__8117 (
            .O(N__33413),
            .I(data_in_17_0));
    LocalMux I__8116 (
            .O(N__33410),
            .I(data_in_17_0));
    InMux I__8115 (
            .O(N__33403),
            .I(N__33399));
    InMux I__8114 (
            .O(N__33402),
            .I(N__33395));
    LocalMux I__8113 (
            .O(N__33399),
            .I(N__33390));
    InMux I__8112 (
            .O(N__33398),
            .I(N__33387));
    LocalMux I__8111 (
            .O(N__33395),
            .I(N__33384));
    InMux I__8110 (
            .O(N__33394),
            .I(N__33381));
    InMux I__8109 (
            .O(N__33393),
            .I(N__33378));
    Span4Mux_h I__8108 (
            .O(N__33390),
            .I(N__33375));
    LocalMux I__8107 (
            .O(N__33387),
            .I(N__33368));
    Span4Mux_v I__8106 (
            .O(N__33384),
            .I(N__33368));
    LocalMux I__8105 (
            .O(N__33381),
            .I(N__33368));
    LocalMux I__8104 (
            .O(N__33378),
            .I(\c0.data_in_field_118 ));
    Odrv4 I__8103 (
            .O(N__33375),
            .I(\c0.data_in_field_118 ));
    Odrv4 I__8102 (
            .O(N__33368),
            .I(\c0.data_in_field_118 ));
    InMux I__8101 (
            .O(N__33361),
            .I(N__33356));
    CascadeMux I__8100 (
            .O(N__33360),
            .I(N__33353));
    InMux I__8099 (
            .O(N__33359),
            .I(N__33350));
    LocalMux I__8098 (
            .O(N__33356),
            .I(N__33347));
    InMux I__8097 (
            .O(N__33353),
            .I(N__33343));
    LocalMux I__8096 (
            .O(N__33350),
            .I(N__33340));
    Span12Mux_h I__8095 (
            .O(N__33347),
            .I(N__33336));
    InMux I__8094 (
            .O(N__33346),
            .I(N__33333));
    LocalMux I__8093 (
            .O(N__33343),
            .I(N__33328));
    Span4Mux_h I__8092 (
            .O(N__33340),
            .I(N__33328));
    InMux I__8091 (
            .O(N__33339),
            .I(N__33325));
    Odrv12 I__8090 (
            .O(N__33336),
            .I(\c0.data_in_field_126 ));
    LocalMux I__8089 (
            .O(N__33333),
            .I(\c0.data_in_field_126 ));
    Odrv4 I__8088 (
            .O(N__33328),
            .I(\c0.data_in_field_126 ));
    LocalMux I__8087 (
            .O(N__33325),
            .I(\c0.data_in_field_126 ));
    InMux I__8086 (
            .O(N__33316),
            .I(N__33312));
    InMux I__8085 (
            .O(N__33315),
            .I(N__33306));
    LocalMux I__8084 (
            .O(N__33312),
            .I(N__33303));
    InMux I__8083 (
            .O(N__33311),
            .I(N__33300));
    InMux I__8082 (
            .O(N__33310),
            .I(N__33295));
    InMux I__8081 (
            .O(N__33309),
            .I(N__33291));
    LocalMux I__8080 (
            .O(N__33306),
            .I(N__33282));
    Span4Mux_v I__8079 (
            .O(N__33303),
            .I(N__33277));
    LocalMux I__8078 (
            .O(N__33300),
            .I(N__33277));
    InMux I__8077 (
            .O(N__33299),
            .I(N__33267));
    InMux I__8076 (
            .O(N__33298),
            .I(N__33264));
    LocalMux I__8075 (
            .O(N__33295),
            .I(N__33260));
    InMux I__8074 (
            .O(N__33294),
            .I(N__33257));
    LocalMux I__8073 (
            .O(N__33291),
            .I(N__33253));
    InMux I__8072 (
            .O(N__33290),
            .I(N__33250));
    InMux I__8071 (
            .O(N__33289),
            .I(N__33247));
    InMux I__8070 (
            .O(N__33288),
            .I(N__33241));
    InMux I__8069 (
            .O(N__33287),
            .I(N__33241));
    InMux I__8068 (
            .O(N__33286),
            .I(N__33238));
    InMux I__8067 (
            .O(N__33285),
            .I(N__33233));
    Span4Mux_v I__8066 (
            .O(N__33282),
            .I(N__33228));
    Span4Mux_h I__8065 (
            .O(N__33277),
            .I(N__33228));
    InMux I__8064 (
            .O(N__33276),
            .I(N__33223));
    InMux I__8063 (
            .O(N__33275),
            .I(N__33223));
    InMux I__8062 (
            .O(N__33274),
            .I(N__33218));
    InMux I__8061 (
            .O(N__33273),
            .I(N__33213));
    InMux I__8060 (
            .O(N__33272),
            .I(N__33213));
    InMux I__8059 (
            .O(N__33271),
            .I(N__33209));
    InMux I__8058 (
            .O(N__33270),
            .I(N__33206));
    LocalMux I__8057 (
            .O(N__33267),
            .I(N__33203));
    LocalMux I__8056 (
            .O(N__33264),
            .I(N__33198));
    InMux I__8055 (
            .O(N__33263),
            .I(N__33195));
    Span4Mux_h I__8054 (
            .O(N__33260),
            .I(N__33190));
    LocalMux I__8053 (
            .O(N__33257),
            .I(N__33190));
    InMux I__8052 (
            .O(N__33256),
            .I(N__33187));
    Span4Mux_s2_v I__8051 (
            .O(N__33253),
            .I(N__33174));
    LocalMux I__8050 (
            .O(N__33250),
            .I(N__33174));
    LocalMux I__8049 (
            .O(N__33247),
            .I(N__33174));
    InMux I__8048 (
            .O(N__33246),
            .I(N__33171));
    LocalMux I__8047 (
            .O(N__33241),
            .I(N__33168));
    LocalMux I__8046 (
            .O(N__33238),
            .I(N__33165));
    InMux I__8045 (
            .O(N__33237),
            .I(N__33162));
    InMux I__8044 (
            .O(N__33236),
            .I(N__33159));
    LocalMux I__8043 (
            .O(N__33233),
            .I(N__33152));
    Span4Mux_h I__8042 (
            .O(N__33228),
            .I(N__33152));
    LocalMux I__8041 (
            .O(N__33223),
            .I(N__33152));
    InMux I__8040 (
            .O(N__33222),
            .I(N__33149));
    InMux I__8039 (
            .O(N__33221),
            .I(N__33146));
    LocalMux I__8038 (
            .O(N__33218),
            .I(N__33143));
    LocalMux I__8037 (
            .O(N__33213),
            .I(N__33140));
    InMux I__8036 (
            .O(N__33212),
            .I(N__33135));
    LocalMux I__8035 (
            .O(N__33209),
            .I(N__33128));
    LocalMux I__8034 (
            .O(N__33206),
            .I(N__33128));
    Span4Mux_v I__8033 (
            .O(N__33203),
            .I(N__33128));
    InMux I__8032 (
            .O(N__33202),
            .I(N__33123));
    InMux I__8031 (
            .O(N__33201),
            .I(N__33123));
    Span4Mux_v I__8030 (
            .O(N__33198),
            .I(N__33118));
    LocalMux I__8029 (
            .O(N__33195),
            .I(N__33118));
    Span4Mux_v I__8028 (
            .O(N__33190),
            .I(N__33112));
    LocalMux I__8027 (
            .O(N__33187),
            .I(N__33109));
    InMux I__8026 (
            .O(N__33186),
            .I(N__33104));
    InMux I__8025 (
            .O(N__33185),
            .I(N__33104));
    InMux I__8024 (
            .O(N__33184),
            .I(N__33101));
    InMux I__8023 (
            .O(N__33183),
            .I(N__33096));
    InMux I__8022 (
            .O(N__33182),
            .I(N__33096));
    InMux I__8021 (
            .O(N__33181),
            .I(N__33093));
    Span4Mux_v I__8020 (
            .O(N__33174),
            .I(N__33090));
    LocalMux I__8019 (
            .O(N__33171),
            .I(N__33079));
    Span4Mux_s2_h I__8018 (
            .O(N__33168),
            .I(N__33079));
    Span4Mux_h I__8017 (
            .O(N__33165),
            .I(N__33079));
    LocalMux I__8016 (
            .O(N__33162),
            .I(N__33079));
    LocalMux I__8015 (
            .O(N__33159),
            .I(N__33079));
    Span4Mux_v I__8014 (
            .O(N__33152),
            .I(N__33076));
    LocalMux I__8013 (
            .O(N__33149),
            .I(N__33067));
    LocalMux I__8012 (
            .O(N__33146),
            .I(N__33067));
    Span4Mux_h I__8011 (
            .O(N__33143),
            .I(N__33067));
    Span4Mux_v I__8010 (
            .O(N__33140),
            .I(N__33067));
    InMux I__8009 (
            .O(N__33139),
            .I(N__33062));
    InMux I__8008 (
            .O(N__33138),
            .I(N__33062));
    LocalMux I__8007 (
            .O(N__33135),
            .I(N__33053));
    Span4Mux_h I__8006 (
            .O(N__33128),
            .I(N__33053));
    LocalMux I__8005 (
            .O(N__33123),
            .I(N__33053));
    Span4Mux_v I__8004 (
            .O(N__33118),
            .I(N__33053));
    InMux I__8003 (
            .O(N__33117),
            .I(N__33050));
    InMux I__8002 (
            .O(N__33116),
            .I(N__33047));
    InMux I__8001 (
            .O(N__33115),
            .I(N__33044));
    Sp12to4 I__8000 (
            .O(N__33112),
            .I(N__33033));
    Span12Mux_s8_v I__7999 (
            .O(N__33109),
            .I(N__33033));
    LocalMux I__7998 (
            .O(N__33104),
            .I(N__33033));
    LocalMux I__7997 (
            .O(N__33101),
            .I(N__33033));
    LocalMux I__7996 (
            .O(N__33096),
            .I(N__33033));
    LocalMux I__7995 (
            .O(N__33093),
            .I(N__33024));
    Span4Mux_h I__7994 (
            .O(N__33090),
            .I(N__33024));
    Span4Mux_v I__7993 (
            .O(N__33079),
            .I(N__33024));
    Span4Mux_h I__7992 (
            .O(N__33076),
            .I(N__33024));
    Span4Mux_v I__7991 (
            .O(N__33067),
            .I(N__33017));
    LocalMux I__7990 (
            .O(N__33062),
            .I(N__33017));
    Span4Mux_h I__7989 (
            .O(N__33053),
            .I(N__33017));
    LocalMux I__7988 (
            .O(N__33050),
            .I(N__33014));
    LocalMux I__7987 (
            .O(N__33047),
            .I(\c0.byte_transmit_counter2_0 ));
    LocalMux I__7986 (
            .O(N__33044),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv12 I__7985 (
            .O(N__33033),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__7984 (
            .O(N__33024),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__7983 (
            .O(N__33017),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv12 I__7982 (
            .O(N__33014),
            .I(\c0.byte_transmit_counter2_0 ));
    InMux I__7981 (
            .O(N__33001),
            .I(N__32998));
    LocalMux I__7980 (
            .O(N__32998),
            .I(N__32995));
    Span4Mux_v I__7979 (
            .O(N__32995),
            .I(N__32991));
    CascadeMux I__7978 (
            .O(N__32994),
            .I(N__32987));
    Sp12to4 I__7977 (
            .O(N__32991),
            .I(N__32982));
    InMux I__7976 (
            .O(N__32990),
            .I(N__32979));
    InMux I__7975 (
            .O(N__32987),
            .I(N__32972));
    InMux I__7974 (
            .O(N__32986),
            .I(N__32972));
    InMux I__7973 (
            .O(N__32985),
            .I(N__32972));
    Odrv12 I__7972 (
            .O(N__32982),
            .I(\c0.data_in_field_86 ));
    LocalMux I__7971 (
            .O(N__32979),
            .I(\c0.data_in_field_86 ));
    LocalMux I__7970 (
            .O(N__32972),
            .I(\c0.data_in_field_86 ));
    InMux I__7969 (
            .O(N__32965),
            .I(N__32961));
    InMux I__7968 (
            .O(N__32964),
            .I(N__32957));
    LocalMux I__7967 (
            .O(N__32961),
            .I(N__32954));
    InMux I__7966 (
            .O(N__32960),
            .I(N__32951));
    LocalMux I__7965 (
            .O(N__32957),
            .I(N__32947));
    Span4Mux_v I__7964 (
            .O(N__32954),
            .I(N__32942));
    LocalMux I__7963 (
            .O(N__32951),
            .I(N__32942));
    CascadeMux I__7962 (
            .O(N__32950),
            .I(N__32939));
    Span4Mux_v I__7961 (
            .O(N__32947),
            .I(N__32933));
    Span4Mux_h I__7960 (
            .O(N__32942),
            .I(N__32933));
    InMux I__7959 (
            .O(N__32939),
            .I(N__32930));
    InMux I__7958 (
            .O(N__32938),
            .I(N__32927));
    Span4Mux_h I__7957 (
            .O(N__32933),
            .I(N__32924));
    LocalMux I__7956 (
            .O(N__32930),
            .I(N__32921));
    LocalMux I__7955 (
            .O(N__32927),
            .I(\c0.data_in_field_94 ));
    Odrv4 I__7954 (
            .O(N__32924),
            .I(\c0.data_in_field_94 ));
    Odrv4 I__7953 (
            .O(N__32921),
            .I(\c0.data_in_field_94 ));
    CascadeMux I__7952 (
            .O(N__32914),
            .I(N__32910));
    InMux I__7951 (
            .O(N__32913),
            .I(N__32906));
    InMux I__7950 (
            .O(N__32910),
            .I(N__32903));
    InMux I__7949 (
            .O(N__32909),
            .I(N__32900));
    LocalMux I__7948 (
            .O(N__32906),
            .I(N__32897));
    LocalMux I__7947 (
            .O(N__32903),
            .I(N__32894));
    LocalMux I__7946 (
            .O(N__32900),
            .I(N__32890));
    Span4Mux_v I__7945 (
            .O(N__32897),
            .I(N__32884));
    Span4Mux_v I__7944 (
            .O(N__32894),
            .I(N__32884));
    InMux I__7943 (
            .O(N__32893),
            .I(N__32881));
    Span4Mux_v I__7942 (
            .O(N__32890),
            .I(N__32878));
    InMux I__7941 (
            .O(N__32889),
            .I(N__32875));
    Sp12to4 I__7940 (
            .O(N__32884),
            .I(N__32872));
    LocalMux I__7939 (
            .O(N__32881),
            .I(\c0.data_in_field_70 ));
    Odrv4 I__7938 (
            .O(N__32878),
            .I(\c0.data_in_field_70 ));
    LocalMux I__7937 (
            .O(N__32875),
            .I(\c0.data_in_field_70 ));
    Odrv12 I__7936 (
            .O(N__32872),
            .I(\c0.data_in_field_70 ));
    CascadeMux I__7935 (
            .O(N__32863),
            .I(\c0.n5899_cascade_ ));
    InMux I__7934 (
            .O(N__32860),
            .I(N__32857));
    LocalMux I__7933 (
            .O(N__32857),
            .I(N__32854));
    Span4Mux_h I__7932 (
            .O(N__32854),
            .I(N__32849));
    InMux I__7931 (
            .O(N__32853),
            .I(N__32844));
    InMux I__7930 (
            .O(N__32852),
            .I(N__32844));
    Odrv4 I__7929 (
            .O(N__32849),
            .I(\c0.data_in_field_78 ));
    LocalMux I__7928 (
            .O(N__32844),
            .I(\c0.data_in_field_78 ));
    InMux I__7927 (
            .O(N__32839),
            .I(N__32836));
    LocalMux I__7926 (
            .O(N__32836),
            .I(N__32833));
    Odrv4 I__7925 (
            .O(N__32833),
            .I(\c0.n5893 ));
    InMux I__7924 (
            .O(N__32830),
            .I(N__32826));
    CascadeMux I__7923 (
            .O(N__32829),
            .I(N__32822));
    LocalMux I__7922 (
            .O(N__32826),
            .I(N__32819));
    InMux I__7921 (
            .O(N__32825),
            .I(N__32816));
    InMux I__7920 (
            .O(N__32822),
            .I(N__32813));
    Span4Mux_v I__7919 (
            .O(N__32819),
            .I(N__32810));
    LocalMux I__7918 (
            .O(N__32816),
            .I(N__32806));
    LocalMux I__7917 (
            .O(N__32813),
            .I(N__32801));
    Span4Mux_h I__7916 (
            .O(N__32810),
            .I(N__32801));
    InMux I__7915 (
            .O(N__32809),
            .I(N__32798));
    Odrv4 I__7914 (
            .O(N__32806),
            .I(\c0.data_in_field_102 ));
    Odrv4 I__7913 (
            .O(N__32801),
            .I(\c0.data_in_field_102 ));
    LocalMux I__7912 (
            .O(N__32798),
            .I(\c0.data_in_field_102 ));
    InMux I__7911 (
            .O(N__32791),
            .I(N__32786));
    CascadeMux I__7910 (
            .O(N__32790),
            .I(N__32782));
    CascadeMux I__7909 (
            .O(N__32789),
            .I(N__32779));
    LocalMux I__7908 (
            .O(N__32786),
            .I(N__32772));
    InMux I__7907 (
            .O(N__32785),
            .I(N__32769));
    InMux I__7906 (
            .O(N__32782),
            .I(N__32766));
    InMux I__7905 (
            .O(N__32779),
            .I(N__32763));
    CascadeMux I__7904 (
            .O(N__32778),
            .I(N__32760));
    CascadeMux I__7903 (
            .O(N__32777),
            .I(N__32757));
    InMux I__7902 (
            .O(N__32776),
            .I(N__32750));
    InMux I__7901 (
            .O(N__32775),
            .I(N__32750));
    Span4Mux_h I__7900 (
            .O(N__32772),
            .I(N__32741));
    LocalMux I__7899 (
            .O(N__32769),
            .I(N__32741));
    LocalMux I__7898 (
            .O(N__32766),
            .I(N__32741));
    LocalMux I__7897 (
            .O(N__32763),
            .I(N__32741));
    InMux I__7896 (
            .O(N__32760),
            .I(N__32736));
    InMux I__7895 (
            .O(N__32757),
            .I(N__32736));
    InMux I__7894 (
            .O(N__32756),
            .I(N__32730));
    InMux I__7893 (
            .O(N__32755),
            .I(N__32727));
    LocalMux I__7892 (
            .O(N__32750),
            .I(N__32720));
    Span4Mux_v I__7891 (
            .O(N__32741),
            .I(N__32720));
    LocalMux I__7890 (
            .O(N__32736),
            .I(N__32720));
    CascadeMux I__7889 (
            .O(N__32735),
            .I(N__32717));
    CascadeMux I__7888 (
            .O(N__32734),
            .I(N__32714));
    InMux I__7887 (
            .O(N__32733),
            .I(N__32709));
    LocalMux I__7886 (
            .O(N__32730),
            .I(N__32702));
    LocalMux I__7885 (
            .O(N__32727),
            .I(N__32702));
    Span4Mux_v I__7884 (
            .O(N__32720),
            .I(N__32702));
    InMux I__7883 (
            .O(N__32717),
            .I(N__32699));
    InMux I__7882 (
            .O(N__32714),
            .I(N__32691));
    InMux I__7881 (
            .O(N__32713),
            .I(N__32691));
    CascadeMux I__7880 (
            .O(N__32712),
            .I(N__32688));
    LocalMux I__7879 (
            .O(N__32709),
            .I(N__32685));
    Span4Mux_v I__7878 (
            .O(N__32702),
            .I(N__32680));
    LocalMux I__7877 (
            .O(N__32699),
            .I(N__32680));
    CascadeMux I__7876 (
            .O(N__32698),
            .I(N__32675));
    CascadeMux I__7875 (
            .O(N__32697),
            .I(N__32671));
    CascadeMux I__7874 (
            .O(N__32696),
            .I(N__32668));
    LocalMux I__7873 (
            .O(N__32691),
            .I(N__32663));
    InMux I__7872 (
            .O(N__32688),
            .I(N__32660));
    Span4Mux_s3_v I__7871 (
            .O(N__32685),
            .I(N__32652));
    Span4Mux_s3_v I__7870 (
            .O(N__32680),
            .I(N__32652));
    CascadeMux I__7869 (
            .O(N__32679),
            .I(N__32649));
    CascadeMux I__7868 (
            .O(N__32678),
            .I(N__32646));
    InMux I__7867 (
            .O(N__32675),
            .I(N__32643));
    InMux I__7866 (
            .O(N__32674),
            .I(N__32634));
    InMux I__7865 (
            .O(N__32671),
            .I(N__32634));
    InMux I__7864 (
            .O(N__32668),
            .I(N__32634));
    InMux I__7863 (
            .O(N__32667),
            .I(N__32634));
    CascadeMux I__7862 (
            .O(N__32666),
            .I(N__32631));
    Span4Mux_h I__7861 (
            .O(N__32663),
            .I(N__32622));
    LocalMux I__7860 (
            .O(N__32660),
            .I(N__32622));
    InMux I__7859 (
            .O(N__32659),
            .I(N__32619));
    CascadeMux I__7858 (
            .O(N__32658),
            .I(N__32616));
    InMux I__7857 (
            .O(N__32657),
            .I(N__32613));
    Span4Mux_h I__7856 (
            .O(N__32652),
            .I(N__32610));
    InMux I__7855 (
            .O(N__32649),
            .I(N__32607));
    InMux I__7854 (
            .O(N__32646),
            .I(N__32604));
    LocalMux I__7853 (
            .O(N__32643),
            .I(N__32599));
    LocalMux I__7852 (
            .O(N__32634),
            .I(N__32599));
    InMux I__7851 (
            .O(N__32631),
            .I(N__32596));
    CascadeMux I__7850 (
            .O(N__32630),
            .I(N__32590));
    CascadeMux I__7849 (
            .O(N__32629),
            .I(N__32583));
    CascadeMux I__7848 (
            .O(N__32628),
            .I(N__32577));
    CascadeMux I__7847 (
            .O(N__32627),
            .I(N__32573));
    Span4Mux_v I__7846 (
            .O(N__32622),
            .I(N__32565));
    LocalMux I__7845 (
            .O(N__32619),
            .I(N__32565));
    InMux I__7844 (
            .O(N__32616),
            .I(N__32561));
    LocalMux I__7843 (
            .O(N__32613),
            .I(N__32554));
    Span4Mux_s3_v I__7842 (
            .O(N__32610),
            .I(N__32554));
    LocalMux I__7841 (
            .O(N__32607),
            .I(N__32554));
    LocalMux I__7840 (
            .O(N__32604),
            .I(N__32547));
    Span4Mux_v I__7839 (
            .O(N__32599),
            .I(N__32547));
    LocalMux I__7838 (
            .O(N__32596),
            .I(N__32547));
    CascadeMux I__7837 (
            .O(N__32595),
            .I(N__32540));
    CascadeMux I__7836 (
            .O(N__32594),
            .I(N__32537));
    CascadeMux I__7835 (
            .O(N__32593),
            .I(N__32534));
    InMux I__7834 (
            .O(N__32590),
            .I(N__32531));
    CascadeMux I__7833 (
            .O(N__32589),
            .I(N__32528));
    CascadeMux I__7832 (
            .O(N__32588),
            .I(N__32519));
    InMux I__7831 (
            .O(N__32587),
            .I(N__32513));
    InMux I__7830 (
            .O(N__32586),
            .I(N__32508));
    InMux I__7829 (
            .O(N__32583),
            .I(N__32508));
    CascadeMux I__7828 (
            .O(N__32582),
            .I(N__32499));
    InMux I__7827 (
            .O(N__32581),
            .I(N__32496));
    InMux I__7826 (
            .O(N__32580),
            .I(N__32493));
    InMux I__7825 (
            .O(N__32577),
            .I(N__32490));
    InMux I__7824 (
            .O(N__32576),
            .I(N__32487));
    InMux I__7823 (
            .O(N__32573),
            .I(N__32484));
    CascadeMux I__7822 (
            .O(N__32572),
            .I(N__32480));
    CascadeMux I__7821 (
            .O(N__32571),
            .I(N__32477));
    CascadeMux I__7820 (
            .O(N__32570),
            .I(N__32472));
    Span4Mux_h I__7819 (
            .O(N__32565),
            .I(N__32469));
    CascadeMux I__7818 (
            .O(N__32564),
            .I(N__32466));
    LocalMux I__7817 (
            .O(N__32561),
            .I(N__32461));
    Span4Mux_v I__7816 (
            .O(N__32554),
            .I(N__32458));
    Span4Mux_v I__7815 (
            .O(N__32547),
            .I(N__32455));
    CascadeMux I__7814 (
            .O(N__32546),
            .I(N__32451));
    CascadeMux I__7813 (
            .O(N__32545),
            .I(N__32448));
    CascadeMux I__7812 (
            .O(N__32544),
            .I(N__32440));
    InMux I__7811 (
            .O(N__32543),
            .I(N__32437));
    InMux I__7810 (
            .O(N__32540),
            .I(N__32434));
    InMux I__7809 (
            .O(N__32537),
            .I(N__32429));
    InMux I__7808 (
            .O(N__32534),
            .I(N__32429));
    LocalMux I__7807 (
            .O(N__32531),
            .I(N__32426));
    InMux I__7806 (
            .O(N__32528),
            .I(N__32423));
    InMux I__7805 (
            .O(N__32527),
            .I(N__32418));
    InMux I__7804 (
            .O(N__32526),
            .I(N__32418));
    InMux I__7803 (
            .O(N__32525),
            .I(N__32413));
    InMux I__7802 (
            .O(N__32524),
            .I(N__32413));
    InMux I__7801 (
            .O(N__32523),
            .I(N__32407));
    InMux I__7800 (
            .O(N__32522),
            .I(N__32407));
    InMux I__7799 (
            .O(N__32519),
            .I(N__32404));
    InMux I__7798 (
            .O(N__32518),
            .I(N__32401));
    InMux I__7797 (
            .O(N__32517),
            .I(N__32396));
    InMux I__7796 (
            .O(N__32516),
            .I(N__32396));
    LocalMux I__7795 (
            .O(N__32513),
            .I(N__32391));
    LocalMux I__7794 (
            .O(N__32508),
            .I(N__32391));
    CascadeMux I__7793 (
            .O(N__32507),
            .I(N__32388));
    CascadeMux I__7792 (
            .O(N__32506),
            .I(N__32385));
    InMux I__7791 (
            .O(N__32505),
            .I(N__32382));
    InMux I__7790 (
            .O(N__32504),
            .I(N__32373));
    InMux I__7789 (
            .O(N__32503),
            .I(N__32373));
    InMux I__7788 (
            .O(N__32502),
            .I(N__32373));
    InMux I__7787 (
            .O(N__32499),
            .I(N__32373));
    LocalMux I__7786 (
            .O(N__32496),
            .I(N__32366));
    LocalMux I__7785 (
            .O(N__32493),
            .I(N__32366));
    LocalMux I__7784 (
            .O(N__32490),
            .I(N__32366));
    LocalMux I__7783 (
            .O(N__32487),
            .I(N__32361));
    LocalMux I__7782 (
            .O(N__32484),
            .I(N__32361));
    InMux I__7781 (
            .O(N__32483),
            .I(N__32356));
    InMux I__7780 (
            .O(N__32480),
            .I(N__32356));
    InMux I__7779 (
            .O(N__32477),
            .I(N__32351));
    InMux I__7778 (
            .O(N__32476),
            .I(N__32351));
    InMux I__7777 (
            .O(N__32475),
            .I(N__32346));
    InMux I__7776 (
            .O(N__32472),
            .I(N__32346));
    Sp12to4 I__7775 (
            .O(N__32469),
            .I(N__32343));
    InMux I__7774 (
            .O(N__32466),
            .I(N__32340));
    InMux I__7773 (
            .O(N__32465),
            .I(N__32337));
    InMux I__7772 (
            .O(N__32464),
            .I(N__32334));
    Span4Mux_v I__7771 (
            .O(N__32461),
            .I(N__32329));
    Span4Mux_h I__7770 (
            .O(N__32458),
            .I(N__32329));
    Span4Mux_v I__7769 (
            .O(N__32455),
            .I(N__32326));
    InMux I__7768 (
            .O(N__32454),
            .I(N__32321));
    InMux I__7767 (
            .O(N__32451),
            .I(N__32321));
    InMux I__7766 (
            .O(N__32448),
            .I(N__32312));
    InMux I__7765 (
            .O(N__32447),
            .I(N__32309));
    InMux I__7764 (
            .O(N__32446),
            .I(N__32306));
    InMux I__7763 (
            .O(N__32445),
            .I(N__32297));
    InMux I__7762 (
            .O(N__32444),
            .I(N__32297));
    InMux I__7761 (
            .O(N__32443),
            .I(N__32297));
    InMux I__7760 (
            .O(N__32440),
            .I(N__32297));
    LocalMux I__7759 (
            .O(N__32437),
            .I(N__32286));
    LocalMux I__7758 (
            .O(N__32434),
            .I(N__32286));
    LocalMux I__7757 (
            .O(N__32429),
            .I(N__32286));
    Span4Mux_h I__7756 (
            .O(N__32426),
            .I(N__32286));
    LocalMux I__7755 (
            .O(N__32423),
            .I(N__32286));
    LocalMux I__7754 (
            .O(N__32418),
            .I(N__32281));
    LocalMux I__7753 (
            .O(N__32413),
            .I(N__32281));
    InMux I__7752 (
            .O(N__32412),
            .I(N__32278));
    LocalMux I__7751 (
            .O(N__32407),
            .I(N__32267));
    LocalMux I__7750 (
            .O(N__32404),
            .I(N__32267));
    LocalMux I__7749 (
            .O(N__32401),
            .I(N__32267));
    LocalMux I__7748 (
            .O(N__32396),
            .I(N__32267));
    Span4Mux_v I__7747 (
            .O(N__32391),
            .I(N__32267));
    InMux I__7746 (
            .O(N__32388),
            .I(N__32262));
    InMux I__7745 (
            .O(N__32385),
            .I(N__32262));
    LocalMux I__7744 (
            .O(N__32382),
            .I(N__32251));
    LocalMux I__7743 (
            .O(N__32373),
            .I(N__32251));
    Span4Mux_v I__7742 (
            .O(N__32366),
            .I(N__32251));
    Span4Mux_h I__7741 (
            .O(N__32361),
            .I(N__32251));
    LocalMux I__7740 (
            .O(N__32356),
            .I(N__32251));
    LocalMux I__7739 (
            .O(N__32351),
            .I(N__32232));
    LocalMux I__7738 (
            .O(N__32346),
            .I(N__32232));
    Span12Mux_s7_v I__7737 (
            .O(N__32343),
            .I(N__32232));
    LocalMux I__7736 (
            .O(N__32340),
            .I(N__32232));
    LocalMux I__7735 (
            .O(N__32337),
            .I(N__32232));
    LocalMux I__7734 (
            .O(N__32334),
            .I(N__32232));
    Sp12to4 I__7733 (
            .O(N__32329),
            .I(N__32232));
    Sp12to4 I__7732 (
            .O(N__32326),
            .I(N__32232));
    LocalMux I__7731 (
            .O(N__32321),
            .I(N__32232));
    InMux I__7730 (
            .O(N__32320),
            .I(N__32229));
    InMux I__7729 (
            .O(N__32319),
            .I(N__32226));
    InMux I__7728 (
            .O(N__32318),
            .I(N__32221));
    InMux I__7727 (
            .O(N__32317),
            .I(N__32221));
    InMux I__7726 (
            .O(N__32316),
            .I(N__32218));
    InMux I__7725 (
            .O(N__32315),
            .I(N__32215));
    LocalMux I__7724 (
            .O(N__32312),
            .I(N__32212));
    LocalMux I__7723 (
            .O(N__32309),
            .I(N__32203));
    LocalMux I__7722 (
            .O(N__32306),
            .I(N__32203));
    LocalMux I__7721 (
            .O(N__32297),
            .I(N__32203));
    Span4Mux_v I__7720 (
            .O(N__32286),
            .I(N__32203));
    Span4Mux_v I__7719 (
            .O(N__32281),
            .I(N__32192));
    LocalMux I__7718 (
            .O(N__32278),
            .I(N__32192));
    Span4Mux_v I__7717 (
            .O(N__32267),
            .I(N__32192));
    LocalMux I__7716 (
            .O(N__32262),
            .I(N__32192));
    Span4Mux_h I__7715 (
            .O(N__32251),
            .I(N__32192));
    Span12Mux_h I__7714 (
            .O(N__32232),
            .I(N__32189));
    LocalMux I__7713 (
            .O(N__32229),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__7712 (
            .O(N__32226),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__7711 (
            .O(N__32221),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__7710 (
            .O(N__32218),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__7709 (
            .O(N__32215),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv12 I__7708 (
            .O(N__32212),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__7707 (
            .O(N__32203),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__7706 (
            .O(N__32192),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv12 I__7705 (
            .O(N__32189),
            .I(\c0.byte_transmit_counter2_1 ));
    InMux I__7704 (
            .O(N__32170),
            .I(N__32167));
    LocalMux I__7703 (
            .O(N__32167),
            .I(N__32163));
    InMux I__7702 (
            .O(N__32166),
            .I(N__32158));
    Span4Mux_h I__7701 (
            .O(N__32163),
            .I(N__32155));
    InMux I__7700 (
            .O(N__32162),
            .I(N__32152));
    InMux I__7699 (
            .O(N__32161),
            .I(N__32149));
    LocalMux I__7698 (
            .O(N__32158),
            .I(\c0.data_in_field_110 ));
    Odrv4 I__7697 (
            .O(N__32155),
            .I(\c0.data_in_field_110 ));
    LocalMux I__7696 (
            .O(N__32152),
            .I(\c0.data_in_field_110 ));
    LocalMux I__7695 (
            .O(N__32149),
            .I(\c0.data_in_field_110 ));
    InMux I__7694 (
            .O(N__32140),
            .I(N__32137));
    LocalMux I__7693 (
            .O(N__32137),
            .I(\c0.n5384 ));
    CascadeMux I__7692 (
            .O(N__32134),
            .I(\c0.n5387_cascade_ ));
    InMux I__7691 (
            .O(N__32131),
            .I(N__32128));
    LocalMux I__7690 (
            .O(N__32128),
            .I(N__32125));
    Span4Mux_v I__7689 (
            .O(N__32125),
            .I(N__32119));
    InMux I__7688 (
            .O(N__32124),
            .I(N__32116));
    InMux I__7687 (
            .O(N__32123),
            .I(N__32112));
    InMux I__7686 (
            .O(N__32122),
            .I(N__32109));
    Span4Mux_h I__7685 (
            .O(N__32119),
            .I(N__32103));
    LocalMux I__7684 (
            .O(N__32116),
            .I(N__32103));
    InMux I__7683 (
            .O(N__32115),
            .I(N__32100));
    LocalMux I__7682 (
            .O(N__32112),
            .I(N__32092));
    LocalMux I__7681 (
            .O(N__32109),
            .I(N__32092));
    InMux I__7680 (
            .O(N__32108),
            .I(N__32089));
    Span4Mux_h I__7679 (
            .O(N__32103),
            .I(N__32086));
    LocalMux I__7678 (
            .O(N__32100),
            .I(N__32083));
    InMux I__7677 (
            .O(N__32099),
            .I(N__32080));
    InMux I__7676 (
            .O(N__32098),
            .I(N__32076));
    InMux I__7675 (
            .O(N__32097),
            .I(N__32073));
    Span4Mux_v I__7674 (
            .O(N__32092),
            .I(N__32070));
    LocalMux I__7673 (
            .O(N__32089),
            .I(N__32061));
    Span4Mux_h I__7672 (
            .O(N__32086),
            .I(N__32061));
    Span4Mux_s2_h I__7671 (
            .O(N__32083),
            .I(N__32061));
    LocalMux I__7670 (
            .O(N__32080),
            .I(N__32061));
    InMux I__7669 (
            .O(N__32079),
            .I(N__32058));
    LocalMux I__7668 (
            .O(N__32076),
            .I(\c0.byte_transmit_counter2_2 ));
    LocalMux I__7667 (
            .O(N__32073),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__7666 (
            .O(N__32070),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__7665 (
            .O(N__32061),
            .I(\c0.byte_transmit_counter2_2 ));
    LocalMux I__7664 (
            .O(N__32058),
            .I(\c0.byte_transmit_counter2_2 ));
    InMux I__7663 (
            .O(N__32047),
            .I(N__32044));
    LocalMux I__7662 (
            .O(N__32044),
            .I(N__32041));
    Odrv4 I__7661 (
            .O(N__32041),
            .I(\c0.n5378 ));
    InMux I__7660 (
            .O(N__32038),
            .I(N__32035));
    LocalMux I__7659 (
            .O(N__32035),
            .I(N__32032));
    Span4Mux_h I__7658 (
            .O(N__32032),
            .I(N__32029));
    Odrv4 I__7657 (
            .O(N__32029),
            .I(\c0.n5381 ));
    InMux I__7656 (
            .O(N__32026),
            .I(N__32023));
    LocalMux I__7655 (
            .O(N__32023),
            .I(N__32019));
    InMux I__7654 (
            .O(N__32022),
            .I(N__32016));
    Span4Mux_s2_h I__7653 (
            .O(N__32019),
            .I(N__32011));
    LocalMux I__7652 (
            .O(N__32016),
            .I(N__32011));
    Span4Mux_v I__7651 (
            .O(N__32011),
            .I(N__32007));
    InMux I__7650 (
            .O(N__32010),
            .I(N__32003));
    Span4Mux_h I__7649 (
            .O(N__32007),
            .I(N__32000));
    InMux I__7648 (
            .O(N__32006),
            .I(N__31996));
    LocalMux I__7647 (
            .O(N__32003),
            .I(N__31993));
    Span4Mux_h I__7646 (
            .O(N__32000),
            .I(N__31990));
    InMux I__7645 (
            .O(N__31999),
            .I(N__31987));
    LocalMux I__7644 (
            .O(N__31996),
            .I(\c0.data_in_field_136 ));
    Odrv4 I__7643 (
            .O(N__31993),
            .I(\c0.data_in_field_136 ));
    Odrv4 I__7642 (
            .O(N__31990),
            .I(\c0.data_in_field_136 ));
    LocalMux I__7641 (
            .O(N__31987),
            .I(\c0.data_in_field_136 ));
    CascadeMux I__7640 (
            .O(N__31978),
            .I(N__31975));
    InMux I__7639 (
            .O(N__31975),
            .I(N__31972));
    LocalMux I__7638 (
            .O(N__31972),
            .I(N__31969));
    Span4Mux_v I__7637 (
            .O(N__31969),
            .I(N__31964));
    InMux I__7636 (
            .O(N__31968),
            .I(N__31959));
    InMux I__7635 (
            .O(N__31967),
            .I(N__31959));
    Odrv4 I__7634 (
            .O(N__31964),
            .I(data_in_15_2));
    LocalMux I__7633 (
            .O(N__31959),
            .I(data_in_15_2));
    InMux I__7632 (
            .O(N__31954),
            .I(N__31950));
    InMux I__7631 (
            .O(N__31953),
            .I(N__31947));
    LocalMux I__7630 (
            .O(N__31950),
            .I(N__31943));
    LocalMux I__7629 (
            .O(N__31947),
            .I(N__31940));
    InMux I__7628 (
            .O(N__31946),
            .I(N__31937));
    Span4Mux_h I__7627 (
            .O(N__31943),
            .I(N__31933));
    Span4Mux_v I__7626 (
            .O(N__31940),
            .I(N__31926));
    LocalMux I__7625 (
            .O(N__31937),
            .I(N__31926));
    InMux I__7624 (
            .O(N__31936),
            .I(N__31923));
    Span4Mux_h I__7623 (
            .O(N__31933),
            .I(N__31920));
    CascadeMux I__7622 (
            .O(N__31932),
            .I(N__31917));
    InMux I__7621 (
            .O(N__31931),
            .I(N__31914));
    Span4Mux_h I__7620 (
            .O(N__31926),
            .I(N__31911));
    LocalMux I__7619 (
            .O(N__31923),
            .I(N__31906));
    Span4Mux_h I__7618 (
            .O(N__31920),
            .I(N__31906));
    InMux I__7617 (
            .O(N__31917),
            .I(N__31903));
    LocalMux I__7616 (
            .O(N__31914),
            .I(\c0.data_in_field_122 ));
    Odrv4 I__7615 (
            .O(N__31911),
            .I(\c0.data_in_field_122 ));
    Odrv4 I__7614 (
            .O(N__31906),
            .I(\c0.data_in_field_122 ));
    LocalMux I__7613 (
            .O(N__31903),
            .I(\c0.data_in_field_122 ));
    InMux I__7612 (
            .O(N__31894),
            .I(N__31891));
    LocalMux I__7611 (
            .O(N__31891),
            .I(N__31888));
    Span4Mux_h I__7610 (
            .O(N__31888),
            .I(N__31885));
    Span4Mux_v I__7609 (
            .O(N__31885),
            .I(N__31880));
    InMux I__7608 (
            .O(N__31884),
            .I(N__31875));
    InMux I__7607 (
            .O(N__31883),
            .I(N__31875));
    Odrv4 I__7606 (
            .O(N__31880),
            .I(data_in_14_3));
    LocalMux I__7605 (
            .O(N__31875),
            .I(data_in_14_3));
    CascadeMux I__7604 (
            .O(N__31870),
            .I(N__31867));
    InMux I__7603 (
            .O(N__31867),
            .I(N__31864));
    LocalMux I__7602 (
            .O(N__31864),
            .I(N__31861));
    Span4Mux_h I__7601 (
            .O(N__31861),
            .I(N__31858));
    Span4Mux_v I__7600 (
            .O(N__31858),
            .I(N__31855));
    Span4Mux_h I__7599 (
            .O(N__31855),
            .I(N__31850));
    InMux I__7598 (
            .O(N__31854),
            .I(N__31845));
    InMux I__7597 (
            .O(N__31853),
            .I(N__31845));
    Odrv4 I__7596 (
            .O(N__31850),
            .I(data_in_13_3));
    LocalMux I__7595 (
            .O(N__31845),
            .I(data_in_13_3));
    CascadeMux I__7594 (
            .O(N__31840),
            .I(N__31837));
    InMux I__7593 (
            .O(N__31837),
            .I(N__31834));
    LocalMux I__7592 (
            .O(N__31834),
            .I(N__31831));
    Span4Mux_h I__7591 (
            .O(N__31831),
            .I(N__31828));
    Span4Mux_h I__7590 (
            .O(N__31828),
            .I(N__31825));
    Span4Mux_h I__7589 (
            .O(N__31825),
            .I(N__31820));
    InMux I__7588 (
            .O(N__31824),
            .I(N__31815));
    InMux I__7587 (
            .O(N__31823),
            .I(N__31815));
    Odrv4 I__7586 (
            .O(N__31820),
            .I(data_in_12_3));
    LocalMux I__7585 (
            .O(N__31815),
            .I(data_in_12_3));
    InMux I__7584 (
            .O(N__31810),
            .I(N__31807));
    LocalMux I__7583 (
            .O(N__31807),
            .I(N__31803));
    CascadeMux I__7582 (
            .O(N__31806),
            .I(N__31800));
    Span4Mux_h I__7581 (
            .O(N__31803),
            .I(N__31796));
    InMux I__7580 (
            .O(N__31800),
            .I(N__31791));
    InMux I__7579 (
            .O(N__31799),
            .I(N__31791));
    Odrv4 I__7578 (
            .O(N__31796),
            .I(data_in_11_3));
    LocalMux I__7577 (
            .O(N__31791),
            .I(data_in_11_3));
    InMux I__7576 (
            .O(N__31786),
            .I(N__31782));
    InMux I__7575 (
            .O(N__31785),
            .I(N__31779));
    LocalMux I__7574 (
            .O(N__31782),
            .I(N__31776));
    LocalMux I__7573 (
            .O(N__31779),
            .I(N__31772));
    Span4Mux_h I__7572 (
            .O(N__31776),
            .I(N__31769));
    InMux I__7571 (
            .O(N__31775),
            .I(N__31764));
    Span4Mux_h I__7570 (
            .O(N__31772),
            .I(N__31759));
    Span4Mux_h I__7569 (
            .O(N__31769),
            .I(N__31759));
    InMux I__7568 (
            .O(N__31768),
            .I(N__31756));
    InMux I__7567 (
            .O(N__31767),
            .I(N__31753));
    LocalMux I__7566 (
            .O(N__31764),
            .I(\c0.data_in_field_91 ));
    Odrv4 I__7565 (
            .O(N__31759),
            .I(\c0.data_in_field_91 ));
    LocalMux I__7564 (
            .O(N__31756),
            .I(\c0.data_in_field_91 ));
    LocalMux I__7563 (
            .O(N__31753),
            .I(\c0.data_in_field_91 ));
    InMux I__7562 (
            .O(N__31744),
            .I(N__31741));
    LocalMux I__7561 (
            .O(N__31741),
            .I(N__31738));
    Span4Mux_v I__7560 (
            .O(N__31738),
            .I(N__31735));
    Span4Mux_h I__7559 (
            .O(N__31735),
            .I(N__31732));
    Span4Mux_h I__7558 (
            .O(N__31732),
            .I(N__31727));
    InMux I__7557 (
            .O(N__31731),
            .I(N__31724));
    InMux I__7556 (
            .O(N__31730),
            .I(N__31721));
    Odrv4 I__7555 (
            .O(N__31727),
            .I(data_in_0_3));
    LocalMux I__7554 (
            .O(N__31724),
            .I(data_in_0_3));
    LocalMux I__7553 (
            .O(N__31721),
            .I(data_in_0_3));
    InMux I__7552 (
            .O(N__31714),
            .I(N__31711));
    LocalMux I__7551 (
            .O(N__31711),
            .I(N__31706));
    InMux I__7550 (
            .O(N__31710),
            .I(N__31703));
    CascadeMux I__7549 (
            .O(N__31709),
            .I(N__31700));
    Span4Mux_h I__7548 (
            .O(N__31706),
            .I(N__31697));
    LocalMux I__7547 (
            .O(N__31703),
            .I(N__31694));
    InMux I__7546 (
            .O(N__31700),
            .I(N__31690));
    Span4Mux_h I__7545 (
            .O(N__31697),
            .I(N__31687));
    Span4Mux_h I__7544 (
            .O(N__31694),
            .I(N__31684));
    InMux I__7543 (
            .O(N__31693),
            .I(N__31681));
    LocalMux I__7542 (
            .O(N__31690),
            .I(\c0.data_in_field_3 ));
    Odrv4 I__7541 (
            .O(N__31687),
            .I(\c0.data_in_field_3 ));
    Odrv4 I__7540 (
            .O(N__31684),
            .I(\c0.data_in_field_3 ));
    LocalMux I__7539 (
            .O(N__31681),
            .I(\c0.data_in_field_3 ));
    InMux I__7538 (
            .O(N__31672),
            .I(N__31668));
    InMux I__7537 (
            .O(N__31671),
            .I(N__31665));
    LocalMux I__7536 (
            .O(N__31668),
            .I(N__31662));
    LocalMux I__7535 (
            .O(N__31665),
            .I(N__31659));
    Span4Mux_v I__7534 (
            .O(N__31662),
            .I(N__31656));
    Span4Mux_h I__7533 (
            .O(N__31659),
            .I(N__31653));
    Span4Mux_h I__7532 (
            .O(N__31656),
            .I(N__31647));
    Span4Mux_v I__7531 (
            .O(N__31653),
            .I(N__31647));
    InMux I__7530 (
            .O(N__31652),
            .I(N__31644));
    Odrv4 I__7529 (
            .O(N__31647),
            .I(data_in_11_2));
    LocalMux I__7528 (
            .O(N__31644),
            .I(data_in_11_2));
    CascadeMux I__7527 (
            .O(N__31639),
            .I(N__31636));
    InMux I__7526 (
            .O(N__31636),
            .I(N__31633));
    LocalMux I__7525 (
            .O(N__31633),
            .I(N__31630));
    Span4Mux_v I__7524 (
            .O(N__31630),
            .I(N__31627));
    Span4Mux_h I__7523 (
            .O(N__31627),
            .I(N__31624));
    Span4Mux_h I__7522 (
            .O(N__31624),
            .I(N__31619));
    InMux I__7521 (
            .O(N__31623),
            .I(N__31614));
    InMux I__7520 (
            .O(N__31622),
            .I(N__31614));
    Odrv4 I__7519 (
            .O(N__31619),
            .I(data_in_10_2));
    LocalMux I__7518 (
            .O(N__31614),
            .I(data_in_10_2));
    CascadeMux I__7517 (
            .O(N__31609),
            .I(N__31606));
    InMux I__7516 (
            .O(N__31606),
            .I(N__31603));
    LocalMux I__7515 (
            .O(N__31603),
            .I(N__31600));
    Span4Mux_v I__7514 (
            .O(N__31600),
            .I(N__31595));
    InMux I__7513 (
            .O(N__31599),
            .I(N__31590));
    InMux I__7512 (
            .O(N__31598),
            .I(N__31590));
    Odrv4 I__7511 (
            .O(N__31595),
            .I(data_in_5_4));
    LocalMux I__7510 (
            .O(N__31590),
            .I(data_in_5_4));
    InMux I__7509 (
            .O(N__31585),
            .I(N__31582));
    LocalMux I__7508 (
            .O(N__31582),
            .I(N__31579));
    Span4Mux_v I__7507 (
            .O(N__31579),
            .I(N__31576));
    Span4Mux_h I__7506 (
            .O(N__31576),
            .I(N__31571));
    InMux I__7505 (
            .O(N__31575),
            .I(N__31568));
    InMux I__7504 (
            .O(N__31574),
            .I(N__31565));
    Span4Mux_h I__7503 (
            .O(N__31571),
            .I(N__31560));
    LocalMux I__7502 (
            .O(N__31568),
            .I(N__31560));
    LocalMux I__7501 (
            .O(N__31565),
            .I(\c0.data_in_field_44 ));
    Odrv4 I__7500 (
            .O(N__31560),
            .I(\c0.data_in_field_44 ));
    InMux I__7499 (
            .O(N__31555),
            .I(N__31551));
    InMux I__7498 (
            .O(N__31554),
            .I(N__31548));
    LocalMux I__7497 (
            .O(N__31551),
            .I(N__31543));
    LocalMux I__7496 (
            .O(N__31548),
            .I(N__31543));
    Span4Mux_v I__7495 (
            .O(N__31543),
            .I(N__31539));
    InMux I__7494 (
            .O(N__31542),
            .I(N__31536));
    Span4Mux_h I__7493 (
            .O(N__31539),
            .I(N__31531));
    LocalMux I__7492 (
            .O(N__31536),
            .I(N__31531));
    Odrv4 I__7491 (
            .O(N__31531),
            .I(\c0.n1962 ));
    InMux I__7490 (
            .O(N__31528),
            .I(N__31525));
    LocalMux I__7489 (
            .O(N__31525),
            .I(N__31521));
    InMux I__7488 (
            .O(N__31524),
            .I(N__31518));
    Span4Mux_s3_v I__7487 (
            .O(N__31521),
            .I(N__31514));
    LocalMux I__7486 (
            .O(N__31518),
            .I(N__31510));
    InMux I__7485 (
            .O(N__31517),
            .I(N__31507));
    Span4Mux_h I__7484 (
            .O(N__31514),
            .I(N__31504));
    InMux I__7483 (
            .O(N__31513),
            .I(N__31501));
    Span4Mux_h I__7482 (
            .O(N__31510),
            .I(N__31496));
    LocalMux I__7481 (
            .O(N__31507),
            .I(N__31496));
    Odrv4 I__7480 (
            .O(N__31504),
            .I(data_in_3_0));
    LocalMux I__7479 (
            .O(N__31501),
            .I(data_in_3_0));
    Odrv4 I__7478 (
            .O(N__31496),
            .I(data_in_3_0));
    CascadeMux I__7477 (
            .O(N__31489),
            .I(N__31485));
    InMux I__7476 (
            .O(N__31488),
            .I(N__31482));
    InMux I__7475 (
            .O(N__31485),
            .I(N__31477));
    LocalMux I__7474 (
            .O(N__31482),
            .I(N__31474));
    InMux I__7473 (
            .O(N__31481),
            .I(N__31471));
    InMux I__7472 (
            .O(N__31480),
            .I(N__31468));
    LocalMux I__7471 (
            .O(N__31477),
            .I(\c0.data_in_field_24 ));
    Odrv4 I__7470 (
            .O(N__31474),
            .I(\c0.data_in_field_24 ));
    LocalMux I__7469 (
            .O(N__31471),
            .I(\c0.data_in_field_24 ));
    LocalMux I__7468 (
            .O(N__31468),
            .I(\c0.data_in_field_24 ));
    CascadeMux I__7467 (
            .O(N__31459),
            .I(N__31455));
    InMux I__7466 (
            .O(N__31458),
            .I(N__31452));
    InMux I__7465 (
            .O(N__31455),
            .I(N__31449));
    LocalMux I__7464 (
            .O(N__31452),
            .I(N__31446));
    LocalMux I__7463 (
            .O(N__31449),
            .I(N__31441));
    Span4Mux_h I__7462 (
            .O(N__31446),
            .I(N__31441));
    Span4Mux_h I__7461 (
            .O(N__31441),
            .I(N__31436));
    CascadeMux I__7460 (
            .O(N__31440),
            .I(N__31433));
    InMux I__7459 (
            .O(N__31439),
            .I(N__31430));
    Span4Mux_h I__7458 (
            .O(N__31436),
            .I(N__31427));
    InMux I__7457 (
            .O(N__31433),
            .I(N__31424));
    LocalMux I__7456 (
            .O(N__31430),
            .I(data_in_2_0));
    Odrv4 I__7455 (
            .O(N__31427),
            .I(data_in_2_0));
    LocalMux I__7454 (
            .O(N__31424),
            .I(data_in_2_0));
    InMux I__7453 (
            .O(N__31417),
            .I(N__31413));
    InMux I__7452 (
            .O(N__31416),
            .I(N__31410));
    LocalMux I__7451 (
            .O(N__31413),
            .I(N__31406));
    LocalMux I__7450 (
            .O(N__31410),
            .I(N__31403));
    CascadeMux I__7449 (
            .O(N__31409),
            .I(N__31399));
    Span4Mux_v I__7448 (
            .O(N__31406),
            .I(N__31394));
    Span4Mux_h I__7447 (
            .O(N__31403),
            .I(N__31394));
    InMux I__7446 (
            .O(N__31402),
            .I(N__31391));
    InMux I__7445 (
            .O(N__31399),
            .I(N__31388));
    Span4Mux_h I__7444 (
            .O(N__31394),
            .I(N__31385));
    LocalMux I__7443 (
            .O(N__31391),
            .I(data_in_1_0));
    LocalMux I__7442 (
            .O(N__31388),
            .I(data_in_1_0));
    Odrv4 I__7441 (
            .O(N__31385),
            .I(data_in_1_0));
    CascadeMux I__7440 (
            .O(N__31378),
            .I(N__31375));
    InMux I__7439 (
            .O(N__31375),
            .I(N__31372));
    LocalMux I__7438 (
            .O(N__31372),
            .I(N__31368));
    InMux I__7437 (
            .O(N__31371),
            .I(N__31365));
    Span4Mux_h I__7436 (
            .O(N__31368),
            .I(N__31361));
    LocalMux I__7435 (
            .O(N__31365),
            .I(N__31358));
    InMux I__7434 (
            .O(N__31364),
            .I(N__31355));
    Odrv4 I__7433 (
            .O(N__31361),
            .I(data_in_15_3));
    Odrv4 I__7432 (
            .O(N__31358),
            .I(data_in_15_3));
    LocalMux I__7431 (
            .O(N__31355),
            .I(data_in_15_3));
    InMux I__7430 (
            .O(N__31348),
            .I(N__31345));
    LocalMux I__7429 (
            .O(N__31345),
            .I(N__31341));
    InMux I__7428 (
            .O(N__31344),
            .I(N__31338));
    Span4Mux_h I__7427 (
            .O(N__31341),
            .I(N__31335));
    LocalMux I__7426 (
            .O(N__31338),
            .I(N__31332));
    Span4Mux_v I__7425 (
            .O(N__31335),
            .I(N__31327));
    Span4Mux_h I__7424 (
            .O(N__31332),
            .I(N__31324));
    InMux I__7423 (
            .O(N__31331),
            .I(N__31321));
    InMux I__7422 (
            .O(N__31330),
            .I(N__31318));
    Span4Mux_h I__7421 (
            .O(N__31327),
            .I(N__31313));
    Span4Mux_h I__7420 (
            .O(N__31324),
            .I(N__31313));
    LocalMux I__7419 (
            .O(N__31321),
            .I(\c0.data_in_field_123 ));
    LocalMux I__7418 (
            .O(N__31318),
            .I(\c0.data_in_field_123 ));
    Odrv4 I__7417 (
            .O(N__31313),
            .I(\c0.data_in_field_123 ));
    InMux I__7416 (
            .O(N__31306),
            .I(N__31300));
    InMux I__7415 (
            .O(N__31305),
            .I(N__31300));
    LocalMux I__7414 (
            .O(N__31300),
            .I(N__31296));
    InMux I__7413 (
            .O(N__31299),
            .I(N__31293));
    Odrv4 I__7412 (
            .O(N__31296),
            .I(data_in_12_6));
    LocalMux I__7411 (
            .O(N__31293),
            .I(data_in_12_6));
    CascadeMux I__7410 (
            .O(N__31288),
            .I(N__31285));
    InMux I__7409 (
            .O(N__31285),
            .I(N__31281));
    InMux I__7408 (
            .O(N__31284),
            .I(N__31278));
    LocalMux I__7407 (
            .O(N__31281),
            .I(N__31275));
    LocalMux I__7406 (
            .O(N__31278),
            .I(N__31271));
    Span4Mux_h I__7405 (
            .O(N__31275),
            .I(N__31268));
    InMux I__7404 (
            .O(N__31274),
            .I(N__31265));
    Span12Mux_v I__7403 (
            .O(N__31271),
            .I(N__31262));
    Span4Mux_h I__7402 (
            .O(N__31268),
            .I(N__31259));
    LocalMux I__7401 (
            .O(N__31265),
            .I(data_in_11_6));
    Odrv12 I__7400 (
            .O(N__31262),
            .I(data_in_11_6));
    Odrv4 I__7399 (
            .O(N__31259),
            .I(data_in_11_6));
    CascadeMux I__7398 (
            .O(N__31252),
            .I(N__31248));
    CascadeMux I__7397 (
            .O(N__31251),
            .I(N__31244));
    InMux I__7396 (
            .O(N__31248),
            .I(N__31241));
    InMux I__7395 (
            .O(N__31247),
            .I(N__31238));
    InMux I__7394 (
            .O(N__31244),
            .I(N__31234));
    LocalMux I__7393 (
            .O(N__31241),
            .I(N__31229));
    LocalMux I__7392 (
            .O(N__31238),
            .I(N__31229));
    CascadeMux I__7391 (
            .O(N__31237),
            .I(N__31226));
    LocalMux I__7390 (
            .O(N__31234),
            .I(N__31223));
    Span4Mux_v I__7389 (
            .O(N__31229),
            .I(N__31220));
    InMux I__7388 (
            .O(N__31226),
            .I(N__31217));
    Sp12to4 I__7387 (
            .O(N__31223),
            .I(N__31214));
    Span4Mux_h I__7386 (
            .O(N__31220),
            .I(N__31211));
    LocalMux I__7385 (
            .O(N__31217),
            .I(data_in_18_2));
    Odrv12 I__7384 (
            .O(N__31214),
            .I(data_in_18_2));
    Odrv4 I__7383 (
            .O(N__31211),
            .I(data_in_18_2));
    InMux I__7382 (
            .O(N__31204),
            .I(N__31200));
    InMux I__7381 (
            .O(N__31203),
            .I(N__31197));
    LocalMux I__7380 (
            .O(N__31200),
            .I(N__31194));
    LocalMux I__7379 (
            .O(N__31197),
            .I(N__31191));
    Span4Mux_v I__7378 (
            .O(N__31194),
            .I(N__31185));
    Span4Mux_h I__7377 (
            .O(N__31191),
            .I(N__31185));
    InMux I__7376 (
            .O(N__31190),
            .I(N__31181));
    Span4Mux_h I__7375 (
            .O(N__31185),
            .I(N__31178));
    InMux I__7374 (
            .O(N__31184),
            .I(N__31175));
    LocalMux I__7373 (
            .O(N__31181),
            .I(\c0.data_in_field_74 ));
    Odrv4 I__7372 (
            .O(N__31178),
            .I(\c0.data_in_field_74 ));
    LocalMux I__7371 (
            .O(N__31175),
            .I(\c0.data_in_field_74 ));
    CascadeMux I__7370 (
            .O(N__31168),
            .I(N__31165));
    InMux I__7369 (
            .O(N__31165),
            .I(N__31162));
    LocalMux I__7368 (
            .O(N__31162),
            .I(N__31159));
    Span4Mux_s2_v I__7367 (
            .O(N__31159),
            .I(N__31156));
    Span4Mux_v I__7366 (
            .O(N__31156),
            .I(N__31151));
    InMux I__7365 (
            .O(N__31155),
            .I(N__31146));
    InMux I__7364 (
            .O(N__31154),
            .I(N__31146));
    Odrv4 I__7363 (
            .O(N__31151),
            .I(data_in_15_1));
    LocalMux I__7362 (
            .O(N__31146),
            .I(data_in_15_1));
    CascadeMux I__7361 (
            .O(N__31141),
            .I(N__31138));
    InMux I__7360 (
            .O(N__31138),
            .I(N__31134));
    InMux I__7359 (
            .O(N__31137),
            .I(N__31131));
    LocalMux I__7358 (
            .O(N__31134),
            .I(N__31127));
    LocalMux I__7357 (
            .O(N__31131),
            .I(N__31124));
    InMux I__7356 (
            .O(N__31130),
            .I(N__31121));
    Odrv4 I__7355 (
            .O(N__31127),
            .I(data_in_14_4));
    Odrv4 I__7354 (
            .O(N__31124),
            .I(data_in_14_4));
    LocalMux I__7353 (
            .O(N__31121),
            .I(data_in_14_4));
    InMux I__7352 (
            .O(N__31114),
            .I(N__31111));
    LocalMux I__7351 (
            .O(N__31111),
            .I(N__31108));
    Span12Mux_h I__7350 (
            .O(N__31108),
            .I(N__31103));
    InMux I__7349 (
            .O(N__31107),
            .I(N__31098));
    InMux I__7348 (
            .O(N__31106),
            .I(N__31098));
    Odrv12 I__7347 (
            .O(N__31103),
            .I(\c0.data_in_field_116 ));
    LocalMux I__7346 (
            .O(N__31098),
            .I(\c0.data_in_field_116 ));
    InMux I__7345 (
            .O(N__31093),
            .I(N__31090));
    LocalMux I__7344 (
            .O(N__31090),
            .I(N__31087));
    Span4Mux_v I__7343 (
            .O(N__31087),
            .I(N__31084));
    Span4Mux_h I__7342 (
            .O(N__31084),
            .I(N__31080));
    InMux I__7341 (
            .O(N__31083),
            .I(N__31077));
    Odrv4 I__7340 (
            .O(N__31080),
            .I(\c0.n1815 ));
    LocalMux I__7339 (
            .O(N__31077),
            .I(\c0.n1815 ));
    CascadeMux I__7338 (
            .O(N__31072),
            .I(\c0.n1815_cascade_ ));
    InMux I__7337 (
            .O(N__31069),
            .I(N__31065));
    InMux I__7336 (
            .O(N__31068),
            .I(N__31062));
    LocalMux I__7335 (
            .O(N__31065),
            .I(N__31059));
    LocalMux I__7334 (
            .O(N__31062),
            .I(N__31056));
    Span4Mux_h I__7333 (
            .O(N__31059),
            .I(N__31053));
    Span4Mux_h I__7332 (
            .O(N__31056),
            .I(N__31050));
    Span4Mux_v I__7331 (
            .O(N__31053),
            .I(N__31045));
    Span4Mux_h I__7330 (
            .O(N__31050),
            .I(N__31042));
    InMux I__7329 (
            .O(N__31049),
            .I(N__31037));
    InMux I__7328 (
            .O(N__31048),
            .I(N__31037));
    Odrv4 I__7327 (
            .O(N__31045),
            .I(\c0.data_in_field_52 ));
    Odrv4 I__7326 (
            .O(N__31042),
            .I(\c0.data_in_field_52 ));
    LocalMux I__7325 (
            .O(N__31037),
            .I(\c0.data_in_field_52 ));
    CascadeMux I__7324 (
            .O(N__31030),
            .I(N__31027));
    InMux I__7323 (
            .O(N__31027),
            .I(N__31024));
    LocalMux I__7322 (
            .O(N__31024),
            .I(N__31021));
    Span4Mux_h I__7321 (
            .O(N__31021),
            .I(N__31018));
    Span4Mux_h I__7320 (
            .O(N__31018),
            .I(N__31015));
    Odrv4 I__7319 (
            .O(N__31015),
            .I(\c0.n27 ));
    CascadeMux I__7318 (
            .O(N__31012),
            .I(N__31009));
    InMux I__7317 (
            .O(N__31009),
            .I(N__31006));
    LocalMux I__7316 (
            .O(N__31006),
            .I(N__31003));
    Span4Mux_h I__7315 (
            .O(N__31003),
            .I(N__31000));
    Span4Mux_h I__7314 (
            .O(N__31000),
            .I(N__30996));
    InMux I__7313 (
            .O(N__30999),
            .I(N__30993));
    Span4Mux_v I__7312 (
            .O(N__30996),
            .I(N__30987));
    LocalMux I__7311 (
            .O(N__30993),
            .I(N__30987));
    InMux I__7310 (
            .O(N__30992),
            .I(N__30984));
    Odrv4 I__7309 (
            .O(N__30987),
            .I(data_in_14_1));
    LocalMux I__7308 (
            .O(N__30984),
            .I(data_in_14_1));
    InMux I__7307 (
            .O(N__30979),
            .I(N__30976));
    LocalMux I__7306 (
            .O(N__30976),
            .I(N__30972));
    InMux I__7305 (
            .O(N__30975),
            .I(N__30969));
    Span4Mux_v I__7304 (
            .O(N__30972),
            .I(N__30966));
    LocalMux I__7303 (
            .O(N__30969),
            .I(N__30963));
    Span4Mux_h I__7302 (
            .O(N__30966),
            .I(N__30960));
    Span4Mux_v I__7301 (
            .O(N__30963),
            .I(N__30957));
    Span4Mux_h I__7300 (
            .O(N__30960),
            .I(N__30953));
    Span4Mux_h I__7299 (
            .O(N__30957),
            .I(N__30950));
    InMux I__7298 (
            .O(N__30956),
            .I(N__30947));
    Odrv4 I__7297 (
            .O(N__30953),
            .I(data_in_13_1));
    Odrv4 I__7296 (
            .O(N__30950),
            .I(data_in_13_1));
    LocalMux I__7295 (
            .O(N__30947),
            .I(data_in_13_1));
    CascadeMux I__7294 (
            .O(N__30940),
            .I(N__30937));
    InMux I__7293 (
            .O(N__30937),
            .I(N__30934));
    LocalMux I__7292 (
            .O(N__30934),
            .I(N__30931));
    Span4Mux_h I__7291 (
            .O(N__30931),
            .I(N__30926));
    InMux I__7290 (
            .O(N__30930),
            .I(N__30921));
    InMux I__7289 (
            .O(N__30929),
            .I(N__30921));
    Odrv4 I__7288 (
            .O(N__30926),
            .I(data_in_7_0));
    LocalMux I__7287 (
            .O(N__30921),
            .I(data_in_7_0));
    InMux I__7286 (
            .O(N__30916),
            .I(N__30912));
    InMux I__7285 (
            .O(N__30915),
            .I(N__30909));
    LocalMux I__7284 (
            .O(N__30912),
            .I(N__30904));
    LocalMux I__7283 (
            .O(N__30909),
            .I(N__30901));
    InMux I__7282 (
            .O(N__30908),
            .I(N__30896));
    InMux I__7281 (
            .O(N__30907),
            .I(N__30896));
    Span4Mux_h I__7280 (
            .O(N__30904),
            .I(N__30893));
    Odrv4 I__7279 (
            .O(N__30901),
            .I(\c0.data_in_field_56 ));
    LocalMux I__7278 (
            .O(N__30896),
            .I(\c0.data_in_field_56 ));
    Odrv4 I__7277 (
            .O(N__30893),
            .I(\c0.data_in_field_56 ));
    InMux I__7276 (
            .O(N__30886),
            .I(N__30882));
    InMux I__7275 (
            .O(N__30885),
            .I(N__30879));
    LocalMux I__7274 (
            .O(N__30882),
            .I(N__30876));
    LocalMux I__7273 (
            .O(N__30879),
            .I(N__30873));
    Span4Mux_v I__7272 (
            .O(N__30876),
            .I(N__30869));
    Span4Mux_v I__7271 (
            .O(N__30873),
            .I(N__30866));
    InMux I__7270 (
            .O(N__30872),
            .I(N__30862));
    Span4Mux_h I__7269 (
            .O(N__30869),
            .I(N__30857));
    Span4Mux_h I__7268 (
            .O(N__30866),
            .I(N__30857));
    InMux I__7267 (
            .O(N__30865),
            .I(N__30854));
    LocalMux I__7266 (
            .O(N__30862),
            .I(N__30851));
    Span4Mux_h I__7265 (
            .O(N__30857),
            .I(N__30844));
    LocalMux I__7264 (
            .O(N__30854),
            .I(N__30844));
    Span4Mux_v I__7263 (
            .O(N__30851),
            .I(N__30841));
    InMux I__7262 (
            .O(N__30850),
            .I(N__30836));
    InMux I__7261 (
            .O(N__30849),
            .I(N__30836));
    Span4Mux_v I__7260 (
            .O(N__30844),
            .I(N__30833));
    Odrv4 I__7259 (
            .O(N__30841),
            .I(\c0.data_in_field_129 ));
    LocalMux I__7258 (
            .O(N__30836),
            .I(\c0.data_in_field_129 ));
    Odrv4 I__7257 (
            .O(N__30833),
            .I(\c0.data_in_field_129 ));
    InMux I__7256 (
            .O(N__30826),
            .I(N__30823));
    LocalMux I__7255 (
            .O(N__30823),
            .I(N__30820));
    Span4Mux_h I__7254 (
            .O(N__30820),
            .I(N__30817));
    Odrv4 I__7253 (
            .O(N__30817),
            .I(\c0.n15_adj_1923 ));
    InMux I__7252 (
            .O(N__30814),
            .I(N__30811));
    LocalMux I__7251 (
            .O(N__30811),
            .I(N__30808));
    Span4Mux_v I__7250 (
            .O(N__30808),
            .I(N__30803));
    InMux I__7249 (
            .O(N__30807),
            .I(N__30798));
    InMux I__7248 (
            .O(N__30806),
            .I(N__30798));
    Odrv4 I__7247 (
            .O(N__30803),
            .I(data_in_6_2));
    LocalMux I__7246 (
            .O(N__30798),
            .I(data_in_6_2));
    InMux I__7245 (
            .O(N__30793),
            .I(N__30789));
    CascadeMux I__7244 (
            .O(N__30792),
            .I(N__30784));
    LocalMux I__7243 (
            .O(N__30789),
            .I(N__30781));
    CascadeMux I__7242 (
            .O(N__30788),
            .I(N__30778));
    CascadeMux I__7241 (
            .O(N__30787),
            .I(N__30775));
    InMux I__7240 (
            .O(N__30784),
            .I(N__30772));
    Span4Mux_h I__7239 (
            .O(N__30781),
            .I(N__30769));
    InMux I__7238 (
            .O(N__30778),
            .I(N__30764));
    InMux I__7237 (
            .O(N__30775),
            .I(N__30764));
    LocalMux I__7236 (
            .O(N__30772),
            .I(\c0.data_in_field_50 ));
    Odrv4 I__7235 (
            .O(N__30769),
            .I(\c0.data_in_field_50 ));
    LocalMux I__7234 (
            .O(N__30764),
            .I(\c0.data_in_field_50 ));
    InMux I__7233 (
            .O(N__30757),
            .I(N__30754));
    LocalMux I__7232 (
            .O(N__30754),
            .I(N__30750));
    InMux I__7231 (
            .O(N__30753),
            .I(N__30746));
    Span4Mux_h I__7230 (
            .O(N__30750),
            .I(N__30743));
    InMux I__7229 (
            .O(N__30749),
            .I(N__30739));
    LocalMux I__7228 (
            .O(N__30746),
            .I(N__30736));
    Span4Mux_h I__7227 (
            .O(N__30743),
            .I(N__30733));
    InMux I__7226 (
            .O(N__30742),
            .I(N__30730));
    LocalMux I__7225 (
            .O(N__30739),
            .I(\c0.data_in_field_8 ));
    Odrv4 I__7224 (
            .O(N__30736),
            .I(\c0.data_in_field_8 ));
    Odrv4 I__7223 (
            .O(N__30733),
            .I(\c0.data_in_field_8 ));
    LocalMux I__7222 (
            .O(N__30730),
            .I(\c0.data_in_field_8 ));
    InMux I__7221 (
            .O(N__30721),
            .I(N__30718));
    LocalMux I__7220 (
            .O(N__30718),
            .I(N__30715));
    Span4Mux_h I__7219 (
            .O(N__30715),
            .I(N__30710));
    InMux I__7218 (
            .O(N__30714),
            .I(N__30705));
    InMux I__7217 (
            .O(N__30713),
            .I(N__30705));
    Odrv4 I__7216 (
            .O(N__30710),
            .I(data_in_8_2));
    LocalMux I__7215 (
            .O(N__30705),
            .I(data_in_8_2));
    CascadeMux I__7214 (
            .O(N__30700),
            .I(N__30696));
    InMux I__7213 (
            .O(N__30699),
            .I(N__30693));
    InMux I__7212 (
            .O(N__30696),
            .I(N__30690));
    LocalMux I__7211 (
            .O(N__30693),
            .I(N__30687));
    LocalMux I__7210 (
            .O(N__30690),
            .I(N__30681));
    Span4Mux_h I__7209 (
            .O(N__30687),
            .I(N__30681));
    InMux I__7208 (
            .O(N__30686),
            .I(N__30678));
    Odrv4 I__7207 (
            .O(N__30681),
            .I(data_in_14_2));
    LocalMux I__7206 (
            .O(N__30678),
            .I(data_in_14_2));
    InMux I__7205 (
            .O(N__30673),
            .I(N__30669));
    CascadeMux I__7204 (
            .O(N__30672),
            .I(N__30665));
    LocalMux I__7203 (
            .O(N__30669),
            .I(N__30661));
    InMux I__7202 (
            .O(N__30668),
            .I(N__30658));
    InMux I__7201 (
            .O(N__30665),
            .I(N__30655));
    InMux I__7200 (
            .O(N__30664),
            .I(N__30652));
    Span4Mux_h I__7199 (
            .O(N__30661),
            .I(N__30649));
    LocalMux I__7198 (
            .O(N__30658),
            .I(N__30645));
    LocalMux I__7197 (
            .O(N__30655),
            .I(N__30642));
    LocalMux I__7196 (
            .O(N__30652),
            .I(N__30639));
    Span4Mux_h I__7195 (
            .O(N__30649),
            .I(N__30636));
    InMux I__7194 (
            .O(N__30648),
            .I(N__30633));
    Span12Mux_v I__7193 (
            .O(N__30645),
            .I(N__30626));
    Span12Mux_s6_v I__7192 (
            .O(N__30642),
            .I(N__30626));
    Span12Mux_s8_h I__7191 (
            .O(N__30639),
            .I(N__30626));
    Span4Mux_h I__7190 (
            .O(N__30636),
            .I(N__30623));
    LocalMux I__7189 (
            .O(N__30633),
            .I(\c0.data_in_field_114 ));
    Odrv12 I__7188 (
            .O(N__30626),
            .I(\c0.data_in_field_114 ));
    Odrv4 I__7187 (
            .O(N__30623),
            .I(\c0.data_in_field_114 ));
    CascadeMux I__7186 (
            .O(N__30616),
            .I(N__30612));
    InMux I__7185 (
            .O(N__30615),
            .I(N__30609));
    InMux I__7184 (
            .O(N__30612),
            .I(N__30606));
    LocalMux I__7183 (
            .O(N__30609),
            .I(N__30603));
    LocalMux I__7182 (
            .O(N__30606),
            .I(N__30600));
    Span4Mux_h I__7181 (
            .O(N__30603),
            .I(N__30597));
    Span4Mux_v I__7180 (
            .O(N__30600),
            .I(N__30593));
    Span4Mux_h I__7179 (
            .O(N__30597),
            .I(N__30590));
    InMux I__7178 (
            .O(N__30596),
            .I(N__30587));
    Odrv4 I__7177 (
            .O(N__30593),
            .I(data_in_4_2));
    Odrv4 I__7176 (
            .O(N__30590),
            .I(data_in_4_2));
    LocalMux I__7175 (
            .O(N__30587),
            .I(data_in_4_2));
    InMux I__7174 (
            .O(N__30580),
            .I(N__30576));
    InMux I__7173 (
            .O(N__30579),
            .I(N__30573));
    LocalMux I__7172 (
            .O(N__30576),
            .I(N__30567));
    LocalMux I__7171 (
            .O(N__30573),
            .I(N__30564));
    InMux I__7170 (
            .O(N__30572),
            .I(N__30561));
    InMux I__7169 (
            .O(N__30571),
            .I(N__30556));
    InMux I__7168 (
            .O(N__30570),
            .I(N__30556));
    Odrv4 I__7167 (
            .O(N__30567),
            .I(\c0.data_in_field_66 ));
    Odrv4 I__7166 (
            .O(N__30564),
            .I(\c0.data_in_field_66 ));
    LocalMux I__7165 (
            .O(N__30561),
            .I(\c0.data_in_field_66 ));
    LocalMux I__7164 (
            .O(N__30556),
            .I(\c0.data_in_field_66 ));
    CascadeMux I__7163 (
            .O(N__30547),
            .I(N__30543));
    InMux I__7162 (
            .O(N__30546),
            .I(N__30540));
    InMux I__7161 (
            .O(N__30543),
            .I(N__30537));
    LocalMux I__7160 (
            .O(N__30540),
            .I(N__30534));
    LocalMux I__7159 (
            .O(N__30537),
            .I(N__30531));
    Span4Mux_h I__7158 (
            .O(N__30534),
            .I(N__30526));
    Span4Mux_h I__7157 (
            .O(N__30531),
            .I(N__30523));
    InMux I__7156 (
            .O(N__30530),
            .I(N__30518));
    InMux I__7155 (
            .O(N__30529),
            .I(N__30518));
    Odrv4 I__7154 (
            .O(N__30526),
            .I(\c0.data_in_field_84 ));
    Odrv4 I__7153 (
            .O(N__30523),
            .I(\c0.data_in_field_84 ));
    LocalMux I__7152 (
            .O(N__30518),
            .I(\c0.data_in_field_84 ));
    InMux I__7151 (
            .O(N__30511),
            .I(N__30508));
    LocalMux I__7150 (
            .O(N__30508),
            .I(N__30505));
    Span4Mux_v I__7149 (
            .O(N__30505),
            .I(N__30501));
    InMux I__7148 (
            .O(N__30504),
            .I(N__30498));
    Span4Mux_h I__7147 (
            .O(N__30501),
            .I(N__30494));
    LocalMux I__7146 (
            .O(N__30498),
            .I(N__30491));
    InMux I__7145 (
            .O(N__30497),
            .I(N__30488));
    Odrv4 I__7144 (
            .O(N__30494),
            .I(\c0.n1969 ));
    Odrv4 I__7143 (
            .O(N__30491),
            .I(\c0.n1969 ));
    LocalMux I__7142 (
            .O(N__30488),
            .I(\c0.n1969 ));
    InMux I__7141 (
            .O(N__30481),
            .I(N__30478));
    LocalMux I__7140 (
            .O(N__30478),
            .I(N__30475));
    Span4Mux_h I__7139 (
            .O(N__30475),
            .I(N__30472));
    Odrv4 I__7138 (
            .O(N__30472),
            .I(\c0.n25 ));
    InMux I__7137 (
            .O(N__30469),
            .I(N__30463));
    InMux I__7136 (
            .O(N__30468),
            .I(N__30463));
    LocalMux I__7135 (
            .O(N__30463),
            .I(N__30459));
    InMux I__7134 (
            .O(N__30462),
            .I(N__30456));
    Odrv4 I__7133 (
            .O(N__30459),
            .I(data_in_5_2));
    LocalMux I__7132 (
            .O(N__30456),
            .I(data_in_5_2));
    InMux I__7131 (
            .O(N__30451),
            .I(N__30445));
    InMux I__7130 (
            .O(N__30450),
            .I(N__30442));
    CascadeMux I__7129 (
            .O(N__30449),
            .I(N__30439));
    InMux I__7128 (
            .O(N__30448),
            .I(N__30436));
    LocalMux I__7127 (
            .O(N__30445),
            .I(N__30433));
    LocalMux I__7126 (
            .O(N__30442),
            .I(N__30430));
    InMux I__7125 (
            .O(N__30439),
            .I(N__30427));
    LocalMux I__7124 (
            .O(N__30436),
            .I(N__30424));
    Span4Mux_h I__7123 (
            .O(N__30433),
            .I(N__30421));
    Span4Mux_v I__7122 (
            .O(N__30430),
            .I(N__30418));
    LocalMux I__7121 (
            .O(N__30427),
            .I(\c0.data_in_field_42 ));
    Odrv4 I__7120 (
            .O(N__30424),
            .I(\c0.data_in_field_42 ));
    Odrv4 I__7119 (
            .O(N__30421),
            .I(\c0.data_in_field_42 ));
    Odrv4 I__7118 (
            .O(N__30418),
            .I(\c0.data_in_field_42 ));
    CascadeMux I__7117 (
            .O(N__30409),
            .I(N__30406));
    InMux I__7116 (
            .O(N__30406),
            .I(N__30401));
    InMux I__7115 (
            .O(N__30405),
            .I(N__30398));
    InMux I__7114 (
            .O(N__30404),
            .I(N__30395));
    LocalMux I__7113 (
            .O(N__30401),
            .I(N__30392));
    LocalMux I__7112 (
            .O(N__30398),
            .I(N__30389));
    LocalMux I__7111 (
            .O(N__30395),
            .I(N__30386));
    Span4Mux_v I__7110 (
            .O(N__30392),
            .I(N__30383));
    Span4Mux_v I__7109 (
            .O(N__30389),
            .I(N__30378));
    Span4Mux_v I__7108 (
            .O(N__30386),
            .I(N__30375));
    Span4Mux_h I__7107 (
            .O(N__30383),
            .I(N__30372));
    InMux I__7106 (
            .O(N__30382),
            .I(N__30367));
    InMux I__7105 (
            .O(N__30381),
            .I(N__30367));
    Odrv4 I__7104 (
            .O(N__30378),
            .I(\c0.data_in_field_107 ));
    Odrv4 I__7103 (
            .O(N__30375),
            .I(\c0.data_in_field_107 ));
    Odrv4 I__7102 (
            .O(N__30372),
            .I(\c0.data_in_field_107 ));
    LocalMux I__7101 (
            .O(N__30367),
            .I(\c0.data_in_field_107 ));
    InMux I__7100 (
            .O(N__30358),
            .I(N__30355));
    LocalMux I__7099 (
            .O(N__30355),
            .I(N__30350));
    InMux I__7098 (
            .O(N__30354),
            .I(N__30347));
    CascadeMux I__7097 (
            .O(N__30353),
            .I(N__30344));
    Sp12to4 I__7096 (
            .O(N__30350),
            .I(N__30341));
    LocalMux I__7095 (
            .O(N__30347),
            .I(N__30338));
    InMux I__7094 (
            .O(N__30344),
            .I(N__30334));
    Span12Mux_v I__7093 (
            .O(N__30341),
            .I(N__30331));
    Span4Mux_h I__7092 (
            .O(N__30338),
            .I(N__30328));
    InMux I__7091 (
            .O(N__30337),
            .I(N__30325));
    LocalMux I__7090 (
            .O(N__30334),
            .I(\c0.data_in_field_15 ));
    Odrv12 I__7089 (
            .O(N__30331),
            .I(\c0.data_in_field_15 ));
    Odrv4 I__7088 (
            .O(N__30328),
            .I(\c0.data_in_field_15 ));
    LocalMux I__7087 (
            .O(N__30325),
            .I(\c0.data_in_field_15 ));
    InMux I__7086 (
            .O(N__30316),
            .I(N__30313));
    LocalMux I__7085 (
            .O(N__30313),
            .I(N__30310));
    Span4Mux_h I__7084 (
            .O(N__30310),
            .I(N__30307));
    Span4Mux_h I__7083 (
            .O(N__30307),
            .I(N__30304));
    Odrv4 I__7082 (
            .O(N__30304),
            .I(\c0.n20_adj_1916 ));
    CascadeMux I__7081 (
            .O(N__30301),
            .I(N__30298));
    InMux I__7080 (
            .O(N__30298),
            .I(N__30294));
    InMux I__7079 (
            .O(N__30297),
            .I(N__30291));
    LocalMux I__7078 (
            .O(N__30294),
            .I(N__30288));
    LocalMux I__7077 (
            .O(N__30291),
            .I(N__30285));
    Span4Mux_v I__7076 (
            .O(N__30288),
            .I(N__30279));
    Span4Mux_v I__7075 (
            .O(N__30285),
            .I(N__30279));
    InMux I__7074 (
            .O(N__30284),
            .I(N__30276));
    Odrv4 I__7073 (
            .O(N__30279),
            .I(data_in_8_1));
    LocalMux I__7072 (
            .O(N__30276),
            .I(data_in_8_1));
    InMux I__7071 (
            .O(N__30271),
            .I(N__30268));
    LocalMux I__7070 (
            .O(N__30268),
            .I(N__30264));
    CascadeMux I__7069 (
            .O(N__30267),
            .I(N__30261));
    Sp12to4 I__7068 (
            .O(N__30264),
            .I(N__30254));
    InMux I__7067 (
            .O(N__30261),
            .I(N__30251));
    InMux I__7066 (
            .O(N__30260),
            .I(N__30248));
    InMux I__7065 (
            .O(N__30259),
            .I(N__30243));
    InMux I__7064 (
            .O(N__30258),
            .I(N__30243));
    InMux I__7063 (
            .O(N__30257),
            .I(N__30240));
    Span12Mux_s6_v I__7062 (
            .O(N__30254),
            .I(N__30233));
    LocalMux I__7061 (
            .O(N__30251),
            .I(N__30233));
    LocalMux I__7060 (
            .O(N__30248),
            .I(N__30233));
    LocalMux I__7059 (
            .O(N__30243),
            .I(N__30230));
    LocalMux I__7058 (
            .O(N__30240),
            .I(\c0.data_in_field_65 ));
    Odrv12 I__7057 (
            .O(N__30233),
            .I(\c0.data_in_field_65 ));
    Odrv4 I__7056 (
            .O(N__30230),
            .I(\c0.data_in_field_65 ));
    CascadeMux I__7055 (
            .O(N__30223),
            .I(N__30220));
    InMux I__7054 (
            .O(N__30220),
            .I(N__30217));
    LocalMux I__7053 (
            .O(N__30217),
            .I(N__30213));
    InMux I__7052 (
            .O(N__30216),
            .I(N__30210));
    Span4Mux_v I__7051 (
            .O(N__30213),
            .I(N__30207));
    LocalMux I__7050 (
            .O(N__30210),
            .I(N__30204));
    Span4Mux_v I__7049 (
            .O(N__30207),
            .I(N__30200));
    Span12Mux_h I__7048 (
            .O(N__30204),
            .I(N__30197));
    InMux I__7047 (
            .O(N__30203),
            .I(N__30194));
    Odrv4 I__7046 (
            .O(N__30200),
            .I(data_in_16_1));
    Odrv12 I__7045 (
            .O(N__30197),
            .I(data_in_16_1));
    LocalMux I__7044 (
            .O(N__30194),
            .I(data_in_16_1));
    InMux I__7043 (
            .O(N__30187),
            .I(N__30182));
    InMux I__7042 (
            .O(N__30186),
            .I(N__30178));
    InMux I__7041 (
            .O(N__30185),
            .I(N__30175));
    LocalMux I__7040 (
            .O(N__30182),
            .I(N__30172));
    InMux I__7039 (
            .O(N__30181),
            .I(N__30169));
    LocalMux I__7038 (
            .O(N__30178),
            .I(N__30164));
    LocalMux I__7037 (
            .O(N__30175),
            .I(N__30164));
    Odrv4 I__7036 (
            .O(N__30172),
            .I(data_in_2_1));
    LocalMux I__7035 (
            .O(N__30169),
            .I(data_in_2_1));
    Odrv12 I__7034 (
            .O(N__30164),
            .I(data_in_2_1));
    InMux I__7033 (
            .O(N__30157),
            .I(N__30154));
    LocalMux I__7032 (
            .O(N__30154),
            .I(N__30150));
    InMux I__7031 (
            .O(N__30153),
            .I(N__30145));
    Span4Mux_h I__7030 (
            .O(N__30150),
            .I(N__30142));
    InMux I__7029 (
            .O(N__30149),
            .I(N__30137));
    InMux I__7028 (
            .O(N__30148),
            .I(N__30137));
    LocalMux I__7027 (
            .O(N__30145),
            .I(N__30134));
    Odrv4 I__7026 (
            .O(N__30142),
            .I(data_in_1_1));
    LocalMux I__7025 (
            .O(N__30137),
            .I(data_in_1_1));
    Odrv12 I__7024 (
            .O(N__30134),
            .I(data_in_1_1));
    CascadeMux I__7023 (
            .O(N__30127),
            .I(N__30124));
    InMux I__7022 (
            .O(N__30124),
            .I(N__30120));
    CascadeMux I__7021 (
            .O(N__30123),
            .I(N__30116));
    LocalMux I__7020 (
            .O(N__30120),
            .I(N__30113));
    CascadeMux I__7019 (
            .O(N__30119),
            .I(N__30110));
    InMux I__7018 (
            .O(N__30116),
            .I(N__30107));
    Span4Mux_h I__7017 (
            .O(N__30113),
            .I(N__30104));
    InMux I__7016 (
            .O(N__30110),
            .I(N__30101));
    LocalMux I__7015 (
            .O(N__30107),
            .I(N__30097));
    Sp12to4 I__7014 (
            .O(N__30104),
            .I(N__30092));
    LocalMux I__7013 (
            .O(N__30101),
            .I(N__30092));
    InMux I__7012 (
            .O(N__30100),
            .I(N__30089));
    Odrv4 I__7011 (
            .O(N__30097),
            .I(\c0.data_in_field_48 ));
    Odrv12 I__7010 (
            .O(N__30092),
            .I(\c0.data_in_field_48 ));
    LocalMux I__7009 (
            .O(N__30089),
            .I(\c0.data_in_field_48 ));
    CascadeMux I__7008 (
            .O(N__30082),
            .I(N__30079));
    InMux I__7007 (
            .O(N__30079),
            .I(N__30076));
    LocalMux I__7006 (
            .O(N__30076),
            .I(\c0.n5701 ));
    InMux I__7005 (
            .O(N__30073),
            .I(N__30069));
    InMux I__7004 (
            .O(N__30072),
            .I(N__30066));
    LocalMux I__7003 (
            .O(N__30069),
            .I(N__30063));
    LocalMux I__7002 (
            .O(N__30066),
            .I(N__30060));
    Sp12to4 I__7001 (
            .O(N__30063),
            .I(N__30057));
    Span4Mux_h I__7000 (
            .O(N__30060),
            .I(N__30054));
    Span12Mux_s7_v I__6999 (
            .O(N__30057),
            .I(N__30050));
    Span4Mux_v I__6998 (
            .O(N__30054),
            .I(N__30047));
    InMux I__6997 (
            .O(N__30053),
            .I(N__30044));
    Odrv12 I__6996 (
            .O(N__30050),
            .I(data_in_4_4));
    Odrv4 I__6995 (
            .O(N__30047),
            .I(data_in_4_4));
    LocalMux I__6994 (
            .O(N__30044),
            .I(data_in_4_4));
    CascadeMux I__6993 (
            .O(N__30037),
            .I(N__30034));
    InMux I__6992 (
            .O(N__30034),
            .I(N__30031));
    LocalMux I__6991 (
            .O(N__30031),
            .I(N__30027));
    InMux I__6990 (
            .O(N__30030),
            .I(N__30024));
    Span4Mux_v I__6989 (
            .O(N__30027),
            .I(N__30021));
    LocalMux I__6988 (
            .O(N__30024),
            .I(N__30018));
    Span4Mux_h I__6987 (
            .O(N__30021),
            .I(N__30013));
    Span4Mux_h I__6986 (
            .O(N__30018),
            .I(N__30013));
    Span4Mux_v I__6985 (
            .O(N__30013),
            .I(N__30009));
    InMux I__6984 (
            .O(N__30012),
            .I(N__30006));
    Odrv4 I__6983 (
            .O(N__30009),
            .I(data_in_6_4));
    LocalMux I__6982 (
            .O(N__30006),
            .I(data_in_6_4));
    InMux I__6981 (
            .O(N__30001),
            .I(N__29998));
    LocalMux I__6980 (
            .O(N__29998),
            .I(N__29995));
    Span4Mux_h I__6979 (
            .O(N__29995),
            .I(N__29990));
    InMux I__6978 (
            .O(N__29994),
            .I(N__29987));
    InMux I__6977 (
            .O(N__29993),
            .I(N__29984));
    Odrv4 I__6976 (
            .O(N__29990),
            .I(data_in_7_2));
    LocalMux I__6975 (
            .O(N__29987),
            .I(data_in_7_2));
    LocalMux I__6974 (
            .O(N__29984),
            .I(data_in_7_2));
    InMux I__6973 (
            .O(N__29977),
            .I(N__29974));
    LocalMux I__6972 (
            .O(N__29974),
            .I(N__29971));
    Span4Mux_v I__6971 (
            .O(N__29971),
            .I(N__29967));
    InMux I__6970 (
            .O(N__29970),
            .I(N__29964));
    Sp12to4 I__6969 (
            .O(N__29967),
            .I(N__29961));
    LocalMux I__6968 (
            .O(N__29964),
            .I(N__29958));
    Span12Mux_s10_h I__6967 (
            .O(N__29961),
            .I(N__29954));
    Span4Mux_h I__6966 (
            .O(N__29958),
            .I(N__29951));
    InMux I__6965 (
            .O(N__29957),
            .I(N__29948));
    Odrv12 I__6964 (
            .O(N__29954),
            .I(data_in_10_6));
    Odrv4 I__6963 (
            .O(N__29951),
            .I(data_in_10_6));
    LocalMux I__6962 (
            .O(N__29948),
            .I(data_in_10_6));
    CascadeMux I__6961 (
            .O(N__29941),
            .I(N__29938));
    InMux I__6960 (
            .O(N__29938),
            .I(N__29935));
    LocalMux I__6959 (
            .O(N__29935),
            .I(N__29932));
    Span4Mux_h I__6958 (
            .O(N__29932),
            .I(N__29929));
    Span4Mux_h I__6957 (
            .O(N__29929),
            .I(N__29924));
    InMux I__6956 (
            .O(N__29928),
            .I(N__29921));
    InMux I__6955 (
            .O(N__29927),
            .I(N__29918));
    Odrv4 I__6954 (
            .O(N__29924),
            .I(data_in_9_6));
    LocalMux I__6953 (
            .O(N__29921),
            .I(data_in_9_6));
    LocalMux I__6952 (
            .O(N__29918),
            .I(data_in_9_6));
    InMux I__6951 (
            .O(N__29911),
            .I(N__29907));
    InMux I__6950 (
            .O(N__29910),
            .I(N__29903));
    LocalMux I__6949 (
            .O(N__29907),
            .I(N__29900));
    InMux I__6948 (
            .O(N__29906),
            .I(N__29897));
    LocalMux I__6947 (
            .O(N__29903),
            .I(data_in_10_0));
    Odrv12 I__6946 (
            .O(N__29900),
            .I(data_in_10_0));
    LocalMux I__6945 (
            .O(N__29897),
            .I(data_in_10_0));
    InMux I__6944 (
            .O(N__29890),
            .I(N__29886));
    InMux I__6943 (
            .O(N__29889),
            .I(N__29882));
    LocalMux I__6942 (
            .O(N__29886),
            .I(N__29879));
    InMux I__6941 (
            .O(N__29885),
            .I(N__29876));
    LocalMux I__6940 (
            .O(N__29882),
            .I(N__29870));
    Span4Mux_v I__6939 (
            .O(N__29879),
            .I(N__29870));
    LocalMux I__6938 (
            .O(N__29876),
            .I(N__29867));
    CascadeMux I__6937 (
            .O(N__29875),
            .I(N__29864));
    Span4Mux_h I__6936 (
            .O(N__29870),
            .I(N__29861));
    Span4Mux_h I__6935 (
            .O(N__29867),
            .I(N__29858));
    InMux I__6934 (
            .O(N__29864),
            .I(N__29854));
    Span4Mux_h I__6933 (
            .O(N__29861),
            .I(N__29849));
    Span4Mux_h I__6932 (
            .O(N__29858),
            .I(N__29849));
    InMux I__6931 (
            .O(N__29857),
            .I(N__29846));
    LocalMux I__6930 (
            .O(N__29854),
            .I(\c0.data_in_field_80 ));
    Odrv4 I__6929 (
            .O(N__29849),
            .I(\c0.data_in_field_80 ));
    LocalMux I__6928 (
            .O(N__29846),
            .I(\c0.data_in_field_80 ));
    InMux I__6927 (
            .O(N__29839),
            .I(N__29834));
    InMux I__6926 (
            .O(N__29838),
            .I(N__29829));
    InMux I__6925 (
            .O(N__29837),
            .I(N__29829));
    LocalMux I__6924 (
            .O(N__29834),
            .I(data_in_13_6));
    LocalMux I__6923 (
            .O(N__29829),
            .I(data_in_13_6));
    InMux I__6922 (
            .O(N__29824),
            .I(N__29821));
    LocalMux I__6921 (
            .O(N__29821),
            .I(n5332));
    CascadeMux I__6920 (
            .O(N__29818),
            .I(n5331_cascade_));
    IoInMux I__6919 (
            .O(N__29815),
            .I(N__29812));
    LocalMux I__6918 (
            .O(N__29812),
            .I(N__29809));
    IoSpan4Mux I__6917 (
            .O(N__29809),
            .I(N__29806));
    IoSpan4Mux I__6916 (
            .O(N__29806),
            .I(N__29803));
    Odrv4 I__6915 (
            .O(N__29803),
            .I(LED_c));
    InMux I__6914 (
            .O(N__29800),
            .I(N__29796));
    InMux I__6913 (
            .O(N__29799),
            .I(N__29791));
    LocalMux I__6912 (
            .O(N__29796),
            .I(N__29787));
    CascadeMux I__6911 (
            .O(N__29795),
            .I(N__29783));
    InMux I__6910 (
            .O(N__29794),
            .I(N__29780));
    LocalMux I__6909 (
            .O(N__29791),
            .I(N__29777));
    InMux I__6908 (
            .O(N__29790),
            .I(N__29774));
    Span4Mux_v I__6907 (
            .O(N__29787),
            .I(N__29771));
    InMux I__6906 (
            .O(N__29786),
            .I(N__29768));
    InMux I__6905 (
            .O(N__29783),
            .I(N__29765));
    LocalMux I__6904 (
            .O(N__29780),
            .I(N__29762));
    Span4Mux_h I__6903 (
            .O(N__29777),
            .I(N__29757));
    LocalMux I__6902 (
            .O(N__29774),
            .I(N__29757));
    Span4Mux_h I__6901 (
            .O(N__29771),
            .I(N__29752));
    LocalMux I__6900 (
            .O(N__29768),
            .I(N__29752));
    LocalMux I__6899 (
            .O(N__29765),
            .I(\c0.data_in_field_97 ));
    Odrv4 I__6898 (
            .O(N__29762),
            .I(\c0.data_in_field_97 ));
    Odrv4 I__6897 (
            .O(N__29757),
            .I(\c0.data_in_field_97 ));
    Odrv4 I__6896 (
            .O(N__29752),
            .I(\c0.data_in_field_97 ));
    CascadeMux I__6895 (
            .O(N__29743),
            .I(N__29740));
    InMux I__6894 (
            .O(N__29740),
            .I(N__29736));
    InMux I__6893 (
            .O(N__29739),
            .I(N__29733));
    LocalMux I__6892 (
            .O(N__29736),
            .I(N__29730));
    LocalMux I__6891 (
            .O(N__29733),
            .I(N__29727));
    Span4Mux_v I__6890 (
            .O(N__29730),
            .I(N__29724));
    Span12Mux_v I__6889 (
            .O(N__29727),
            .I(N__29721));
    Span4Mux_h I__6888 (
            .O(N__29724),
            .I(N__29718));
    Odrv12 I__6887 (
            .O(N__29721),
            .I(\c0.n1972 ));
    Odrv4 I__6886 (
            .O(N__29718),
            .I(\c0.n1972 ));
    CascadeMux I__6885 (
            .O(N__29713),
            .I(N__29710));
    InMux I__6884 (
            .O(N__29710),
            .I(N__29707));
    LocalMux I__6883 (
            .O(N__29707),
            .I(N__29704));
    Span4Mux_v I__6882 (
            .O(N__29704),
            .I(N__29699));
    InMux I__6881 (
            .O(N__29703),
            .I(N__29696));
    InMux I__6880 (
            .O(N__29702),
            .I(N__29693));
    Odrv4 I__6879 (
            .O(N__29699),
            .I(data_in_9_4));
    LocalMux I__6878 (
            .O(N__29696),
            .I(data_in_9_4));
    LocalMux I__6877 (
            .O(N__29693),
            .I(data_in_9_4));
    InMux I__6876 (
            .O(N__29686),
            .I(N__29683));
    LocalMux I__6875 (
            .O(N__29683),
            .I(N__29680));
    Span4Mux_v I__6874 (
            .O(N__29680),
            .I(N__29677));
    Span4Mux_h I__6873 (
            .O(N__29677),
            .I(N__29671));
    InMux I__6872 (
            .O(N__29676),
            .I(N__29666));
    InMux I__6871 (
            .O(N__29675),
            .I(N__29666));
    InMux I__6870 (
            .O(N__29674),
            .I(N__29663));
    Odrv4 I__6869 (
            .O(N__29671),
            .I(\c0.data_in_field_76 ));
    LocalMux I__6868 (
            .O(N__29666),
            .I(\c0.data_in_field_76 ));
    LocalMux I__6867 (
            .O(N__29663),
            .I(\c0.data_in_field_76 ));
    CascadeMux I__6866 (
            .O(N__29656),
            .I(N__29652));
    InMux I__6865 (
            .O(N__29655),
            .I(N__29649));
    InMux I__6864 (
            .O(N__29652),
            .I(N__29646));
    LocalMux I__6863 (
            .O(N__29649),
            .I(N__29640));
    LocalMux I__6862 (
            .O(N__29646),
            .I(N__29640));
    InMux I__6861 (
            .O(N__29645),
            .I(N__29637));
    Span4Mux_h I__6860 (
            .O(N__29640),
            .I(N__29634));
    LocalMux I__6859 (
            .O(N__29637),
            .I(data_in_0_1));
    Odrv4 I__6858 (
            .O(N__29634),
            .I(data_in_0_1));
    CascadeMux I__6857 (
            .O(N__29629),
            .I(N__29626));
    InMux I__6856 (
            .O(N__29626),
            .I(N__29621));
    InMux I__6855 (
            .O(N__29625),
            .I(N__29618));
    InMux I__6854 (
            .O(N__29624),
            .I(N__29615));
    LocalMux I__6853 (
            .O(N__29621),
            .I(data_in_5_5));
    LocalMux I__6852 (
            .O(N__29618),
            .I(data_in_5_5));
    LocalMux I__6851 (
            .O(N__29615),
            .I(data_in_5_5));
    InMux I__6850 (
            .O(N__29608),
            .I(N__29604));
    InMux I__6849 (
            .O(N__29607),
            .I(N__29601));
    LocalMux I__6848 (
            .O(N__29604),
            .I(N__29598));
    LocalMux I__6847 (
            .O(N__29601),
            .I(N__29594));
    Span4Mux_h I__6846 (
            .O(N__29598),
            .I(N__29591));
    InMux I__6845 (
            .O(N__29597),
            .I(N__29587));
    Span4Mux_h I__6844 (
            .O(N__29594),
            .I(N__29584));
    Span4Mux_h I__6843 (
            .O(N__29591),
            .I(N__29581));
    InMux I__6842 (
            .O(N__29590),
            .I(N__29578));
    LocalMux I__6841 (
            .O(N__29587),
            .I(\c0.data_in_field_45 ));
    Odrv4 I__6840 (
            .O(N__29584),
            .I(\c0.data_in_field_45 ));
    Odrv4 I__6839 (
            .O(N__29581),
            .I(\c0.data_in_field_45 ));
    LocalMux I__6838 (
            .O(N__29578),
            .I(\c0.data_in_field_45 ));
    CascadeMux I__6837 (
            .O(N__29569),
            .I(N__29566));
    InMux I__6836 (
            .O(N__29566),
            .I(N__29563));
    LocalMux I__6835 (
            .O(N__29563),
            .I(N__29559));
    InMux I__6834 (
            .O(N__29562),
            .I(N__29556));
    Span4Mux_v I__6833 (
            .O(N__29559),
            .I(N__29551));
    LocalMux I__6832 (
            .O(N__29556),
            .I(N__29551));
    Span4Mux_v I__6831 (
            .O(N__29551),
            .I(N__29547));
    InMux I__6830 (
            .O(N__29550),
            .I(N__29544));
    Odrv4 I__6829 (
            .O(N__29547),
            .I(data_in_9_0));
    LocalMux I__6828 (
            .O(N__29544),
            .I(data_in_9_0));
    InMux I__6827 (
            .O(N__29539),
            .I(N__29536));
    LocalMux I__6826 (
            .O(N__29536),
            .I(N__29531));
    InMux I__6825 (
            .O(N__29535),
            .I(N__29528));
    InMux I__6824 (
            .O(N__29534),
            .I(N__29524));
    Span4Mux_v I__6823 (
            .O(N__29531),
            .I(N__29519));
    LocalMux I__6822 (
            .O(N__29528),
            .I(N__29519));
    InMux I__6821 (
            .O(N__29527),
            .I(N__29516));
    LocalMux I__6820 (
            .O(N__29524),
            .I(N__29512));
    Span4Mux_h I__6819 (
            .O(N__29519),
            .I(N__29509));
    LocalMux I__6818 (
            .O(N__29516),
            .I(N__29506));
    InMux I__6817 (
            .O(N__29515),
            .I(N__29503));
    Span12Mux_s9_h I__6816 (
            .O(N__29512),
            .I(N__29500));
    Span4Mux_h I__6815 (
            .O(N__29509),
            .I(N__29495));
    Span4Mux_h I__6814 (
            .O(N__29506),
            .I(N__29495));
    LocalMux I__6813 (
            .O(N__29503),
            .I(\c0.data_in_field_128 ));
    Odrv12 I__6812 (
            .O(N__29500),
            .I(\c0.data_in_field_128 ));
    Odrv4 I__6811 (
            .O(N__29495),
            .I(\c0.data_in_field_128 ));
    CascadeMux I__6810 (
            .O(N__29488),
            .I(N__29485));
    InMux I__6809 (
            .O(N__29485),
            .I(N__29480));
    InMux I__6808 (
            .O(N__29484),
            .I(N__29475));
    InMux I__6807 (
            .O(N__29483),
            .I(N__29475));
    LocalMux I__6806 (
            .O(N__29480),
            .I(N__29472));
    LocalMux I__6805 (
            .O(N__29475),
            .I(\c0.data_in_field_16 ));
    Odrv4 I__6804 (
            .O(N__29472),
            .I(\c0.data_in_field_16 ));
    CascadeMux I__6803 (
            .O(N__29467),
            .I(N__29464));
    InMux I__6802 (
            .O(N__29464),
            .I(N__29461));
    LocalMux I__6801 (
            .O(N__29461),
            .I(N__29458));
    Span4Mux_h I__6800 (
            .O(N__29458),
            .I(N__29452));
    InMux I__6799 (
            .O(N__29457),
            .I(N__29447));
    InMux I__6798 (
            .O(N__29456),
            .I(N__29447));
    InMux I__6797 (
            .O(N__29455),
            .I(N__29444));
    Odrv4 I__6796 (
            .O(N__29452),
            .I(\c0.data_in_field_72 ));
    LocalMux I__6795 (
            .O(N__29447),
            .I(\c0.data_in_field_72 ));
    LocalMux I__6794 (
            .O(N__29444),
            .I(\c0.data_in_field_72 ));
    InMux I__6793 (
            .O(N__29437),
            .I(N__29433));
    InMux I__6792 (
            .O(N__29436),
            .I(N__29430));
    LocalMux I__6791 (
            .O(N__29433),
            .I(\c0.n5188 ));
    LocalMux I__6790 (
            .O(N__29430),
            .I(\c0.n5188 ));
    CascadeMux I__6789 (
            .O(N__29425),
            .I(\c0.n5138_cascade_ ));
    InMux I__6788 (
            .O(N__29422),
            .I(N__29419));
    LocalMux I__6787 (
            .O(N__29419),
            .I(N__29416));
    Odrv12 I__6786 (
            .O(N__29416),
            .I(\c0.n15_adj_1968 ));
    InMux I__6785 (
            .O(N__29413),
            .I(N__29409));
    InMux I__6784 (
            .O(N__29412),
            .I(N__29406));
    LocalMux I__6783 (
            .O(N__29409),
            .I(N__29403));
    LocalMux I__6782 (
            .O(N__29406),
            .I(N__29400));
    Span4Mux_h I__6781 (
            .O(N__29403),
            .I(N__29393));
    Span4Mux_h I__6780 (
            .O(N__29400),
            .I(N__29393));
    CascadeMux I__6779 (
            .O(N__29399),
            .I(N__29390));
    InMux I__6778 (
            .O(N__29398),
            .I(N__29387));
    Span4Mux_v I__6777 (
            .O(N__29393),
            .I(N__29384));
    InMux I__6776 (
            .O(N__29390),
            .I(N__29381));
    LocalMux I__6775 (
            .O(N__29387),
            .I(data_in_3_2));
    Odrv4 I__6774 (
            .O(N__29384),
            .I(data_in_3_2));
    LocalMux I__6773 (
            .O(N__29381),
            .I(data_in_3_2));
    InMux I__6772 (
            .O(N__29374),
            .I(N__29371));
    LocalMux I__6771 (
            .O(N__29371),
            .I(N__29368));
    Span4Mux_h I__6770 (
            .O(N__29368),
            .I(N__29362));
    InMux I__6769 (
            .O(N__29367),
            .I(N__29356));
    InMux I__6768 (
            .O(N__29366),
            .I(N__29356));
    InMux I__6767 (
            .O(N__29365),
            .I(N__29353));
    Span4Mux_v I__6766 (
            .O(N__29362),
            .I(N__29350));
    InMux I__6765 (
            .O(N__29361),
            .I(N__29347));
    LocalMux I__6764 (
            .O(N__29356),
            .I(N__29344));
    LocalMux I__6763 (
            .O(N__29353),
            .I(\c0.data_in_field_26 ));
    Odrv4 I__6762 (
            .O(N__29350),
            .I(\c0.data_in_field_26 ));
    LocalMux I__6761 (
            .O(N__29347),
            .I(\c0.data_in_field_26 ));
    Odrv12 I__6760 (
            .O(N__29344),
            .I(\c0.data_in_field_26 ));
    InMux I__6759 (
            .O(N__29335),
            .I(N__29331));
    InMux I__6758 (
            .O(N__29334),
            .I(N__29328));
    LocalMux I__6757 (
            .O(N__29331),
            .I(N__29325));
    LocalMux I__6756 (
            .O(N__29328),
            .I(N__29321));
    Span4Mux_s3_v I__6755 (
            .O(N__29325),
            .I(N__29318));
    InMux I__6754 (
            .O(N__29324),
            .I(N__29315));
    Span12Mux_h I__6753 (
            .O(N__29321),
            .I(N__29312));
    Span4Mux_h I__6752 (
            .O(N__29318),
            .I(N__29309));
    LocalMux I__6751 (
            .O(N__29315),
            .I(data_in_4_1));
    Odrv12 I__6750 (
            .O(N__29312),
            .I(data_in_4_1));
    Odrv4 I__6749 (
            .O(N__29309),
            .I(data_in_4_1));
    InMux I__6748 (
            .O(N__29302),
            .I(N__29299));
    LocalMux I__6747 (
            .O(N__29299),
            .I(N__29295));
    CascadeMux I__6746 (
            .O(N__29298),
            .I(N__29291));
    Span4Mux_v I__6745 (
            .O(N__29295),
            .I(N__29288));
    InMux I__6744 (
            .O(N__29294),
            .I(N__29285));
    InMux I__6743 (
            .O(N__29291),
            .I(N__29281));
    Span4Mux_h I__6742 (
            .O(N__29288),
            .I(N__29276));
    LocalMux I__6741 (
            .O(N__29285),
            .I(N__29276));
    CascadeMux I__6740 (
            .O(N__29284),
            .I(N__29273));
    LocalMux I__6739 (
            .O(N__29281),
            .I(N__29270));
    Span4Mux_h I__6738 (
            .O(N__29276),
            .I(N__29267));
    InMux I__6737 (
            .O(N__29273),
            .I(N__29264));
    Odrv4 I__6736 (
            .O(N__29270),
            .I(\c0.data_in_field_33 ));
    Odrv4 I__6735 (
            .O(N__29267),
            .I(\c0.data_in_field_33 ));
    LocalMux I__6734 (
            .O(N__29264),
            .I(\c0.data_in_field_33 ));
    CascadeMux I__6733 (
            .O(N__29257),
            .I(N__29254));
    InMux I__6732 (
            .O(N__29254),
            .I(N__29251));
    LocalMux I__6731 (
            .O(N__29251),
            .I(N__29247));
    InMux I__6730 (
            .O(N__29250),
            .I(N__29243));
    Span4Mux_h I__6729 (
            .O(N__29247),
            .I(N__29240));
    InMux I__6728 (
            .O(N__29246),
            .I(N__29236));
    LocalMux I__6727 (
            .O(N__29243),
            .I(N__29233));
    Span4Mux_h I__6726 (
            .O(N__29240),
            .I(N__29230));
    InMux I__6725 (
            .O(N__29239),
            .I(N__29227));
    LocalMux I__6724 (
            .O(N__29236),
            .I(data_in_2_2));
    Odrv4 I__6723 (
            .O(N__29233),
            .I(data_in_2_2));
    Odrv4 I__6722 (
            .O(N__29230),
            .I(data_in_2_2));
    LocalMux I__6721 (
            .O(N__29227),
            .I(data_in_2_2));
    CascadeMux I__6720 (
            .O(N__29218),
            .I(N__29214));
    InMux I__6719 (
            .O(N__29217),
            .I(N__29211));
    InMux I__6718 (
            .O(N__29214),
            .I(N__29208));
    LocalMux I__6717 (
            .O(N__29211),
            .I(N__29205));
    LocalMux I__6716 (
            .O(N__29208),
            .I(N__29202));
    Span4Mux_h I__6715 (
            .O(N__29205),
            .I(N__29199));
    Span4Mux_h I__6714 (
            .O(N__29202),
            .I(N__29196));
    Span4Mux_v I__6713 (
            .O(N__29199),
            .I(N__29191));
    Span4Mux_h I__6712 (
            .O(N__29196),
            .I(N__29188));
    InMux I__6711 (
            .O(N__29195),
            .I(N__29183));
    InMux I__6710 (
            .O(N__29194),
            .I(N__29183));
    Odrv4 I__6709 (
            .O(N__29191),
            .I(\c0.data_in_field_18 ));
    Odrv4 I__6708 (
            .O(N__29188),
            .I(\c0.data_in_field_18 ));
    LocalMux I__6707 (
            .O(N__29183),
            .I(\c0.data_in_field_18 ));
    InMux I__6706 (
            .O(N__29176),
            .I(N__29173));
    LocalMux I__6705 (
            .O(N__29173),
            .I(\c0.n6 ));
    InMux I__6704 (
            .O(N__29170),
            .I(N__29166));
    InMux I__6703 (
            .O(N__29169),
            .I(N__29163));
    LocalMux I__6702 (
            .O(N__29166),
            .I(N__29160));
    LocalMux I__6701 (
            .O(N__29163),
            .I(N__29157));
    Span4Mux_v I__6700 (
            .O(N__29160),
            .I(N__29152));
    Span4Mux_v I__6699 (
            .O(N__29157),
            .I(N__29152));
    Sp12to4 I__6698 (
            .O(N__29152),
            .I(N__29148));
    InMux I__6697 (
            .O(N__29151),
            .I(N__29145));
    Odrv12 I__6696 (
            .O(N__29148),
            .I(data_in_4_0));
    LocalMux I__6695 (
            .O(N__29145),
            .I(data_in_4_0));
    InMux I__6694 (
            .O(N__29140),
            .I(N__29136));
    InMux I__6693 (
            .O(N__29139),
            .I(N__29133));
    LocalMux I__6692 (
            .O(N__29136),
            .I(N__29130));
    LocalMux I__6691 (
            .O(N__29133),
            .I(N__29126));
    Span4Mux_h I__6690 (
            .O(N__29130),
            .I(N__29123));
    InMux I__6689 (
            .O(N__29129),
            .I(N__29120));
    Span4Mux_v I__6688 (
            .O(N__29126),
            .I(N__29115));
    Span4Mux_v I__6687 (
            .O(N__29123),
            .I(N__29115));
    LocalMux I__6686 (
            .O(N__29120),
            .I(N__29110));
    Span4Mux_h I__6685 (
            .O(N__29115),
            .I(N__29107));
    InMux I__6684 (
            .O(N__29114),
            .I(N__29102));
    InMux I__6683 (
            .O(N__29113),
            .I(N__29102));
    Odrv12 I__6682 (
            .O(N__29110),
            .I(\c0.data_in_field_32 ));
    Odrv4 I__6681 (
            .O(N__29107),
            .I(\c0.data_in_field_32 ));
    LocalMux I__6680 (
            .O(N__29102),
            .I(\c0.data_in_field_32 ));
    CascadeMux I__6679 (
            .O(N__29095),
            .I(N__29092));
    InMux I__6678 (
            .O(N__29092),
            .I(N__29088));
    InMux I__6677 (
            .O(N__29091),
            .I(N__29085));
    LocalMux I__6676 (
            .O(N__29088),
            .I(N__29082));
    LocalMux I__6675 (
            .O(N__29085),
            .I(N__29079));
    Span4Mux_v I__6674 (
            .O(N__29082),
            .I(N__29073));
    Span4Mux_h I__6673 (
            .O(N__29079),
            .I(N__29073));
    InMux I__6672 (
            .O(N__29078),
            .I(N__29070));
    Odrv4 I__6671 (
            .O(N__29073),
            .I(data_in_13_2));
    LocalMux I__6670 (
            .O(N__29070),
            .I(data_in_13_2));
    CascadeMux I__6669 (
            .O(N__29065),
            .I(N__29062));
    InMux I__6668 (
            .O(N__29062),
            .I(N__29059));
    LocalMux I__6667 (
            .O(N__29059),
            .I(N__29056));
    Span4Mux_h I__6666 (
            .O(N__29056),
            .I(N__29052));
    InMux I__6665 (
            .O(N__29055),
            .I(N__29049));
    Span4Mux_v I__6664 (
            .O(N__29052),
            .I(N__29044));
    LocalMux I__6663 (
            .O(N__29049),
            .I(N__29044));
    Span4Mux_h I__6662 (
            .O(N__29044),
            .I(N__29040));
    InMux I__6661 (
            .O(N__29043),
            .I(N__29037));
    Odrv4 I__6660 (
            .O(N__29040),
            .I(data_in_12_2));
    LocalMux I__6659 (
            .O(N__29037),
            .I(data_in_12_2));
    InMux I__6658 (
            .O(N__29032),
            .I(N__29026));
    InMux I__6657 (
            .O(N__29031),
            .I(N__29023));
    InMux I__6656 (
            .O(N__29030),
            .I(N__29020));
    InMux I__6655 (
            .O(N__29029),
            .I(N__29016));
    LocalMux I__6654 (
            .O(N__29026),
            .I(N__29012));
    LocalMux I__6653 (
            .O(N__29023),
            .I(N__29009));
    LocalMux I__6652 (
            .O(N__29020),
            .I(N__29006));
    InMux I__6651 (
            .O(N__29019),
            .I(N__29003));
    LocalMux I__6650 (
            .O(N__29016),
            .I(N__29000));
    InMux I__6649 (
            .O(N__29015),
            .I(N__28997));
    Span4Mux_h I__6648 (
            .O(N__29012),
            .I(N__28994));
    Span4Mux_h I__6647 (
            .O(N__29009),
            .I(N__28991));
    Span12Mux_v I__6646 (
            .O(N__29006),
            .I(N__28984));
    LocalMux I__6645 (
            .O(N__29003),
            .I(N__28984));
    Sp12to4 I__6644 (
            .O(N__29000),
            .I(N__28984));
    LocalMux I__6643 (
            .O(N__28997),
            .I(\c0.data_in_field_64 ));
    Odrv4 I__6642 (
            .O(N__28994),
            .I(\c0.data_in_field_64 ));
    Odrv4 I__6641 (
            .O(N__28991),
            .I(\c0.data_in_field_64 ));
    Odrv12 I__6640 (
            .O(N__28984),
            .I(\c0.data_in_field_64 ));
    InMux I__6639 (
            .O(N__28975),
            .I(N__28970));
    InMux I__6638 (
            .O(N__28974),
            .I(N__28965));
    InMux I__6637 (
            .O(N__28973),
            .I(N__28965));
    LocalMux I__6636 (
            .O(N__28970),
            .I(\c0.n5179 ));
    LocalMux I__6635 (
            .O(N__28965),
            .I(\c0.n5179 ));
    InMux I__6634 (
            .O(N__28960),
            .I(N__28956));
    InMux I__6633 (
            .O(N__28959),
            .I(N__28951));
    LocalMux I__6632 (
            .O(N__28956),
            .I(N__28948));
    InMux I__6631 (
            .O(N__28955),
            .I(N__28945));
    InMux I__6630 (
            .O(N__28954),
            .I(N__28942));
    LocalMux I__6629 (
            .O(N__28951),
            .I(N__28939));
    Span4Mux_h I__6628 (
            .O(N__28948),
            .I(N__28936));
    LocalMux I__6627 (
            .O(N__28945),
            .I(N__28933));
    LocalMux I__6626 (
            .O(N__28942),
            .I(\c0.data_in_field_46 ));
    Odrv4 I__6625 (
            .O(N__28939),
            .I(\c0.data_in_field_46 ));
    Odrv4 I__6624 (
            .O(N__28936),
            .I(\c0.data_in_field_46 ));
    Odrv4 I__6623 (
            .O(N__28933),
            .I(\c0.data_in_field_46 ));
    CascadeMux I__6622 (
            .O(N__28924),
            .I(N__28921));
    InMux I__6621 (
            .O(N__28921),
            .I(N__28918));
    LocalMux I__6620 (
            .O(N__28918),
            .I(N__28911));
    InMux I__6619 (
            .O(N__28917),
            .I(N__28908));
    InMux I__6618 (
            .O(N__28916),
            .I(N__28905));
    InMux I__6617 (
            .O(N__28915),
            .I(N__28902));
    InMux I__6616 (
            .O(N__28914),
            .I(N__28899));
    Span12Mux_s6_v I__6615 (
            .O(N__28911),
            .I(N__28896));
    LocalMux I__6614 (
            .O(N__28908),
            .I(\c0.data_in_field_4 ));
    LocalMux I__6613 (
            .O(N__28905),
            .I(\c0.data_in_field_4 ));
    LocalMux I__6612 (
            .O(N__28902),
            .I(\c0.data_in_field_4 ));
    LocalMux I__6611 (
            .O(N__28899),
            .I(\c0.data_in_field_4 ));
    Odrv12 I__6610 (
            .O(N__28896),
            .I(\c0.data_in_field_4 ));
    CascadeMux I__6609 (
            .O(N__28885),
            .I(\c0.n1767_cascade_ ));
    InMux I__6608 (
            .O(N__28882),
            .I(N__28879));
    LocalMux I__6607 (
            .O(N__28879),
            .I(N__28875));
    InMux I__6606 (
            .O(N__28878),
            .I(N__28872));
    Odrv4 I__6605 (
            .O(N__28875),
            .I(\c0.n1899 ));
    LocalMux I__6604 (
            .O(N__28872),
            .I(\c0.n1899 ));
    InMux I__6603 (
            .O(N__28867),
            .I(N__28864));
    LocalMux I__6602 (
            .O(N__28864),
            .I(\c0.n5126 ));
    InMux I__6601 (
            .O(N__28861),
            .I(N__28858));
    LocalMux I__6600 (
            .O(N__28858),
            .I(N__28855));
    Span4Mux_h I__6599 (
            .O(N__28855),
            .I(N__28850));
    InMux I__6598 (
            .O(N__28854),
            .I(N__28845));
    InMux I__6597 (
            .O(N__28853),
            .I(N__28841));
    Span4Mux_h I__6596 (
            .O(N__28850),
            .I(N__28838));
    InMux I__6595 (
            .O(N__28849),
            .I(N__28835));
    InMux I__6594 (
            .O(N__28848),
            .I(N__28832));
    LocalMux I__6593 (
            .O(N__28845),
            .I(N__28829));
    InMux I__6592 (
            .O(N__28844),
            .I(N__28826));
    LocalMux I__6591 (
            .O(N__28841),
            .I(\c0.data_in_field_140 ));
    Odrv4 I__6590 (
            .O(N__28838),
            .I(\c0.data_in_field_140 ));
    LocalMux I__6589 (
            .O(N__28835),
            .I(\c0.data_in_field_140 ));
    LocalMux I__6588 (
            .O(N__28832),
            .I(\c0.data_in_field_140 ));
    Odrv4 I__6587 (
            .O(N__28829),
            .I(\c0.data_in_field_140 ));
    LocalMux I__6586 (
            .O(N__28826),
            .I(\c0.data_in_field_140 ));
    CascadeMux I__6585 (
            .O(N__28813),
            .I(\c0.n5126_cascade_ ));
    InMux I__6584 (
            .O(N__28810),
            .I(N__28805));
    InMux I__6583 (
            .O(N__28809),
            .I(N__28802));
    InMux I__6582 (
            .O(N__28808),
            .I(N__28799));
    LocalMux I__6581 (
            .O(N__28805),
            .I(N__28796));
    LocalMux I__6580 (
            .O(N__28802),
            .I(N__28793));
    LocalMux I__6579 (
            .O(N__28799),
            .I(N__28790));
    Span4Mux_h I__6578 (
            .O(N__28796),
            .I(N__28783));
    Span4Mux_v I__6577 (
            .O(N__28793),
            .I(N__28783));
    Span4Mux_h I__6576 (
            .O(N__28790),
            .I(N__28780));
    InMux I__6575 (
            .O(N__28789),
            .I(N__28777));
    CascadeMux I__6574 (
            .O(N__28788),
            .I(N__28774));
    Span4Mux_h I__6573 (
            .O(N__28783),
            .I(N__28769));
    Span4Mux_v I__6572 (
            .O(N__28780),
            .I(N__28769));
    LocalMux I__6571 (
            .O(N__28777),
            .I(N__28766));
    InMux I__6570 (
            .O(N__28774),
            .I(N__28763));
    Odrv4 I__6569 (
            .O(N__28769),
            .I(\c0.data_in_field_125 ));
    Odrv4 I__6568 (
            .O(N__28766),
            .I(\c0.data_in_field_125 ));
    LocalMux I__6567 (
            .O(N__28763),
            .I(\c0.data_in_field_125 ));
    InMux I__6566 (
            .O(N__28756),
            .I(N__28753));
    LocalMux I__6565 (
            .O(N__28753),
            .I(N__28750));
    Span4Mux_h I__6564 (
            .O(N__28750),
            .I(N__28747));
    Span4Mux_h I__6563 (
            .O(N__28747),
            .I(N__28744));
    Odrv4 I__6562 (
            .O(N__28744),
            .I(\c0.n20_adj_1899 ));
    CascadeMux I__6561 (
            .O(N__28741),
            .I(N__28738));
    InMux I__6560 (
            .O(N__28738),
            .I(N__28734));
    InMux I__6559 (
            .O(N__28737),
            .I(N__28731));
    LocalMux I__6558 (
            .O(N__28734),
            .I(N__28726));
    LocalMux I__6557 (
            .O(N__28731),
            .I(N__28726));
    Span4Mux_h I__6556 (
            .O(N__28726),
            .I(N__28722));
    InMux I__6555 (
            .O(N__28725),
            .I(N__28719));
    Odrv4 I__6554 (
            .O(N__28722),
            .I(data_in_14_6));
    LocalMux I__6553 (
            .O(N__28719),
            .I(data_in_14_6));
    InMux I__6552 (
            .O(N__28714),
            .I(N__28711));
    LocalMux I__6551 (
            .O(N__28711),
            .I(\c0.n10_adj_1872 ));
    InMux I__6550 (
            .O(N__28708),
            .I(N__28704));
    CascadeMux I__6549 (
            .O(N__28707),
            .I(N__28701));
    LocalMux I__6548 (
            .O(N__28704),
            .I(N__28698));
    InMux I__6547 (
            .O(N__28701),
            .I(N__28695));
    Span4Mux_h I__6546 (
            .O(N__28698),
            .I(N__28692));
    LocalMux I__6545 (
            .O(N__28695),
            .I(N__28689));
    Span4Mux_v I__6544 (
            .O(N__28692),
            .I(N__28686));
    Span4Mux_h I__6543 (
            .O(N__28689),
            .I(N__28682));
    Span4Mux_h I__6542 (
            .O(N__28686),
            .I(N__28679));
    InMux I__6541 (
            .O(N__28685),
            .I(N__28676));
    Odrv4 I__6540 (
            .O(N__28682),
            .I(data_in_12_4));
    Odrv4 I__6539 (
            .O(N__28679),
            .I(data_in_12_4));
    LocalMux I__6538 (
            .O(N__28676),
            .I(data_in_12_4));
    InMux I__6537 (
            .O(N__28669),
            .I(N__28666));
    LocalMux I__6536 (
            .O(N__28666),
            .I(N__28662));
    InMux I__6535 (
            .O(N__28665),
            .I(N__28659));
    Span4Mux_v I__6534 (
            .O(N__28662),
            .I(N__28656));
    LocalMux I__6533 (
            .O(N__28659),
            .I(N__28651));
    Span4Mux_h I__6532 (
            .O(N__28656),
            .I(N__28648));
    InMux I__6531 (
            .O(N__28655),
            .I(N__28643));
    InMux I__6530 (
            .O(N__28654),
            .I(N__28643));
    Odrv4 I__6529 (
            .O(N__28651),
            .I(\c0.data_in_field_100 ));
    Odrv4 I__6528 (
            .O(N__28648),
            .I(\c0.data_in_field_100 ));
    LocalMux I__6527 (
            .O(N__28643),
            .I(\c0.data_in_field_100 ));
    InMux I__6526 (
            .O(N__28636),
            .I(N__28632));
    InMux I__6525 (
            .O(N__28635),
            .I(N__28627));
    LocalMux I__6524 (
            .O(N__28632),
            .I(N__28624));
    InMux I__6523 (
            .O(N__28631),
            .I(N__28621));
    InMux I__6522 (
            .O(N__28630),
            .I(N__28618));
    LocalMux I__6521 (
            .O(N__28627),
            .I(\c0.data_in_field_40 ));
    Odrv4 I__6520 (
            .O(N__28624),
            .I(\c0.data_in_field_40 ));
    LocalMux I__6519 (
            .O(N__28621),
            .I(\c0.data_in_field_40 ));
    LocalMux I__6518 (
            .O(N__28618),
            .I(\c0.data_in_field_40 ));
    CascadeMux I__6517 (
            .O(N__28609),
            .I(N__28605));
    InMux I__6516 (
            .O(N__28608),
            .I(N__28602));
    InMux I__6515 (
            .O(N__28605),
            .I(N__28599));
    LocalMux I__6514 (
            .O(N__28602),
            .I(N__28596));
    LocalMux I__6513 (
            .O(N__28599),
            .I(N__28593));
    Span4Mux_h I__6512 (
            .O(N__28596),
            .I(N__28590));
    Span4Mux_h I__6511 (
            .O(N__28593),
            .I(N__28586));
    Span4Mux_h I__6510 (
            .O(N__28590),
            .I(N__28583));
    InMux I__6509 (
            .O(N__28589),
            .I(N__28580));
    Odrv4 I__6508 (
            .O(N__28586),
            .I(data_in_11_1));
    Odrv4 I__6507 (
            .O(N__28583),
            .I(data_in_11_1));
    LocalMux I__6506 (
            .O(N__28580),
            .I(data_in_11_1));
    InMux I__6505 (
            .O(N__28573),
            .I(N__28570));
    LocalMux I__6504 (
            .O(N__28570),
            .I(N__28567));
    Span4Mux_h I__6503 (
            .O(N__28567),
            .I(N__28564));
    Span4Mux_h I__6502 (
            .O(N__28564),
            .I(N__28559));
    InMux I__6501 (
            .O(N__28563),
            .I(N__28556));
    InMux I__6500 (
            .O(N__28562),
            .I(N__28553));
    Span4Mux_v I__6499 (
            .O(N__28559),
            .I(N__28550));
    LocalMux I__6498 (
            .O(N__28556),
            .I(data_in_10_1));
    LocalMux I__6497 (
            .O(N__28553),
            .I(data_in_10_1));
    Odrv4 I__6496 (
            .O(N__28550),
            .I(data_in_10_1));
    CascadeMux I__6495 (
            .O(N__28543),
            .I(N__28540));
    InMux I__6494 (
            .O(N__28540),
            .I(N__28537));
    LocalMux I__6493 (
            .O(N__28537),
            .I(N__28533));
    InMux I__6492 (
            .O(N__28536),
            .I(N__28530));
    Span4Mux_v I__6491 (
            .O(N__28533),
            .I(N__28527));
    LocalMux I__6490 (
            .O(N__28530),
            .I(N__28524));
    Span4Mux_v I__6489 (
            .O(N__28527),
            .I(N__28518));
    Span4Mux_h I__6488 (
            .O(N__28524),
            .I(N__28518));
    InMux I__6487 (
            .O(N__28523),
            .I(N__28515));
    Odrv4 I__6486 (
            .O(N__28518),
            .I(data_in_11_0));
    LocalMux I__6485 (
            .O(N__28515),
            .I(data_in_11_0));
    InMux I__6484 (
            .O(N__28510),
            .I(N__28506));
    CascadeMux I__6483 (
            .O(N__28509),
            .I(N__28502));
    LocalMux I__6482 (
            .O(N__28506),
            .I(N__28499));
    CascadeMux I__6481 (
            .O(N__28505),
            .I(N__28496));
    InMux I__6480 (
            .O(N__28502),
            .I(N__28493));
    Span4Mux_h I__6479 (
            .O(N__28499),
            .I(N__28490));
    InMux I__6478 (
            .O(N__28496),
            .I(N__28487));
    LocalMux I__6477 (
            .O(N__28493),
            .I(\c0.data_in_field_14 ));
    Odrv4 I__6476 (
            .O(N__28490),
            .I(\c0.data_in_field_14 ));
    LocalMux I__6475 (
            .O(N__28487),
            .I(\c0.data_in_field_14 ));
    CascadeMux I__6474 (
            .O(N__28480),
            .I(N__28477));
    InMux I__6473 (
            .O(N__28477),
            .I(N__28474));
    LocalMux I__6472 (
            .O(N__28474),
            .I(N__28471));
    Span4Mux_h I__6471 (
            .O(N__28471),
            .I(N__28468));
    Span4Mux_h I__6470 (
            .O(N__28468),
            .I(N__28465));
    Odrv4 I__6469 (
            .O(N__28465),
            .I(\c0.n5911 ));
    InMux I__6468 (
            .O(N__28462),
            .I(N__28459));
    LocalMux I__6467 (
            .O(N__28459),
            .I(N__28453));
    InMux I__6466 (
            .O(N__28458),
            .I(N__28448));
    InMux I__6465 (
            .O(N__28457),
            .I(N__28448));
    InMux I__6464 (
            .O(N__28456),
            .I(N__28445));
    Odrv4 I__6463 (
            .O(N__28453),
            .I(\c0.data_in_field_6 ));
    LocalMux I__6462 (
            .O(N__28448),
            .I(\c0.data_in_field_6 ));
    LocalMux I__6461 (
            .O(N__28445),
            .I(\c0.data_in_field_6 ));
    InMux I__6460 (
            .O(N__28438),
            .I(N__28434));
    InMux I__6459 (
            .O(N__28437),
            .I(N__28431));
    LocalMux I__6458 (
            .O(N__28434),
            .I(N__28428));
    LocalMux I__6457 (
            .O(N__28431),
            .I(N__28425));
    Span4Mux_v I__6456 (
            .O(N__28428),
            .I(N__28419));
    Span4Mux_s3_h I__6455 (
            .O(N__28425),
            .I(N__28419));
    InMux I__6454 (
            .O(N__28424),
            .I(N__28416));
    Span4Mux_h I__6453 (
            .O(N__28419),
            .I(N__28411));
    LocalMux I__6452 (
            .O(N__28416),
            .I(N__28411));
    Span4Mux_h I__6451 (
            .O(N__28411),
            .I(N__28406));
    InMux I__6450 (
            .O(N__28410),
            .I(N__28401));
    InMux I__6449 (
            .O(N__28409),
            .I(N__28401));
    Odrv4 I__6448 (
            .O(N__28406),
            .I(\c0.data_in_field_138 ));
    LocalMux I__6447 (
            .O(N__28401),
            .I(\c0.data_in_field_138 ));
    InMux I__6446 (
            .O(N__28396),
            .I(N__28392));
    InMux I__6445 (
            .O(N__28395),
            .I(N__28389));
    LocalMux I__6444 (
            .O(N__28392),
            .I(N__28386));
    LocalMux I__6443 (
            .O(N__28389),
            .I(N__28383));
    Span4Mux_s3_h I__6442 (
            .O(N__28386),
            .I(N__28377));
    Span4Mux_v I__6441 (
            .O(N__28383),
            .I(N__28377));
    CascadeMux I__6440 (
            .O(N__28382),
            .I(N__28374));
    Span4Mux_h I__6439 (
            .O(N__28377),
            .I(N__28371));
    InMux I__6438 (
            .O(N__28374),
            .I(N__28368));
    Span4Mux_h I__6437 (
            .O(N__28371),
            .I(N__28361));
    LocalMux I__6436 (
            .O(N__28368),
            .I(N__28361));
    InMux I__6435 (
            .O(N__28367),
            .I(N__28356));
    InMux I__6434 (
            .O(N__28366),
            .I(N__28356));
    Odrv4 I__6433 (
            .O(N__28361),
            .I(\c0.data_in_field_130 ));
    LocalMux I__6432 (
            .O(N__28356),
            .I(\c0.data_in_field_130 ));
    InMux I__6431 (
            .O(N__28351),
            .I(N__28348));
    LocalMux I__6430 (
            .O(N__28348),
            .I(N__28345));
    Span4Mux_h I__6429 (
            .O(N__28345),
            .I(N__28342));
    Span4Mux_h I__6428 (
            .O(N__28342),
            .I(N__28339));
    Odrv4 I__6427 (
            .O(N__28339),
            .I(\c0.n5123 ));
    CascadeMux I__6426 (
            .O(N__28336),
            .I(\c0.n5123_cascade_ ));
    InMux I__6425 (
            .O(N__28333),
            .I(N__28330));
    LocalMux I__6424 (
            .O(N__28330),
            .I(N__28327));
    Span4Mux_h I__6423 (
            .O(N__28327),
            .I(N__28323));
    InMux I__6422 (
            .O(N__28326),
            .I(N__28320));
    Span4Mux_h I__6421 (
            .O(N__28323),
            .I(N__28317));
    LocalMux I__6420 (
            .O(N__28320),
            .I(N__28314));
    Span4Mux_h I__6419 (
            .O(N__28317),
            .I(N__28311));
    Odrv12 I__6418 (
            .O(N__28314),
            .I(\c0.n5231 ));
    Odrv4 I__6417 (
            .O(N__28311),
            .I(\c0.n5231 ));
    InMux I__6416 (
            .O(N__28306),
            .I(N__28301));
    InMux I__6415 (
            .O(N__28305),
            .I(N__28298));
    InMux I__6414 (
            .O(N__28304),
            .I(N__28295));
    LocalMux I__6413 (
            .O(N__28301),
            .I(N__28291));
    LocalMux I__6412 (
            .O(N__28298),
            .I(N__28288));
    LocalMux I__6411 (
            .O(N__28295),
            .I(N__28285));
    InMux I__6410 (
            .O(N__28294),
            .I(N__28281));
    Span4Mux_h I__6409 (
            .O(N__28291),
            .I(N__28278));
    Span4Mux_v I__6408 (
            .O(N__28288),
            .I(N__28273));
    Span4Mux_h I__6407 (
            .O(N__28285),
            .I(N__28273));
    InMux I__6406 (
            .O(N__28284),
            .I(N__28270));
    LocalMux I__6405 (
            .O(N__28281),
            .I(\c0.data_in_field_58 ));
    Odrv4 I__6404 (
            .O(N__28278),
            .I(\c0.data_in_field_58 ));
    Odrv4 I__6403 (
            .O(N__28273),
            .I(\c0.data_in_field_58 ));
    LocalMux I__6402 (
            .O(N__28270),
            .I(\c0.data_in_field_58 ));
    CascadeMux I__6401 (
            .O(N__28261),
            .I(\c0.n5773_cascade_ ));
    InMux I__6400 (
            .O(N__28258),
            .I(N__28254));
    InMux I__6399 (
            .O(N__28257),
            .I(N__28251));
    LocalMux I__6398 (
            .O(N__28254),
            .I(N__28246));
    LocalMux I__6397 (
            .O(N__28251),
            .I(N__28243));
    InMux I__6396 (
            .O(N__28250),
            .I(N__28240));
    InMux I__6395 (
            .O(N__28249),
            .I(N__28237));
    Span4Mux_v I__6394 (
            .O(N__28246),
            .I(N__28234));
    Span4Mux_h I__6393 (
            .O(N__28243),
            .I(N__28231));
    LocalMux I__6392 (
            .O(N__28240),
            .I(N__28228));
    LocalMux I__6391 (
            .O(N__28237),
            .I(\c0.data_in_field_34 ));
    Odrv4 I__6390 (
            .O(N__28234),
            .I(\c0.data_in_field_34 ));
    Odrv4 I__6389 (
            .O(N__28231),
            .I(\c0.data_in_field_34 ));
    Odrv12 I__6388 (
            .O(N__28228),
            .I(\c0.data_in_field_34 ));
    InMux I__6387 (
            .O(N__28219),
            .I(N__28216));
    LocalMux I__6386 (
            .O(N__28216),
            .I(N__28213));
    Span4Mux_h I__6385 (
            .O(N__28213),
            .I(N__28210));
    Odrv4 I__6384 (
            .O(N__28210),
            .I(\c0.n5441 ));
    InMux I__6383 (
            .O(N__28207),
            .I(N__28204));
    LocalMux I__6382 (
            .O(N__28204),
            .I(N__28201));
    Span12Mux_v I__6381 (
            .O(N__28201),
            .I(N__28198));
    Odrv12 I__6380 (
            .O(N__28198),
            .I(\c0.n5477 ));
    CascadeMux I__6379 (
            .O(N__28195),
            .I(N__28192));
    InMux I__6378 (
            .O(N__28192),
            .I(N__28189));
    LocalMux I__6377 (
            .O(N__28189),
            .I(N__28185));
    InMux I__6376 (
            .O(N__28188),
            .I(N__28182));
    Span4Mux_h I__6375 (
            .O(N__28185),
            .I(N__28179));
    LocalMux I__6374 (
            .O(N__28182),
            .I(N__28173));
    Span4Mux_h I__6373 (
            .O(N__28179),
            .I(N__28173));
    InMux I__6372 (
            .O(N__28178),
            .I(N__28170));
    Span4Mux_v I__6371 (
            .O(N__28173),
            .I(N__28167));
    LocalMux I__6370 (
            .O(N__28170),
            .I(data_in_16_4));
    Odrv4 I__6369 (
            .O(N__28167),
            .I(data_in_16_4));
    CascadeMux I__6368 (
            .O(N__28162),
            .I(N__28159));
    InMux I__6367 (
            .O(N__28159),
            .I(N__28156));
    LocalMux I__6366 (
            .O(N__28156),
            .I(N__28152));
    CascadeMux I__6365 (
            .O(N__28155),
            .I(N__28149));
    Span4Mux_h I__6364 (
            .O(N__28152),
            .I(N__28145));
    InMux I__6363 (
            .O(N__28149),
            .I(N__28140));
    InMux I__6362 (
            .O(N__28148),
            .I(N__28140));
    Span4Mux_h I__6361 (
            .O(N__28145),
            .I(N__28137));
    LocalMux I__6360 (
            .O(N__28140),
            .I(data_in_15_4));
    Odrv4 I__6359 (
            .O(N__28137),
            .I(data_in_15_4));
    CascadeMux I__6358 (
            .O(N__28132),
            .I(N__28127));
    InMux I__6357 (
            .O(N__28131),
            .I(N__28124));
    InMux I__6356 (
            .O(N__28130),
            .I(N__28121));
    InMux I__6355 (
            .O(N__28127),
            .I(N__28118));
    LocalMux I__6354 (
            .O(N__28124),
            .I(N__28115));
    LocalMux I__6353 (
            .O(N__28121),
            .I(data_in_8_6));
    LocalMux I__6352 (
            .O(N__28118),
            .I(data_in_8_6));
    Odrv4 I__6351 (
            .O(N__28115),
            .I(data_in_8_6));
    InMux I__6350 (
            .O(N__28108),
            .I(N__28104));
    InMux I__6349 (
            .O(N__28107),
            .I(N__28101));
    LocalMux I__6348 (
            .O(N__28104),
            .I(N__28097));
    LocalMux I__6347 (
            .O(N__28101),
            .I(N__28094));
    InMux I__6346 (
            .O(N__28100),
            .I(N__28091));
    Span4Mux_h I__6345 (
            .O(N__28097),
            .I(N__28088));
    Span4Mux_h I__6344 (
            .O(N__28094),
            .I(N__28085));
    LocalMux I__6343 (
            .O(N__28091),
            .I(data_in_6_5));
    Odrv4 I__6342 (
            .O(N__28088),
            .I(data_in_6_5));
    Odrv4 I__6341 (
            .O(N__28085),
            .I(data_in_6_5));
    InMux I__6340 (
            .O(N__28078),
            .I(N__28075));
    LocalMux I__6339 (
            .O(N__28075),
            .I(N__28070));
    InMux I__6338 (
            .O(N__28074),
            .I(N__28067));
    InMux I__6337 (
            .O(N__28073),
            .I(N__28064));
    Odrv4 I__6336 (
            .O(N__28070),
            .I(data_in_4_6));
    LocalMux I__6335 (
            .O(N__28067),
            .I(data_in_4_6));
    LocalMux I__6334 (
            .O(N__28064),
            .I(data_in_4_6));
    InMux I__6333 (
            .O(N__28057),
            .I(N__28054));
    LocalMux I__6332 (
            .O(N__28054),
            .I(N__28051));
    Span4Mux_h I__6331 (
            .O(N__28051),
            .I(N__28047));
    CascadeMux I__6330 (
            .O(N__28050),
            .I(N__28043));
    Sp12to4 I__6329 (
            .O(N__28047),
            .I(N__28040));
    InMux I__6328 (
            .O(N__28046),
            .I(N__28035));
    InMux I__6327 (
            .O(N__28043),
            .I(N__28035));
    Odrv12 I__6326 (
            .O(N__28040),
            .I(data_in_6_0));
    LocalMux I__6325 (
            .O(N__28035),
            .I(data_in_6_0));
    InMux I__6324 (
            .O(N__28030),
            .I(N__28026));
    InMux I__6323 (
            .O(N__28029),
            .I(N__28021));
    LocalMux I__6322 (
            .O(N__28026),
            .I(N__28018));
    InMux I__6321 (
            .O(N__28025),
            .I(N__28015));
    InMux I__6320 (
            .O(N__28024),
            .I(N__28012));
    LocalMux I__6319 (
            .O(N__28021),
            .I(N__28009));
    Span4Mux_v I__6318 (
            .O(N__28018),
            .I(N__28004));
    LocalMux I__6317 (
            .O(N__28015),
            .I(N__28004));
    LocalMux I__6316 (
            .O(N__28012),
            .I(N__28000));
    Span4Mux_v I__6315 (
            .O(N__28009),
            .I(N__27995));
    Span4Mux_h I__6314 (
            .O(N__28004),
            .I(N__27995));
    InMux I__6313 (
            .O(N__28003),
            .I(N__27991));
    Span12Mux_v I__6312 (
            .O(N__28000),
            .I(N__27988));
    Span4Mux_h I__6311 (
            .O(N__27995),
            .I(N__27985));
    InMux I__6310 (
            .O(N__27994),
            .I(N__27982));
    LocalMux I__6309 (
            .O(N__27991),
            .I(\c0.data_in_field_60 ));
    Odrv12 I__6308 (
            .O(N__27988),
            .I(\c0.data_in_field_60 ));
    Odrv4 I__6307 (
            .O(N__27985),
            .I(\c0.data_in_field_60 ));
    LocalMux I__6306 (
            .O(N__27982),
            .I(\c0.data_in_field_60 ));
    InMux I__6305 (
            .O(N__27973),
            .I(N__27970));
    LocalMux I__6304 (
            .O(N__27970),
            .I(\c0.n6_adj_1875 ));
    InMux I__6303 (
            .O(N__27967),
            .I(N__27963));
    InMux I__6302 (
            .O(N__27966),
            .I(N__27960));
    LocalMux I__6301 (
            .O(N__27963),
            .I(N__27957));
    LocalMux I__6300 (
            .O(N__27960),
            .I(N__27953));
    Span4Mux_s2_v I__6299 (
            .O(N__27957),
            .I(N__27950));
    InMux I__6298 (
            .O(N__27956),
            .I(N__27946));
    Span4Mux_h I__6297 (
            .O(N__27953),
            .I(N__27943));
    Span4Mux_h I__6296 (
            .O(N__27950),
            .I(N__27940));
    InMux I__6295 (
            .O(N__27949),
            .I(N__27937));
    LocalMux I__6294 (
            .O(N__27946),
            .I(data_in_3_5));
    Odrv4 I__6293 (
            .O(N__27943),
            .I(data_in_3_5));
    Odrv4 I__6292 (
            .O(N__27940),
            .I(data_in_3_5));
    LocalMux I__6291 (
            .O(N__27937),
            .I(data_in_3_5));
    InMux I__6290 (
            .O(N__27928),
            .I(N__27923));
    CascadeMux I__6289 (
            .O(N__27927),
            .I(N__27920));
    InMux I__6288 (
            .O(N__27926),
            .I(N__27916));
    LocalMux I__6287 (
            .O(N__27923),
            .I(N__27913));
    InMux I__6286 (
            .O(N__27920),
            .I(N__27910));
    InMux I__6285 (
            .O(N__27919),
            .I(N__27907));
    LocalMux I__6284 (
            .O(N__27916),
            .I(N__27904));
    Span4Mux_v I__6283 (
            .O(N__27913),
            .I(N__27899));
    LocalMux I__6282 (
            .O(N__27910),
            .I(N__27899));
    LocalMux I__6281 (
            .O(N__27907),
            .I(data_in_3_4));
    Odrv12 I__6280 (
            .O(N__27904),
            .I(data_in_3_4));
    Odrv4 I__6279 (
            .O(N__27899),
            .I(data_in_3_4));
    InMux I__6278 (
            .O(N__27892),
            .I(N__27888));
    InMux I__6277 (
            .O(N__27891),
            .I(N__27885));
    LocalMux I__6276 (
            .O(N__27888),
            .I(N__27882));
    LocalMux I__6275 (
            .O(N__27885),
            .I(N__27879));
    Span4Mux_h I__6274 (
            .O(N__27882),
            .I(N__27876));
    Span4Mux_h I__6273 (
            .O(N__27879),
            .I(N__27873));
    Span4Mux_h I__6272 (
            .O(N__27876),
            .I(N__27870));
    Span4Mux_h I__6271 (
            .O(N__27873),
            .I(N__27865));
    Sp12to4 I__6270 (
            .O(N__27870),
            .I(N__27862));
    InMux I__6269 (
            .O(N__27869),
            .I(N__27857));
    InMux I__6268 (
            .O(N__27868),
            .I(N__27857));
    Odrv4 I__6267 (
            .O(N__27865),
            .I(data_in_2_6));
    Odrv12 I__6266 (
            .O(N__27862),
            .I(data_in_2_6));
    LocalMux I__6265 (
            .O(N__27857),
            .I(data_in_2_6));
    CascadeMux I__6264 (
            .O(N__27850),
            .I(N__27847));
    InMux I__6263 (
            .O(N__27847),
            .I(N__27844));
    LocalMux I__6262 (
            .O(N__27844),
            .I(N__27841));
    Span4Mux_h I__6261 (
            .O(N__27841),
            .I(N__27838));
    Span4Mux_h I__6260 (
            .O(N__27838),
            .I(N__27832));
    InMux I__6259 (
            .O(N__27837),
            .I(N__27825));
    InMux I__6258 (
            .O(N__27836),
            .I(N__27825));
    InMux I__6257 (
            .O(N__27835),
            .I(N__27825));
    Odrv4 I__6256 (
            .O(N__27832),
            .I(data_in_3_6));
    LocalMux I__6255 (
            .O(N__27825),
            .I(data_in_3_6));
    CascadeMux I__6254 (
            .O(N__27820),
            .I(\c0.n28_adj_1953_cascade_ ));
    InMux I__6253 (
            .O(N__27817),
            .I(N__27814));
    LocalMux I__6252 (
            .O(N__27814),
            .I(\c0.n22_adj_1952 ));
    InMux I__6251 (
            .O(N__27811),
            .I(N__27808));
    LocalMux I__6250 (
            .O(N__27808),
            .I(N__27805));
    Odrv12 I__6249 (
            .O(N__27805),
            .I(\c0.n30_adj_1959 ));
    CascadeMux I__6248 (
            .O(N__27802),
            .I(N__27799));
    InMux I__6247 (
            .O(N__27799),
            .I(N__27796));
    LocalMux I__6246 (
            .O(N__27796),
            .I(N__27792));
    InMux I__6245 (
            .O(N__27795),
            .I(N__27789));
    Span4Mux_h I__6244 (
            .O(N__27792),
            .I(N__27785));
    LocalMux I__6243 (
            .O(N__27789),
            .I(N__27782));
    InMux I__6242 (
            .O(N__27788),
            .I(N__27779));
    Odrv4 I__6241 (
            .O(N__27785),
            .I(data_in_4_5));
    Odrv4 I__6240 (
            .O(N__27782),
            .I(data_in_4_5));
    LocalMux I__6239 (
            .O(N__27779),
            .I(data_in_4_5));
    CascadeMux I__6238 (
            .O(N__27772),
            .I(N__27769));
    InMux I__6237 (
            .O(N__27769),
            .I(N__27763));
    InMux I__6236 (
            .O(N__27768),
            .I(N__27763));
    LocalMux I__6235 (
            .O(N__27763),
            .I(N__27760));
    Span4Mux_h I__6234 (
            .O(N__27760),
            .I(N__27756));
    InMux I__6233 (
            .O(N__27759),
            .I(N__27753));
    Odrv4 I__6232 (
            .O(N__27756),
            .I(data_in_8_0));
    LocalMux I__6231 (
            .O(N__27753),
            .I(data_in_8_0));
    CascadeMux I__6230 (
            .O(N__27748),
            .I(N__27745));
    InMux I__6229 (
            .O(N__27745),
            .I(N__27741));
    InMux I__6228 (
            .O(N__27744),
            .I(N__27738));
    LocalMux I__6227 (
            .O(N__27741),
            .I(N__27734));
    LocalMux I__6226 (
            .O(N__27738),
            .I(N__27731));
    InMux I__6225 (
            .O(N__27737),
            .I(N__27728));
    Odrv12 I__6224 (
            .O(N__27734),
            .I(data_in_5_7));
    Odrv4 I__6223 (
            .O(N__27731),
            .I(data_in_5_7));
    LocalMux I__6222 (
            .O(N__27728),
            .I(data_in_5_7));
    InMux I__6221 (
            .O(N__27721),
            .I(N__27717));
    InMux I__6220 (
            .O(N__27720),
            .I(N__27714));
    LocalMux I__6219 (
            .O(N__27717),
            .I(N__27710));
    LocalMux I__6218 (
            .O(N__27714),
            .I(N__27707));
    InMux I__6217 (
            .O(N__27713),
            .I(N__27703));
    Span4Mux_h I__6216 (
            .O(N__27710),
            .I(N__27698));
    Span4Mux_v I__6215 (
            .O(N__27707),
            .I(N__27698));
    InMux I__6214 (
            .O(N__27706),
            .I(N__27695));
    LocalMux I__6213 (
            .O(N__27703),
            .I(\c0.data_in_field_47 ));
    Odrv4 I__6212 (
            .O(N__27698),
            .I(\c0.data_in_field_47 ));
    LocalMux I__6211 (
            .O(N__27695),
            .I(\c0.data_in_field_47 ));
    InMux I__6210 (
            .O(N__27688),
            .I(N__27684));
    CascadeMux I__6209 (
            .O(N__27687),
            .I(N__27681));
    LocalMux I__6208 (
            .O(N__27684),
            .I(N__27678));
    InMux I__6207 (
            .O(N__27681),
            .I(N__27674));
    Span4Mux_h I__6206 (
            .O(N__27678),
            .I(N__27671));
    InMux I__6205 (
            .O(N__27677),
            .I(N__27668));
    LocalMux I__6204 (
            .O(N__27674),
            .I(data_in_15_7));
    Odrv4 I__6203 (
            .O(N__27671),
            .I(data_in_15_7));
    LocalMux I__6202 (
            .O(N__27668),
            .I(data_in_15_7));
    InMux I__6201 (
            .O(N__27661),
            .I(N__27658));
    LocalMux I__6200 (
            .O(N__27658),
            .I(N__27654));
    InMux I__6199 (
            .O(N__27657),
            .I(N__27651));
    Span4Mux_h I__6198 (
            .O(N__27654),
            .I(N__27645));
    LocalMux I__6197 (
            .O(N__27651),
            .I(N__27645));
    InMux I__6196 (
            .O(N__27650),
            .I(N__27642));
    Span4Mux_v I__6195 (
            .O(N__27645),
            .I(N__27637));
    LocalMux I__6194 (
            .O(N__27642),
            .I(N__27634));
    InMux I__6193 (
            .O(N__27641),
            .I(N__27631));
    InMux I__6192 (
            .O(N__27640),
            .I(N__27628));
    Span4Mux_h I__6191 (
            .O(N__27637),
            .I(N__27625));
    Span4Mux_h I__6190 (
            .O(N__27634),
            .I(N__27622));
    LocalMux I__6189 (
            .O(N__27631),
            .I(\c0.data_in_field_127 ));
    LocalMux I__6188 (
            .O(N__27628),
            .I(\c0.data_in_field_127 ));
    Odrv4 I__6187 (
            .O(N__27625),
            .I(\c0.data_in_field_127 ));
    Odrv4 I__6186 (
            .O(N__27622),
            .I(\c0.data_in_field_127 ));
    InMux I__6185 (
            .O(N__27613),
            .I(N__27609));
    CascadeMux I__6184 (
            .O(N__27612),
            .I(N__27605));
    LocalMux I__6183 (
            .O(N__27609),
            .I(N__27602));
    InMux I__6182 (
            .O(N__27608),
            .I(N__27599));
    InMux I__6181 (
            .O(N__27605),
            .I(N__27596));
    Span4Mux_h I__6180 (
            .O(N__27602),
            .I(N__27593));
    LocalMux I__6179 (
            .O(N__27599),
            .I(data_in_16_0));
    LocalMux I__6178 (
            .O(N__27596),
            .I(data_in_16_0));
    Odrv4 I__6177 (
            .O(N__27593),
            .I(data_in_16_0));
    InMux I__6176 (
            .O(N__27586),
            .I(N__27582));
    CascadeMux I__6175 (
            .O(N__27585),
            .I(N__27579));
    LocalMux I__6174 (
            .O(N__27582),
            .I(N__27574));
    InMux I__6173 (
            .O(N__27579),
            .I(N__27571));
    InMux I__6172 (
            .O(N__27578),
            .I(N__27568));
    InMux I__6171 (
            .O(N__27577),
            .I(N__27565));
    Span12Mux_h I__6170 (
            .O(N__27574),
            .I(N__27562));
    LocalMux I__6169 (
            .O(N__27571),
            .I(N__27559));
    LocalMux I__6168 (
            .O(N__27568),
            .I(data_in_1_7));
    LocalMux I__6167 (
            .O(N__27565),
            .I(data_in_1_7));
    Odrv12 I__6166 (
            .O(N__27562),
            .I(data_in_1_7));
    Odrv4 I__6165 (
            .O(N__27559),
            .I(data_in_1_7));
    CascadeMux I__6164 (
            .O(N__27550),
            .I(N__27547));
    InMux I__6163 (
            .O(N__27547),
            .I(N__27543));
    InMux I__6162 (
            .O(N__27546),
            .I(N__27540));
    LocalMux I__6161 (
            .O(N__27543),
            .I(N__27537));
    LocalMux I__6160 (
            .O(N__27540),
            .I(N__27534));
    Span4Mux_v I__6159 (
            .O(N__27537),
            .I(N__27529));
    Span4Mux_v I__6158 (
            .O(N__27534),
            .I(N__27529));
    Sp12to4 I__6157 (
            .O(N__27529),
            .I(N__27525));
    InMux I__6156 (
            .O(N__27528),
            .I(N__27522));
    Odrv12 I__6155 (
            .O(N__27525),
            .I(data_in_10_5));
    LocalMux I__6154 (
            .O(N__27522),
            .I(data_in_10_5));
    InMux I__6153 (
            .O(N__27517),
            .I(N__27514));
    LocalMux I__6152 (
            .O(N__27514),
            .I(N__27510));
    InMux I__6151 (
            .O(N__27513),
            .I(N__27506));
    Span4Mux_h I__6150 (
            .O(N__27510),
            .I(N__27503));
    InMux I__6149 (
            .O(N__27509),
            .I(N__27500));
    LocalMux I__6148 (
            .O(N__27506),
            .I(data_in_9_5));
    Odrv4 I__6147 (
            .O(N__27503),
            .I(data_in_9_5));
    LocalMux I__6146 (
            .O(N__27500),
            .I(data_in_9_5));
    CascadeMux I__6145 (
            .O(N__27493),
            .I(N__27490));
    InMux I__6144 (
            .O(N__27490),
            .I(N__27485));
    InMux I__6143 (
            .O(N__27489),
            .I(N__27482));
    InMux I__6142 (
            .O(N__27488),
            .I(N__27479));
    LocalMux I__6141 (
            .O(N__27485),
            .I(N__27476));
    LocalMux I__6140 (
            .O(N__27482),
            .I(N__27473));
    LocalMux I__6139 (
            .O(N__27479),
            .I(data_in_0_5));
    Odrv4 I__6138 (
            .O(N__27476),
            .I(data_in_0_5));
    Odrv12 I__6137 (
            .O(N__27473),
            .I(data_in_0_5));
    InMux I__6136 (
            .O(N__27466),
            .I(N__27463));
    LocalMux I__6135 (
            .O(N__27463),
            .I(N__27460));
    Span4Mux_h I__6134 (
            .O(N__27460),
            .I(N__27457));
    Span4Mux_h I__6133 (
            .O(N__27457),
            .I(N__27451));
    InMux I__6132 (
            .O(N__27456),
            .I(N__27446));
    InMux I__6131 (
            .O(N__27455),
            .I(N__27446));
    InMux I__6130 (
            .O(N__27454),
            .I(N__27443));
    Odrv4 I__6129 (
            .O(N__27451),
            .I(data_in_1_2));
    LocalMux I__6128 (
            .O(N__27446),
            .I(data_in_1_2));
    LocalMux I__6127 (
            .O(N__27443),
            .I(data_in_1_2));
    CascadeMux I__6126 (
            .O(N__27436),
            .I(\c0.n6_adj_1876_cascade_ ));
    InMux I__6125 (
            .O(N__27433),
            .I(N__27430));
    LocalMux I__6124 (
            .O(N__27430),
            .I(N__27427));
    Span4Mux_v I__6123 (
            .O(N__27427),
            .I(N__27421));
    InMux I__6122 (
            .O(N__27426),
            .I(N__27418));
    InMux I__6121 (
            .O(N__27425),
            .I(N__27415));
    InMux I__6120 (
            .O(N__27424),
            .I(N__27411));
    Span4Mux_h I__6119 (
            .O(N__27421),
            .I(N__27406));
    LocalMux I__6118 (
            .O(N__27418),
            .I(N__27406));
    LocalMux I__6117 (
            .O(N__27415),
            .I(N__27403));
    InMux I__6116 (
            .O(N__27414),
            .I(N__27400));
    LocalMux I__6115 (
            .O(N__27411),
            .I(\c0.data_in_field_132 ));
    Odrv4 I__6114 (
            .O(N__27406),
            .I(\c0.data_in_field_132 ));
    Odrv12 I__6113 (
            .O(N__27403),
            .I(\c0.data_in_field_132 ));
    LocalMux I__6112 (
            .O(N__27400),
            .I(\c0.data_in_field_132 ));
    InMux I__6111 (
            .O(N__27391),
            .I(N__27388));
    LocalMux I__6110 (
            .O(N__27388),
            .I(N__27385));
    Span4Mux_h I__6109 (
            .O(N__27385),
            .I(N__27382));
    Span4Mux_h I__6108 (
            .O(N__27382),
            .I(N__27378));
    InMux I__6107 (
            .O(N__27381),
            .I(N__27375));
    Odrv4 I__6106 (
            .O(N__27378),
            .I(\c0.n5129 ));
    LocalMux I__6105 (
            .O(N__27375),
            .I(\c0.n5129 ));
    InMux I__6104 (
            .O(N__27370),
            .I(N__27367));
    LocalMux I__6103 (
            .O(N__27367),
            .I(N__27364));
    Odrv4 I__6102 (
            .O(N__27364),
            .I(\c0.n6_adj_1874 ));
    InMux I__6101 (
            .O(N__27361),
            .I(N__27358));
    LocalMux I__6100 (
            .O(N__27358),
            .I(N__27355));
    Span4Mux_h I__6099 (
            .O(N__27355),
            .I(N__27350));
    InMux I__6098 (
            .O(N__27354),
            .I(N__27345));
    InMux I__6097 (
            .O(N__27353),
            .I(N__27345));
    Odrv4 I__6096 (
            .O(N__27350),
            .I(data_in_0_0));
    LocalMux I__6095 (
            .O(N__27345),
            .I(data_in_0_0));
    InMux I__6094 (
            .O(N__27340),
            .I(N__27337));
    LocalMux I__6093 (
            .O(N__27337),
            .I(N__27331));
    InMux I__6092 (
            .O(N__27336),
            .I(N__27324));
    InMux I__6091 (
            .O(N__27335),
            .I(N__27324));
    InMux I__6090 (
            .O(N__27334),
            .I(N__27324));
    Odrv4 I__6089 (
            .O(N__27331),
            .I(\c0.data_in_field_0 ));
    LocalMux I__6088 (
            .O(N__27324),
            .I(\c0.data_in_field_0 ));
    InMux I__6087 (
            .O(N__27319),
            .I(N__27315));
    CascadeMux I__6086 (
            .O(N__27318),
            .I(N__27312));
    LocalMux I__6085 (
            .O(N__27315),
            .I(N__27307));
    InMux I__6084 (
            .O(N__27312),
            .I(N__27304));
    InMux I__6083 (
            .O(N__27311),
            .I(N__27301));
    CascadeMux I__6082 (
            .O(N__27310),
            .I(N__27298));
    Span4Mux_v I__6081 (
            .O(N__27307),
            .I(N__27291));
    LocalMux I__6080 (
            .O(N__27304),
            .I(N__27291));
    LocalMux I__6079 (
            .O(N__27301),
            .I(N__27288));
    InMux I__6078 (
            .O(N__27298),
            .I(N__27285));
    InMux I__6077 (
            .O(N__27297),
            .I(N__27282));
    InMux I__6076 (
            .O(N__27296),
            .I(N__27279));
    Span4Mux_h I__6075 (
            .O(N__27291),
            .I(N__27276));
    Span4Mux_h I__6074 (
            .O(N__27288),
            .I(N__27273));
    LocalMux I__6073 (
            .O(N__27285),
            .I(\c0.data_in_field_90 ));
    LocalMux I__6072 (
            .O(N__27282),
            .I(\c0.data_in_field_90 ));
    LocalMux I__6071 (
            .O(N__27279),
            .I(\c0.data_in_field_90 ));
    Odrv4 I__6070 (
            .O(N__27276),
            .I(\c0.data_in_field_90 ));
    Odrv4 I__6069 (
            .O(N__27273),
            .I(\c0.data_in_field_90 ));
    InMux I__6068 (
            .O(N__27262),
            .I(N__27259));
    LocalMux I__6067 (
            .O(N__27259),
            .I(N__27256));
    Span4Mux_h I__6066 (
            .O(N__27256),
            .I(N__27253));
    Odrv4 I__6065 (
            .O(N__27253),
            .I(\c0.n22_adj_1935 ));
    CascadeMux I__6064 (
            .O(N__27250),
            .I(N__27247));
    InMux I__6063 (
            .O(N__27247),
            .I(N__27244));
    LocalMux I__6062 (
            .O(N__27244),
            .I(N__27241));
    Span4Mux_h I__6061 (
            .O(N__27241),
            .I(N__27236));
    InMux I__6060 (
            .O(N__27240),
            .I(N__27231));
    InMux I__6059 (
            .O(N__27239),
            .I(N__27231));
    Odrv4 I__6058 (
            .O(N__27236),
            .I(data_in_5_6));
    LocalMux I__6057 (
            .O(N__27231),
            .I(data_in_5_6));
    InMux I__6056 (
            .O(N__27226),
            .I(N__27222));
    InMux I__6055 (
            .O(N__27225),
            .I(N__27219));
    LocalMux I__6054 (
            .O(N__27222),
            .I(N__27214));
    LocalMux I__6053 (
            .O(N__27219),
            .I(N__27211));
    InMux I__6052 (
            .O(N__27218),
            .I(N__27208));
    InMux I__6051 (
            .O(N__27217),
            .I(N__27205));
    Span4Mux_v I__6050 (
            .O(N__27214),
            .I(N__27202));
    Span12Mux_s9_h I__6049 (
            .O(N__27211),
            .I(N__27199));
    LocalMux I__6048 (
            .O(N__27208),
            .I(N__27196));
    LocalMux I__6047 (
            .O(N__27205),
            .I(\c0.data_in_field_2 ));
    Odrv4 I__6046 (
            .O(N__27202),
            .I(\c0.data_in_field_2 ));
    Odrv12 I__6045 (
            .O(N__27199),
            .I(\c0.data_in_field_2 ));
    Odrv4 I__6044 (
            .O(N__27196),
            .I(\c0.data_in_field_2 ));
    InMux I__6043 (
            .O(N__27187),
            .I(N__27184));
    LocalMux I__6042 (
            .O(N__27184),
            .I(N__27181));
    Span4Mux_v I__6041 (
            .O(N__27181),
            .I(N__27175));
    InMux I__6040 (
            .O(N__27180),
            .I(N__27172));
    InMux I__6039 (
            .O(N__27179),
            .I(N__27169));
    InMux I__6038 (
            .O(N__27178),
            .I(N__27166));
    Span4Mux_h I__6037 (
            .O(N__27175),
            .I(N__27161));
    LocalMux I__6036 (
            .O(N__27172),
            .I(N__27161));
    LocalMux I__6035 (
            .O(N__27169),
            .I(\c0.data_in_field_108 ));
    LocalMux I__6034 (
            .O(N__27166),
            .I(\c0.data_in_field_108 ));
    Odrv4 I__6033 (
            .O(N__27161),
            .I(\c0.data_in_field_108 ));
    InMux I__6032 (
            .O(N__27154),
            .I(N__27151));
    LocalMux I__6031 (
            .O(N__27151),
            .I(N__27147));
    InMux I__6030 (
            .O(N__27150),
            .I(N__27144));
    Odrv12 I__6029 (
            .O(N__27147),
            .I(\c0.n5102 ));
    LocalMux I__6028 (
            .O(N__27144),
            .I(\c0.n5102 ));
    InMux I__6027 (
            .O(N__27139),
            .I(N__27134));
    InMux I__6026 (
            .O(N__27138),
            .I(N__27131));
    InMux I__6025 (
            .O(N__27137),
            .I(N__27127));
    LocalMux I__6024 (
            .O(N__27134),
            .I(N__27123));
    LocalMux I__6023 (
            .O(N__27131),
            .I(N__27120));
    InMux I__6022 (
            .O(N__27130),
            .I(N__27117));
    LocalMux I__6021 (
            .O(N__27127),
            .I(N__27114));
    CascadeMux I__6020 (
            .O(N__27126),
            .I(N__27110));
    Span12Mux_v I__6019 (
            .O(N__27123),
            .I(N__27107));
    Span4Mux_v I__6018 (
            .O(N__27120),
            .I(N__27104));
    LocalMux I__6017 (
            .O(N__27117),
            .I(N__27099));
    Span4Mux_h I__6016 (
            .O(N__27114),
            .I(N__27099));
    InMux I__6015 (
            .O(N__27113),
            .I(N__27094));
    InMux I__6014 (
            .O(N__27110),
            .I(N__27094));
    Odrv12 I__6013 (
            .O(N__27107),
            .I(\c0.data_in_field_142 ));
    Odrv4 I__6012 (
            .O(N__27104),
            .I(\c0.data_in_field_142 ));
    Odrv4 I__6011 (
            .O(N__27099),
            .I(\c0.data_in_field_142 ));
    LocalMux I__6010 (
            .O(N__27094),
            .I(\c0.data_in_field_142 ));
    InMux I__6009 (
            .O(N__27085),
            .I(N__27082));
    LocalMux I__6008 (
            .O(N__27082),
            .I(N__27078));
    CascadeMux I__6007 (
            .O(N__27081),
            .I(N__27075));
    Span12Mux_v I__6006 (
            .O(N__27078),
            .I(N__27072));
    InMux I__6005 (
            .O(N__27075),
            .I(N__27069));
    Odrv12 I__6004 (
            .O(N__27072),
            .I(\c0.n1795 ));
    LocalMux I__6003 (
            .O(N__27069),
            .I(\c0.n1795 ));
    InMux I__6002 (
            .O(N__27064),
            .I(N__27061));
    LocalMux I__6001 (
            .O(N__27061),
            .I(N__27058));
    Odrv12 I__6000 (
            .O(N__27058),
            .I(\c0.n11_adj_1913 ));
    InMux I__5999 (
            .O(N__27055),
            .I(N__27051));
    InMux I__5998 (
            .O(N__27054),
            .I(N__27048));
    LocalMux I__5997 (
            .O(N__27051),
            .I(N__27045));
    LocalMux I__5996 (
            .O(N__27048),
            .I(N__27042));
    Span4Mux_v I__5995 (
            .O(N__27045),
            .I(N__27039));
    Span4Mux_h I__5994 (
            .O(N__27042),
            .I(N__27035));
    Span4Mux_h I__5993 (
            .O(N__27039),
            .I(N__27032));
    InMux I__5992 (
            .O(N__27038),
            .I(N__27029));
    Span4Mux_h I__5991 (
            .O(N__27035),
            .I(N__27026));
    Span4Mux_h I__5990 (
            .O(N__27032),
            .I(N__27023));
    LocalMux I__5989 (
            .O(N__27029),
            .I(data_in_11_4));
    Odrv4 I__5988 (
            .O(N__27026),
            .I(data_in_11_4));
    Odrv4 I__5987 (
            .O(N__27023),
            .I(data_in_11_4));
    InMux I__5986 (
            .O(N__27016),
            .I(N__27013));
    LocalMux I__5985 (
            .O(N__27013),
            .I(N__27009));
    InMux I__5984 (
            .O(N__27012),
            .I(N__27006));
    Span4Mux_h I__5983 (
            .O(N__27009),
            .I(N__27003));
    LocalMux I__5982 (
            .O(N__27006),
            .I(N__27000));
    Span4Mux_v I__5981 (
            .O(N__27003),
            .I(N__26993));
    Span4Mux_v I__5980 (
            .O(N__27000),
            .I(N__26993));
    InMux I__5979 (
            .O(N__26999),
            .I(N__26988));
    InMux I__5978 (
            .O(N__26998),
            .I(N__26988));
    Odrv4 I__5977 (
            .O(N__26993),
            .I(\c0.data_in_field_92 ));
    LocalMux I__5976 (
            .O(N__26988),
            .I(\c0.data_in_field_92 ));
    CascadeMux I__5975 (
            .O(N__26983),
            .I(N__26979));
    InMux I__5974 (
            .O(N__26982),
            .I(N__26975));
    InMux I__5973 (
            .O(N__26979),
            .I(N__26970));
    InMux I__5972 (
            .O(N__26978),
            .I(N__26970));
    LocalMux I__5971 (
            .O(N__26975),
            .I(N__26967));
    LocalMux I__5970 (
            .O(N__26970),
            .I(N__26964));
    Span4Mux_v I__5969 (
            .O(N__26967),
            .I(N__26961));
    Span4Mux_v I__5968 (
            .O(N__26964),
            .I(N__26956));
    Span4Mux_h I__5967 (
            .O(N__26961),
            .I(N__26956));
    Odrv4 I__5966 (
            .O(N__26956),
            .I(data_in_11_5));
    InMux I__5965 (
            .O(N__26953),
            .I(N__26950));
    LocalMux I__5964 (
            .O(N__26950),
            .I(N__26947));
    Span4Mux_v I__5963 (
            .O(N__26947),
            .I(N__26942));
    InMux I__5962 (
            .O(N__26946),
            .I(N__26937));
    InMux I__5961 (
            .O(N__26945),
            .I(N__26937));
    Span4Mux_h I__5960 (
            .O(N__26942),
            .I(N__26931));
    LocalMux I__5959 (
            .O(N__26937),
            .I(N__26931));
    InMux I__5958 (
            .O(N__26936),
            .I(N__26927));
    Span4Mux_h I__5957 (
            .O(N__26931),
            .I(N__26924));
    InMux I__5956 (
            .O(N__26930),
            .I(N__26921));
    LocalMux I__5955 (
            .O(N__26927),
            .I(\c0.data_in_field_93 ));
    Odrv4 I__5954 (
            .O(N__26924),
            .I(\c0.data_in_field_93 ));
    LocalMux I__5953 (
            .O(N__26921),
            .I(\c0.data_in_field_93 ));
    CascadeMux I__5952 (
            .O(N__26914),
            .I(N__26911));
    InMux I__5951 (
            .O(N__26911),
            .I(N__26908));
    LocalMux I__5950 (
            .O(N__26908),
            .I(\c0.n5707 ));
    InMux I__5949 (
            .O(N__26905),
            .I(N__26902));
    LocalMux I__5948 (
            .O(N__26902),
            .I(N__26898));
    InMux I__5947 (
            .O(N__26901),
            .I(N__26895));
    Span4Mux_v I__5946 (
            .O(N__26898),
            .I(N__26891));
    LocalMux I__5945 (
            .O(N__26895),
            .I(N__26888));
    InMux I__5944 (
            .O(N__26894),
            .I(N__26885));
    Odrv4 I__5943 (
            .O(N__26891),
            .I(\c0.n1838 ));
    Odrv12 I__5942 (
            .O(N__26888),
            .I(\c0.n1838 ));
    LocalMux I__5941 (
            .O(N__26885),
            .I(\c0.n1838 ));
    CascadeMux I__5940 (
            .O(N__26878),
            .I(N__26875));
    InMux I__5939 (
            .O(N__26875),
            .I(N__26871));
    InMux I__5938 (
            .O(N__26874),
            .I(N__26868));
    LocalMux I__5937 (
            .O(N__26871),
            .I(N__26865));
    LocalMux I__5936 (
            .O(N__26868),
            .I(N__26862));
    Span4Mux_h I__5935 (
            .O(N__26865),
            .I(N__26858));
    Span4Mux_s3_v I__5934 (
            .O(N__26862),
            .I(N__26855));
    InMux I__5933 (
            .O(N__26861),
            .I(N__26852));
    Odrv4 I__5932 (
            .O(N__26858),
            .I(data_in_5_0));
    Odrv4 I__5931 (
            .O(N__26855),
            .I(data_in_5_0));
    LocalMux I__5930 (
            .O(N__26852),
            .I(data_in_5_0));
    InMux I__5929 (
            .O(N__26845),
            .I(N__26842));
    LocalMux I__5928 (
            .O(N__26842),
            .I(N__26839));
    Span4Mux_v I__5927 (
            .O(N__26839),
            .I(N__26836));
    Span4Mux_h I__5926 (
            .O(N__26836),
            .I(N__26832));
    CascadeMux I__5925 (
            .O(N__26835),
            .I(N__26828));
    Span4Mux_h I__5924 (
            .O(N__26832),
            .I(N__26825));
    InMux I__5923 (
            .O(N__26831),
            .I(N__26822));
    InMux I__5922 (
            .O(N__26828),
            .I(N__26819));
    Span4Mux_h I__5921 (
            .O(N__26825),
            .I(N__26816));
    LocalMux I__5920 (
            .O(N__26822),
            .I(data_in_16_3));
    LocalMux I__5919 (
            .O(N__26819),
            .I(data_in_16_3));
    Odrv4 I__5918 (
            .O(N__26816),
            .I(data_in_16_3));
    CascadeMux I__5917 (
            .O(N__26809),
            .I(N__26804));
    CascadeMux I__5916 (
            .O(N__26808),
            .I(N__26801));
    InMux I__5915 (
            .O(N__26807),
            .I(N__26796));
    InMux I__5914 (
            .O(N__26804),
            .I(N__26796));
    InMux I__5913 (
            .O(N__26801),
            .I(N__26792));
    LocalMux I__5912 (
            .O(N__26796),
            .I(N__26789));
    InMux I__5911 (
            .O(N__26795),
            .I(N__26786));
    LocalMux I__5910 (
            .O(N__26792),
            .I(N__26783));
    Sp12to4 I__5909 (
            .O(N__26789),
            .I(N__26780));
    LocalMux I__5908 (
            .O(N__26786),
            .I(N__26777));
    Span4Mux_h I__5907 (
            .O(N__26783),
            .I(N__26774));
    Span12Mux_v I__5906 (
            .O(N__26780),
            .I(N__26771));
    Odrv4 I__5905 (
            .O(N__26777),
            .I(data_in_18_4));
    Odrv4 I__5904 (
            .O(N__26774),
            .I(data_in_18_4));
    Odrv12 I__5903 (
            .O(N__26771),
            .I(data_in_18_4));
    InMux I__5902 (
            .O(N__26764),
            .I(N__26760));
    CascadeMux I__5901 (
            .O(N__26763),
            .I(N__26756));
    LocalMux I__5900 (
            .O(N__26760),
            .I(N__26753));
    InMux I__5899 (
            .O(N__26759),
            .I(N__26748));
    InMux I__5898 (
            .O(N__26756),
            .I(N__26748));
    Span4Mux_h I__5897 (
            .O(N__26753),
            .I(N__26745));
    LocalMux I__5896 (
            .O(N__26748),
            .I(data_in_17_4));
    Odrv4 I__5895 (
            .O(N__26745),
            .I(data_in_17_4));
    CascadeMux I__5894 (
            .O(N__26740),
            .I(N__26737));
    InMux I__5893 (
            .O(N__26737),
            .I(N__26734));
    LocalMux I__5892 (
            .O(N__26734),
            .I(N__26731));
    Span4Mux_h I__5891 (
            .O(N__26731),
            .I(N__26725));
    InMux I__5890 (
            .O(N__26730),
            .I(N__26722));
    InMux I__5889 (
            .O(N__26729),
            .I(N__26719));
    InMux I__5888 (
            .O(N__26728),
            .I(N__26716));
    Span4Mux_v I__5887 (
            .O(N__26725),
            .I(N__26712));
    LocalMux I__5886 (
            .O(N__26722),
            .I(N__26709));
    LocalMux I__5885 (
            .O(N__26719),
            .I(N__26706));
    LocalMux I__5884 (
            .O(N__26716),
            .I(N__26703));
    InMux I__5883 (
            .O(N__26715),
            .I(N__26699));
    IoSpan4Mux I__5882 (
            .O(N__26712),
            .I(N__26696));
    Span4Mux_h I__5881 (
            .O(N__26709),
            .I(N__26693));
    Span4Mux_v I__5880 (
            .O(N__26706),
            .I(N__26690));
    Span4Mux_h I__5879 (
            .O(N__26703),
            .I(N__26687));
    InMux I__5878 (
            .O(N__26702),
            .I(N__26684));
    LocalMux I__5877 (
            .O(N__26699),
            .I(\c0.data_in_field_63 ));
    Odrv4 I__5876 (
            .O(N__26696),
            .I(\c0.data_in_field_63 ));
    Odrv4 I__5875 (
            .O(N__26693),
            .I(\c0.data_in_field_63 ));
    Odrv4 I__5874 (
            .O(N__26690),
            .I(\c0.data_in_field_63 ));
    Odrv4 I__5873 (
            .O(N__26687),
            .I(\c0.data_in_field_63 ));
    LocalMux I__5872 (
            .O(N__26684),
            .I(\c0.data_in_field_63 ));
    CascadeMux I__5871 (
            .O(N__26671),
            .I(N__26668));
    InMux I__5870 (
            .O(N__26668),
            .I(N__26665));
    LocalMux I__5869 (
            .O(N__26665),
            .I(N__26660));
    InMux I__5868 (
            .O(N__26664),
            .I(N__26657));
    InMux I__5867 (
            .O(N__26663),
            .I(N__26652));
    Span4Mux_h I__5866 (
            .O(N__26660),
            .I(N__26647));
    LocalMux I__5865 (
            .O(N__26657),
            .I(N__26647));
    InMux I__5864 (
            .O(N__26656),
            .I(N__26644));
    InMux I__5863 (
            .O(N__26655),
            .I(N__26641));
    LocalMux I__5862 (
            .O(N__26652),
            .I(\c0.data_in_field_62 ));
    Odrv4 I__5861 (
            .O(N__26647),
            .I(\c0.data_in_field_62 ));
    LocalMux I__5860 (
            .O(N__26644),
            .I(\c0.data_in_field_62 ));
    LocalMux I__5859 (
            .O(N__26641),
            .I(\c0.data_in_field_62 ));
    CascadeMux I__5858 (
            .O(N__26632),
            .I(\c0.n1795_cascade_ ));
    InMux I__5857 (
            .O(N__26629),
            .I(N__26626));
    LocalMux I__5856 (
            .O(N__26626),
            .I(N__26623));
    Odrv12 I__5855 (
            .O(N__26623),
            .I(\c0.n6097 ));
    CascadeMux I__5854 (
            .O(N__26620),
            .I(N__26616));
    InMux I__5853 (
            .O(N__26619),
            .I(N__26613));
    InMux I__5852 (
            .O(N__26616),
            .I(N__26610));
    LocalMux I__5851 (
            .O(N__26613),
            .I(N__26607));
    LocalMux I__5850 (
            .O(N__26610),
            .I(N__26604));
    Span4Mux_h I__5849 (
            .O(N__26607),
            .I(N__26601));
    Span12Mux_h I__5848 (
            .O(N__26604),
            .I(N__26597));
    Span4Mux_v I__5847 (
            .O(N__26601),
            .I(N__26594));
    InMux I__5846 (
            .O(N__26600),
            .I(N__26591));
    Odrv12 I__5845 (
            .O(N__26597),
            .I(data_in_6_3));
    Odrv4 I__5844 (
            .O(N__26594),
            .I(data_in_6_3));
    LocalMux I__5843 (
            .O(N__26591),
            .I(data_in_6_3));
    InMux I__5842 (
            .O(N__26584),
            .I(N__26581));
    LocalMux I__5841 (
            .O(N__26581),
            .I(N__26578));
    Span4Mux_s1_v I__5840 (
            .O(N__26578),
            .I(N__26575));
    Sp12to4 I__5839 (
            .O(N__26575),
            .I(N__26571));
    InMux I__5838 (
            .O(N__26574),
            .I(N__26567));
    Span12Mux_s10_h I__5837 (
            .O(N__26571),
            .I(N__26564));
    InMux I__5836 (
            .O(N__26570),
            .I(N__26561));
    LocalMux I__5835 (
            .O(N__26567),
            .I(data_in_5_3));
    Odrv12 I__5834 (
            .O(N__26564),
            .I(data_in_5_3));
    LocalMux I__5833 (
            .O(N__26561),
            .I(data_in_5_3));
    CascadeMux I__5832 (
            .O(N__26554),
            .I(N__26551));
    InMux I__5831 (
            .O(N__26551),
            .I(N__26548));
    LocalMux I__5830 (
            .O(N__26548),
            .I(N__26545));
    Span4Mux_h I__5829 (
            .O(N__26545),
            .I(N__26542));
    Span4Mux_h I__5828 (
            .O(N__26542),
            .I(N__26539));
    Span4Mux_v I__5827 (
            .O(N__26539),
            .I(N__26534));
    InMux I__5826 (
            .O(N__26538),
            .I(N__26529));
    InMux I__5825 (
            .O(N__26537),
            .I(N__26529));
    Odrv4 I__5824 (
            .O(N__26534),
            .I(data_in_9_1));
    LocalMux I__5823 (
            .O(N__26529),
            .I(data_in_9_1));
    CascadeMux I__5822 (
            .O(N__26524),
            .I(N__26520));
    InMux I__5821 (
            .O(N__26523),
            .I(N__26517));
    InMux I__5820 (
            .O(N__26520),
            .I(N__26514));
    LocalMux I__5819 (
            .O(N__26517),
            .I(N__26511));
    LocalMux I__5818 (
            .O(N__26514),
            .I(N__26505));
    Span4Mux_h I__5817 (
            .O(N__26511),
            .I(N__26505));
    InMux I__5816 (
            .O(N__26510),
            .I(N__26502));
    Odrv4 I__5815 (
            .O(N__26505),
            .I(data_in_7_6));
    LocalMux I__5814 (
            .O(N__26502),
            .I(data_in_7_6));
    CascadeMux I__5813 (
            .O(N__26497),
            .I(N__26493));
    InMux I__5812 (
            .O(N__26496),
            .I(N__26490));
    InMux I__5811 (
            .O(N__26493),
            .I(N__26486));
    LocalMux I__5810 (
            .O(N__26490),
            .I(N__26483));
    InMux I__5809 (
            .O(N__26489),
            .I(N__26480));
    LocalMux I__5808 (
            .O(N__26486),
            .I(data_in_10_4));
    Odrv12 I__5807 (
            .O(N__26483),
            .I(data_in_10_4));
    LocalMux I__5806 (
            .O(N__26480),
            .I(data_in_10_4));
    CascadeMux I__5805 (
            .O(N__26473),
            .I(N__26470));
    InMux I__5804 (
            .O(N__26470),
            .I(N__26467));
    LocalMux I__5803 (
            .O(N__26467),
            .I(N__26464));
    Span4Mux_h I__5802 (
            .O(N__26464),
            .I(N__26461));
    Span4Mux_h I__5801 (
            .O(N__26461),
            .I(N__26458));
    Span4Mux_v I__5800 (
            .O(N__26458),
            .I(N__26453));
    InMux I__5799 (
            .O(N__26457),
            .I(N__26448));
    InMux I__5798 (
            .O(N__26456),
            .I(N__26448));
    Odrv4 I__5797 (
            .O(N__26453),
            .I(data_in_10_3));
    LocalMux I__5796 (
            .O(N__26448),
            .I(data_in_10_3));
    InMux I__5795 (
            .O(N__26443),
            .I(N__26439));
    InMux I__5794 (
            .O(N__26442),
            .I(N__26436));
    LocalMux I__5793 (
            .O(N__26439),
            .I(N__26433));
    LocalMux I__5792 (
            .O(N__26436),
            .I(N__26429));
    Sp12to4 I__5791 (
            .O(N__26433),
            .I(N__26426));
    InMux I__5790 (
            .O(N__26432),
            .I(N__26423));
    Odrv4 I__5789 (
            .O(N__26429),
            .I(data_in_9_3));
    Odrv12 I__5788 (
            .O(N__26426),
            .I(data_in_9_3));
    LocalMux I__5787 (
            .O(N__26423),
            .I(data_in_9_3));
    InMux I__5786 (
            .O(N__26416),
            .I(N__26413));
    LocalMux I__5785 (
            .O(N__26413),
            .I(N__26410));
    Span4Mux_h I__5784 (
            .O(N__26410),
            .I(N__26407));
    Odrv4 I__5783 (
            .O(N__26407),
            .I(\c0.n26_adj_1878 ));
    InMux I__5782 (
            .O(N__26404),
            .I(N__26401));
    LocalMux I__5781 (
            .O(N__26401),
            .I(N__26398));
    Span4Mux_h I__5780 (
            .O(N__26398),
            .I(N__26395));
    Span4Mux_v I__5779 (
            .O(N__26395),
            .I(N__26390));
    InMux I__5778 (
            .O(N__26394),
            .I(N__26385));
    InMux I__5777 (
            .O(N__26393),
            .I(N__26385));
    Odrv4 I__5776 (
            .O(N__26390),
            .I(data_in_0_4));
    LocalMux I__5775 (
            .O(N__26385),
            .I(data_in_0_4));
    InMux I__5774 (
            .O(N__26380),
            .I(N__26376));
    InMux I__5773 (
            .O(N__26379),
            .I(N__26372));
    LocalMux I__5772 (
            .O(N__26376),
            .I(N__26369));
    InMux I__5771 (
            .O(N__26375),
            .I(N__26366));
    LocalMux I__5770 (
            .O(N__26372),
            .I(N__26361));
    Span4Mux_h I__5769 (
            .O(N__26369),
            .I(N__26356));
    LocalMux I__5768 (
            .O(N__26366),
            .I(N__26356));
    InMux I__5767 (
            .O(N__26365),
            .I(N__26352));
    InMux I__5766 (
            .O(N__26364),
            .I(N__26349));
    Span4Mux_v I__5765 (
            .O(N__26361),
            .I(N__26344));
    Span4Mux_v I__5764 (
            .O(N__26356),
            .I(N__26344));
    InMux I__5763 (
            .O(N__26355),
            .I(N__26341));
    LocalMux I__5762 (
            .O(N__26352),
            .I(N__26338));
    LocalMux I__5761 (
            .O(N__26349),
            .I(\c0.data_in_field_68 ));
    Odrv4 I__5760 (
            .O(N__26344),
            .I(\c0.data_in_field_68 ));
    LocalMux I__5759 (
            .O(N__26341),
            .I(\c0.data_in_field_68 ));
    Odrv12 I__5758 (
            .O(N__26338),
            .I(\c0.data_in_field_68 ));
    CascadeMux I__5757 (
            .O(N__26329),
            .I(N__26326));
    InMux I__5756 (
            .O(N__26326),
            .I(N__26322));
    InMux I__5755 (
            .O(N__26325),
            .I(N__26319));
    LocalMux I__5754 (
            .O(N__26322),
            .I(N__26316));
    LocalMux I__5753 (
            .O(N__26319),
            .I(N__26313));
    Span4Mux_h I__5752 (
            .O(N__26316),
            .I(N__26310));
    Span4Mux_h I__5751 (
            .O(N__26313),
            .I(N__26307));
    Odrv4 I__5750 (
            .O(N__26310),
            .I(\c0.n5105 ));
    Odrv4 I__5749 (
            .O(N__26307),
            .I(\c0.n5105 ));
    InMux I__5748 (
            .O(N__26302),
            .I(N__26299));
    LocalMux I__5747 (
            .O(N__26299),
            .I(N__26296));
    Span4Mux_v I__5746 (
            .O(N__26296),
            .I(N__26292));
    InMux I__5745 (
            .O(N__26295),
            .I(N__26289));
    Odrv4 I__5744 (
            .O(N__26292),
            .I(\c0.n5111 ));
    LocalMux I__5743 (
            .O(N__26289),
            .I(\c0.n5111 ));
    InMux I__5742 (
            .O(N__26284),
            .I(N__26281));
    LocalMux I__5741 (
            .O(N__26281),
            .I(N__26278));
    Span12Mux_s10_h I__5740 (
            .O(N__26278),
            .I(N__26275));
    Odrv12 I__5739 (
            .O(N__26275),
            .I(\c0.n35 ));
    CascadeMux I__5738 (
            .O(N__26272),
            .I(N__26268));
    InMux I__5737 (
            .O(N__26271),
            .I(N__26265));
    InMux I__5736 (
            .O(N__26268),
            .I(N__26261));
    LocalMux I__5735 (
            .O(N__26265),
            .I(N__26257));
    InMux I__5734 (
            .O(N__26264),
            .I(N__26254));
    LocalMux I__5733 (
            .O(N__26261),
            .I(N__26251));
    InMux I__5732 (
            .O(N__26260),
            .I(N__26248));
    Span4Mux_v I__5731 (
            .O(N__26257),
            .I(N__26242));
    LocalMux I__5730 (
            .O(N__26254),
            .I(N__26242));
    Span4Mux_h I__5729 (
            .O(N__26251),
            .I(N__26237));
    LocalMux I__5728 (
            .O(N__26248),
            .I(N__26237));
    CascadeMux I__5727 (
            .O(N__26247),
            .I(N__26234));
    Span4Mux_h I__5726 (
            .O(N__26242),
            .I(N__26229));
    Span4Mux_v I__5725 (
            .O(N__26237),
            .I(N__26229));
    InMux I__5724 (
            .O(N__26234),
            .I(N__26226));
    Span4Mux_h I__5723 (
            .O(N__26229),
            .I(N__26223));
    LocalMux I__5722 (
            .O(N__26226),
            .I(\c0.data_in_field_59 ));
    Odrv4 I__5721 (
            .O(N__26223),
            .I(\c0.data_in_field_59 ));
    CascadeMux I__5720 (
            .O(N__26218),
            .I(N__26215));
    InMux I__5719 (
            .O(N__26215),
            .I(N__26211));
    InMux I__5718 (
            .O(N__26214),
            .I(N__26208));
    LocalMux I__5717 (
            .O(N__26211),
            .I(N__26205));
    LocalMux I__5716 (
            .O(N__26208),
            .I(N__26202));
    Span4Mux_v I__5715 (
            .O(N__26205),
            .I(N__26199));
    Span4Mux_s1_v I__5714 (
            .O(N__26202),
            .I(N__26196));
    Span4Mux_h I__5713 (
            .O(N__26199),
            .I(N__26190));
    Span4Mux_v I__5712 (
            .O(N__26196),
            .I(N__26190));
    InMux I__5711 (
            .O(N__26195),
            .I(N__26187));
    Odrv4 I__5710 (
            .O(N__26190),
            .I(data_in_6_6));
    LocalMux I__5709 (
            .O(N__26187),
            .I(data_in_6_6));
    CascadeMux I__5708 (
            .O(N__26182),
            .I(N__26179));
    InMux I__5707 (
            .O(N__26179),
            .I(N__26175));
    InMux I__5706 (
            .O(N__26178),
            .I(N__26172));
    LocalMux I__5705 (
            .O(N__26175),
            .I(N__26167));
    LocalMux I__5704 (
            .O(N__26172),
            .I(N__26167));
    Span12Mux_s10_v I__5703 (
            .O(N__26167),
            .I(N__26163));
    InMux I__5702 (
            .O(N__26166),
            .I(N__26160));
    Odrv12 I__5701 (
            .O(N__26163),
            .I(data_in_13_4));
    LocalMux I__5700 (
            .O(N__26160),
            .I(data_in_13_4));
    InMux I__5699 (
            .O(N__26155),
            .I(N__26151));
    InMux I__5698 (
            .O(N__26154),
            .I(N__26147));
    LocalMux I__5697 (
            .O(N__26151),
            .I(N__26144));
    InMux I__5696 (
            .O(N__26150),
            .I(N__26140));
    LocalMux I__5695 (
            .O(N__26147),
            .I(N__26137));
    Span4Mux_v I__5694 (
            .O(N__26144),
            .I(N__26134));
    InMux I__5693 (
            .O(N__26143),
            .I(N__26131));
    LocalMux I__5692 (
            .O(N__26140),
            .I(N__26128));
    Span12Mux_s8_v I__5691 (
            .O(N__26137),
            .I(N__26125));
    Span4Mux_h I__5690 (
            .O(N__26134),
            .I(N__26118));
    LocalMux I__5689 (
            .O(N__26131),
            .I(N__26118));
    Span4Mux_v I__5688 (
            .O(N__26128),
            .I(N__26118));
    Odrv12 I__5687 (
            .O(N__26125),
            .I(data_in_2_4));
    Odrv4 I__5686 (
            .O(N__26118),
            .I(data_in_2_4));
    CascadeMux I__5685 (
            .O(N__26113),
            .I(N__26108));
    InMux I__5684 (
            .O(N__26112),
            .I(N__26105));
    InMux I__5683 (
            .O(N__26111),
            .I(N__26102));
    InMux I__5682 (
            .O(N__26108),
            .I(N__26098));
    LocalMux I__5681 (
            .O(N__26105),
            .I(N__26095));
    LocalMux I__5680 (
            .O(N__26102),
            .I(N__26092));
    InMux I__5679 (
            .O(N__26101),
            .I(N__26088));
    LocalMux I__5678 (
            .O(N__26098),
            .I(N__26085));
    Span4Mux_v I__5677 (
            .O(N__26095),
            .I(N__26082));
    Span4Mux_h I__5676 (
            .O(N__26092),
            .I(N__26079));
    CascadeMux I__5675 (
            .O(N__26091),
            .I(N__26076));
    LocalMux I__5674 (
            .O(N__26088),
            .I(N__26071));
    Span4Mux_v I__5673 (
            .O(N__26085),
            .I(N__26071));
    Span4Mux_h I__5672 (
            .O(N__26082),
            .I(N__26066));
    Span4Mux_h I__5671 (
            .O(N__26079),
            .I(N__26066));
    InMux I__5670 (
            .O(N__26076),
            .I(N__26063));
    Span4Mux_h I__5669 (
            .O(N__26071),
            .I(N__26060));
    Span4Mux_v I__5668 (
            .O(N__26066),
            .I(N__26057));
    LocalMux I__5667 (
            .O(N__26063),
            .I(\c0.data_in_field_115 ));
    Odrv4 I__5666 (
            .O(N__26060),
            .I(\c0.data_in_field_115 ));
    Odrv4 I__5665 (
            .O(N__26057),
            .I(\c0.data_in_field_115 ));
    InMux I__5664 (
            .O(N__26050),
            .I(N__26047));
    LocalMux I__5663 (
            .O(N__26047),
            .I(N__26044));
    Span4Mux_s2_v I__5662 (
            .O(N__26044),
            .I(N__26040));
    InMux I__5661 (
            .O(N__26043),
            .I(N__26035));
    Span4Mux_h I__5660 (
            .O(N__26040),
            .I(N__26032));
    InMux I__5659 (
            .O(N__26039),
            .I(N__26027));
    InMux I__5658 (
            .O(N__26038),
            .I(N__26027));
    LocalMux I__5657 (
            .O(N__26035),
            .I(data_in_18_7));
    Odrv4 I__5656 (
            .O(N__26032),
            .I(data_in_18_7));
    LocalMux I__5655 (
            .O(N__26027),
            .I(data_in_18_7));
    InMux I__5654 (
            .O(N__26020),
            .I(N__26013));
    InMux I__5653 (
            .O(N__26019),
            .I(N__26013));
    InMux I__5652 (
            .O(N__26018),
            .I(N__26010));
    LocalMux I__5651 (
            .O(N__26013),
            .I(data_in_17_7));
    LocalMux I__5650 (
            .O(N__26010),
            .I(data_in_17_7));
    InMux I__5649 (
            .O(N__26005),
            .I(N__25999));
    InMux I__5648 (
            .O(N__26004),
            .I(N__25999));
    LocalMux I__5647 (
            .O(N__25999),
            .I(N__25994));
    InMux I__5646 (
            .O(N__25998),
            .I(N__25991));
    CascadeMux I__5645 (
            .O(N__25997),
            .I(N__25988));
    Span4Mux_v I__5644 (
            .O(N__25994),
            .I(N__25985));
    LocalMux I__5643 (
            .O(N__25991),
            .I(N__25982));
    InMux I__5642 (
            .O(N__25988),
            .I(N__25978));
    Span4Mux_s2_v I__5641 (
            .O(N__25985),
            .I(N__25975));
    Span12Mux_v I__5640 (
            .O(N__25982),
            .I(N__25972));
    InMux I__5639 (
            .O(N__25981),
            .I(N__25969));
    LocalMux I__5638 (
            .O(N__25978),
            .I(\c0.data_in_field_49 ));
    Odrv4 I__5637 (
            .O(N__25975),
            .I(\c0.data_in_field_49 ));
    Odrv12 I__5636 (
            .O(N__25972),
            .I(\c0.data_in_field_49 ));
    LocalMux I__5635 (
            .O(N__25969),
            .I(\c0.data_in_field_49 ));
    CascadeMux I__5634 (
            .O(N__25960),
            .I(\c0.n2092_cascade_ ));
    InMux I__5633 (
            .O(N__25957),
            .I(N__25953));
    InMux I__5632 (
            .O(N__25956),
            .I(N__25950));
    LocalMux I__5631 (
            .O(N__25953),
            .I(N__25947));
    LocalMux I__5630 (
            .O(N__25950),
            .I(N__25944));
    Odrv4 I__5629 (
            .O(N__25947),
            .I(\c0.n2043 ));
    Odrv12 I__5628 (
            .O(N__25944),
            .I(\c0.n2043 ));
    InMux I__5627 (
            .O(N__25939),
            .I(N__25935));
    InMux I__5626 (
            .O(N__25938),
            .I(N__25932));
    LocalMux I__5625 (
            .O(N__25935),
            .I(N__25929));
    LocalMux I__5624 (
            .O(N__25932),
            .I(N__25926));
    Span4Mux_h I__5623 (
            .O(N__25929),
            .I(N__25923));
    Span4Mux_v I__5622 (
            .O(N__25926),
            .I(N__25920));
    Span4Mux_h I__5621 (
            .O(N__25923),
            .I(N__25917));
    Odrv4 I__5620 (
            .O(N__25920),
            .I(\c0.n5246 ));
    Odrv4 I__5619 (
            .O(N__25917),
            .I(\c0.n5246 ));
    CascadeMux I__5618 (
            .O(N__25912),
            .I(N__25908));
    InMux I__5617 (
            .O(N__25911),
            .I(N__25904));
    InMux I__5616 (
            .O(N__25908),
            .I(N__25901));
    InMux I__5615 (
            .O(N__25907),
            .I(N__25898));
    LocalMux I__5614 (
            .O(N__25904),
            .I(N__25895));
    LocalMux I__5613 (
            .O(N__25901),
            .I(N__25892));
    LocalMux I__5612 (
            .O(N__25898),
            .I(data_in_0_2));
    Odrv4 I__5611 (
            .O(N__25895),
            .I(data_in_0_2));
    Odrv12 I__5610 (
            .O(N__25892),
            .I(data_in_0_2));
    InMux I__5609 (
            .O(N__25885),
            .I(N__25882));
    LocalMux I__5608 (
            .O(N__25882),
            .I(N__25878));
    InMux I__5607 (
            .O(N__25881),
            .I(N__25875));
    Span4Mux_v I__5606 (
            .O(N__25878),
            .I(N__25872));
    LocalMux I__5605 (
            .O(N__25875),
            .I(N__25867));
    Span4Mux_h I__5604 (
            .O(N__25872),
            .I(N__25864));
    InMux I__5603 (
            .O(N__25871),
            .I(N__25859));
    InMux I__5602 (
            .O(N__25870),
            .I(N__25859));
    Odrv4 I__5601 (
            .O(N__25867),
            .I(\c0.data_in_field_9 ));
    Odrv4 I__5600 (
            .O(N__25864),
            .I(\c0.data_in_field_9 ));
    LocalMux I__5599 (
            .O(N__25859),
            .I(\c0.data_in_field_9 ));
    CascadeMux I__5598 (
            .O(N__25852),
            .I(N__25849));
    InMux I__5597 (
            .O(N__25849),
            .I(N__25846));
    LocalMux I__5596 (
            .O(N__25846),
            .I(N__25843));
    Span4Mux_h I__5595 (
            .O(N__25843),
            .I(N__25840));
    Odrv4 I__5594 (
            .O(N__25840),
            .I(\c0.n5749 ));
    InMux I__5593 (
            .O(N__25837),
            .I(N__25832));
    InMux I__5592 (
            .O(N__25836),
            .I(N__25827));
    InMux I__5591 (
            .O(N__25835),
            .I(N__25827));
    LocalMux I__5590 (
            .O(N__25832),
            .I(\c0.data_in_field_1 ));
    LocalMux I__5589 (
            .O(N__25827),
            .I(\c0.data_in_field_1 ));
    InMux I__5588 (
            .O(N__25822),
            .I(N__25819));
    LocalMux I__5587 (
            .O(N__25819),
            .I(N__25816));
    Span12Mux_v I__5586 (
            .O(N__25816),
            .I(N__25813));
    Odrv12 I__5585 (
            .O(N__25813),
            .I(\c0.n5453 ));
    InMux I__5584 (
            .O(N__25810),
            .I(N__25806));
    InMux I__5583 (
            .O(N__25809),
            .I(N__25803));
    LocalMux I__5582 (
            .O(N__25806),
            .I(N__25800));
    LocalMux I__5581 (
            .O(N__25803),
            .I(N__25797));
    Span4Mux_h I__5580 (
            .O(N__25800),
            .I(N__25792));
    Span4Mux_v I__5579 (
            .O(N__25797),
            .I(N__25792));
    Span4Mux_h I__5578 (
            .O(N__25792),
            .I(N__25788));
    InMux I__5577 (
            .O(N__25791),
            .I(N__25785));
    Odrv4 I__5576 (
            .O(N__25788),
            .I(\c0.n1830 ));
    LocalMux I__5575 (
            .O(N__25785),
            .I(\c0.n1830 ));
    InMux I__5574 (
            .O(N__25780),
            .I(N__25777));
    LocalMux I__5573 (
            .O(N__25777),
            .I(\c0.n5141 ));
    InMux I__5572 (
            .O(N__25774),
            .I(N__25771));
    LocalMux I__5571 (
            .O(N__25771),
            .I(N__25767));
    InMux I__5570 (
            .O(N__25770),
            .I(N__25764));
    Span4Mux_h I__5569 (
            .O(N__25767),
            .I(N__25760));
    LocalMux I__5568 (
            .O(N__25764),
            .I(N__25756));
    InMux I__5567 (
            .O(N__25763),
            .I(N__25753));
    Span4Mux_v I__5566 (
            .O(N__25760),
            .I(N__25750));
    InMux I__5565 (
            .O(N__25759),
            .I(N__25746));
    Span4Mux_v I__5564 (
            .O(N__25756),
            .I(N__25741));
    LocalMux I__5563 (
            .O(N__25753),
            .I(N__25741));
    Span4Mux_h I__5562 (
            .O(N__25750),
            .I(N__25738));
    InMux I__5561 (
            .O(N__25749),
            .I(N__25735));
    LocalMux I__5560 (
            .O(N__25746),
            .I(\c0.data_in_field_106 ));
    Odrv4 I__5559 (
            .O(N__25741),
            .I(\c0.data_in_field_106 ));
    Odrv4 I__5558 (
            .O(N__25738),
            .I(\c0.data_in_field_106 ));
    LocalMux I__5557 (
            .O(N__25735),
            .I(\c0.data_in_field_106 ));
    InMux I__5556 (
            .O(N__25726),
            .I(N__25722));
    InMux I__5555 (
            .O(N__25725),
            .I(N__25719));
    LocalMux I__5554 (
            .O(N__25722),
            .I(N__25715));
    LocalMux I__5553 (
            .O(N__25719),
            .I(N__25712));
    InMux I__5552 (
            .O(N__25718),
            .I(N__25709));
    Odrv12 I__5551 (
            .O(N__25715),
            .I(data_in_13_7));
    Odrv4 I__5550 (
            .O(N__25712),
            .I(data_in_13_7));
    LocalMux I__5549 (
            .O(N__25709),
            .I(data_in_13_7));
    InMux I__5548 (
            .O(N__25702),
            .I(N__25699));
    LocalMux I__5547 (
            .O(N__25699),
            .I(N__25696));
    Span4Mux_h I__5546 (
            .O(N__25696),
            .I(N__25693));
    Span4Mux_h I__5545 (
            .O(N__25693),
            .I(N__25688));
    InMux I__5544 (
            .O(N__25692),
            .I(N__25683));
    InMux I__5543 (
            .O(N__25691),
            .I(N__25683));
    Odrv4 I__5542 (
            .O(N__25688),
            .I(\c0.data_in_field_111 ));
    LocalMux I__5541 (
            .O(N__25683),
            .I(\c0.data_in_field_111 ));
    InMux I__5540 (
            .O(N__25678),
            .I(N__25673));
    InMux I__5539 (
            .O(N__25677),
            .I(N__25669));
    InMux I__5538 (
            .O(N__25676),
            .I(N__25665));
    LocalMux I__5537 (
            .O(N__25673),
            .I(N__25662));
    CascadeMux I__5536 (
            .O(N__25672),
            .I(N__25659));
    LocalMux I__5535 (
            .O(N__25669),
            .I(N__25656));
    InMux I__5534 (
            .O(N__25668),
            .I(N__25653));
    LocalMux I__5533 (
            .O(N__25665),
            .I(N__25649));
    Span4Mux_h I__5532 (
            .O(N__25662),
            .I(N__25646));
    InMux I__5531 (
            .O(N__25659),
            .I(N__25643));
    Span12Mux_v I__5530 (
            .O(N__25656),
            .I(N__25640));
    LocalMux I__5529 (
            .O(N__25653),
            .I(N__25637));
    InMux I__5528 (
            .O(N__25652),
            .I(N__25634));
    Span4Mux_h I__5527 (
            .O(N__25649),
            .I(N__25629));
    Span4Mux_v I__5526 (
            .O(N__25646),
            .I(N__25629));
    LocalMux I__5525 (
            .O(N__25643),
            .I(\c0.data_in_field_143 ));
    Odrv12 I__5524 (
            .O(N__25640),
            .I(\c0.data_in_field_143 ));
    Odrv4 I__5523 (
            .O(N__25637),
            .I(\c0.data_in_field_143 ));
    LocalMux I__5522 (
            .O(N__25634),
            .I(\c0.data_in_field_143 ));
    Odrv4 I__5521 (
            .O(N__25629),
            .I(\c0.data_in_field_143 ));
    CascadeMux I__5520 (
            .O(N__25618),
            .I(N__25615));
    InMux I__5519 (
            .O(N__25615),
            .I(N__25612));
    LocalMux I__5518 (
            .O(N__25612),
            .I(N__25609));
    Span4Mux_h I__5517 (
            .O(N__25609),
            .I(N__25605));
    InMux I__5516 (
            .O(N__25608),
            .I(N__25602));
    Span4Mux_s0_v I__5515 (
            .O(N__25605),
            .I(N__25596));
    LocalMux I__5514 (
            .O(N__25602),
            .I(N__25596));
    InMux I__5513 (
            .O(N__25601),
            .I(N__25593));
    Odrv4 I__5512 (
            .O(N__25596),
            .I(data_in_16_7));
    LocalMux I__5511 (
            .O(N__25593),
            .I(data_in_16_7));
    CascadeMux I__5510 (
            .O(N__25588),
            .I(N__25585));
    InMux I__5509 (
            .O(N__25585),
            .I(N__25582));
    LocalMux I__5508 (
            .O(N__25582),
            .I(N__25579));
    Span4Mux_h I__5507 (
            .O(N__25579),
            .I(N__25574));
    InMux I__5506 (
            .O(N__25578),
            .I(N__25569));
    InMux I__5505 (
            .O(N__25577),
            .I(N__25569));
    Odrv4 I__5504 (
            .O(N__25574),
            .I(data_in_4_7));
    LocalMux I__5503 (
            .O(N__25569),
            .I(data_in_4_7));
    InMux I__5502 (
            .O(N__25564),
            .I(N__25561));
    LocalMux I__5501 (
            .O(N__25561),
            .I(N__25557));
    InMux I__5500 (
            .O(N__25560),
            .I(N__25554));
    Span4Mux_v I__5499 (
            .O(N__25557),
            .I(N__25549));
    LocalMux I__5498 (
            .O(N__25554),
            .I(N__25546));
    InMux I__5497 (
            .O(N__25553),
            .I(N__25541));
    InMux I__5496 (
            .O(N__25552),
            .I(N__25541));
    Odrv4 I__5495 (
            .O(N__25549),
            .I(\c0.data_in_field_39 ));
    Odrv4 I__5494 (
            .O(N__25546),
            .I(\c0.data_in_field_39 ));
    LocalMux I__5493 (
            .O(N__25541),
            .I(\c0.data_in_field_39 ));
    InMux I__5492 (
            .O(N__25534),
            .I(N__25530));
    InMux I__5491 (
            .O(N__25533),
            .I(N__25527));
    LocalMux I__5490 (
            .O(N__25530),
            .I(N__25523));
    LocalMux I__5489 (
            .O(N__25527),
            .I(N__25520));
    InMux I__5488 (
            .O(N__25526),
            .I(N__25516));
    Span4Mux_h I__5487 (
            .O(N__25523),
            .I(N__25511));
    Span4Mux_h I__5486 (
            .O(N__25520),
            .I(N__25511));
    InMux I__5485 (
            .O(N__25519),
            .I(N__25508));
    LocalMux I__5484 (
            .O(N__25516),
            .I(\c0.data_in_field_5 ));
    Odrv4 I__5483 (
            .O(N__25511),
            .I(\c0.data_in_field_5 ));
    LocalMux I__5482 (
            .O(N__25508),
            .I(\c0.data_in_field_5 ));
    InMux I__5481 (
            .O(N__25501),
            .I(N__25498));
    LocalMux I__5480 (
            .O(N__25498),
            .I(N__25494));
    CascadeMux I__5479 (
            .O(N__25497),
            .I(N__25488));
    Span4Mux_v I__5478 (
            .O(N__25494),
            .I(N__25485));
    InMux I__5477 (
            .O(N__25493),
            .I(N__25480));
    InMux I__5476 (
            .O(N__25492),
            .I(N__25480));
    CascadeMux I__5475 (
            .O(N__25491),
            .I(N__25477));
    InMux I__5474 (
            .O(N__25488),
            .I(N__25474));
    Span4Mux_h I__5473 (
            .O(N__25485),
            .I(N__25469));
    LocalMux I__5472 (
            .O(N__25480),
            .I(N__25469));
    InMux I__5471 (
            .O(N__25477),
            .I(N__25466));
    LocalMux I__5470 (
            .O(N__25474),
            .I(\c0.data_in_field_79 ));
    Odrv4 I__5469 (
            .O(N__25469),
            .I(\c0.data_in_field_79 ));
    LocalMux I__5468 (
            .O(N__25466),
            .I(\c0.data_in_field_79 ));
    InMux I__5467 (
            .O(N__25459),
            .I(N__25456));
    LocalMux I__5466 (
            .O(N__25456),
            .I(N__25453));
    Span4Mux_s1_h I__5465 (
            .O(N__25453),
            .I(N__25448));
    InMux I__5464 (
            .O(N__25452),
            .I(N__25445));
    CascadeMux I__5463 (
            .O(N__25451),
            .I(N__25442));
    Span4Mux_h I__5462 (
            .O(N__25448),
            .I(N__25439));
    LocalMux I__5461 (
            .O(N__25445),
            .I(N__25436));
    InMux I__5460 (
            .O(N__25442),
            .I(N__25432));
    Span4Mux_h I__5459 (
            .O(N__25439),
            .I(N__25427));
    Span4Mux_h I__5458 (
            .O(N__25436),
            .I(N__25427));
    InMux I__5457 (
            .O(N__25435),
            .I(N__25424));
    LocalMux I__5456 (
            .O(N__25432),
            .I(\c0.data_in_field_77 ));
    Odrv4 I__5455 (
            .O(N__25427),
            .I(\c0.data_in_field_77 ));
    LocalMux I__5454 (
            .O(N__25424),
            .I(\c0.data_in_field_77 ));
    CascadeMux I__5453 (
            .O(N__25417),
            .I(\c0.n10_adj_1871_cascade_ ));
    InMux I__5452 (
            .O(N__25414),
            .I(N__25411));
    LocalMux I__5451 (
            .O(N__25411),
            .I(N__25407));
    InMux I__5450 (
            .O(N__25410),
            .I(N__25404));
    Span4Mux_h I__5449 (
            .O(N__25407),
            .I(N__25399));
    LocalMux I__5448 (
            .O(N__25404),
            .I(N__25399));
    Odrv4 I__5447 (
            .O(N__25399),
            .I(\c0.n5234 ));
    InMux I__5446 (
            .O(N__25396),
            .I(N__25393));
    LocalMux I__5445 (
            .O(N__25393),
            .I(N__25389));
    InMux I__5444 (
            .O(N__25392),
            .I(N__25386));
    Odrv12 I__5443 (
            .O(N__25389),
            .I(\c0.n1975 ));
    LocalMux I__5442 (
            .O(N__25386),
            .I(\c0.n1975 ));
    InMux I__5441 (
            .O(N__25381),
            .I(N__25378));
    LocalMux I__5440 (
            .O(N__25378),
            .I(N__25374));
    InMux I__5439 (
            .O(N__25377),
            .I(N__25371));
    Span4Mux_h I__5438 (
            .O(N__25374),
            .I(N__25368));
    LocalMux I__5437 (
            .O(N__25371),
            .I(N__25362));
    Span4Mux_h I__5436 (
            .O(N__25368),
            .I(N__25359));
    InMux I__5435 (
            .O(N__25367),
            .I(N__25356));
    InMux I__5434 (
            .O(N__25366),
            .I(N__25351));
    InMux I__5433 (
            .O(N__25365),
            .I(N__25351));
    Odrv12 I__5432 (
            .O(N__25362),
            .I(\c0.data_in_field_38 ));
    Odrv4 I__5431 (
            .O(N__25359),
            .I(\c0.data_in_field_38 ));
    LocalMux I__5430 (
            .O(N__25356),
            .I(\c0.data_in_field_38 ));
    LocalMux I__5429 (
            .O(N__25351),
            .I(\c0.data_in_field_38 ));
    InMux I__5428 (
            .O(N__25342),
            .I(N__25339));
    LocalMux I__5427 (
            .O(N__25339),
            .I(N__25336));
    Span4Mux_v I__5426 (
            .O(N__25336),
            .I(N__25333));
    Span4Mux_h I__5425 (
            .O(N__25333),
            .I(N__25328));
    InMux I__5424 (
            .O(N__25332),
            .I(N__25325));
    InMux I__5423 (
            .O(N__25331),
            .I(N__25322));
    Odrv4 I__5422 (
            .O(N__25328),
            .I(data_in_12_1));
    LocalMux I__5421 (
            .O(N__25325),
            .I(data_in_12_1));
    LocalMux I__5420 (
            .O(N__25322),
            .I(data_in_12_1));
    InMux I__5419 (
            .O(N__25315),
            .I(N__25312));
    LocalMux I__5418 (
            .O(N__25312),
            .I(N__25308));
    InMux I__5417 (
            .O(N__25311),
            .I(N__25305));
    Span4Mux_h I__5416 (
            .O(N__25308),
            .I(N__25302));
    LocalMux I__5415 (
            .O(N__25305),
            .I(N__25299));
    Odrv4 I__5414 (
            .O(N__25302),
            .I(\c0.n2062 ));
    Odrv12 I__5413 (
            .O(N__25299),
            .I(\c0.n2062 ));
    CascadeMux I__5412 (
            .O(N__25294),
            .I(N__25289));
    InMux I__5411 (
            .O(N__25293),
            .I(N__25286));
    InMux I__5410 (
            .O(N__25292),
            .I(N__25283));
    InMux I__5409 (
            .O(N__25289),
            .I(N__25279));
    LocalMux I__5408 (
            .O(N__25286),
            .I(N__25276));
    LocalMux I__5407 (
            .O(N__25283),
            .I(N__25273));
    InMux I__5406 (
            .O(N__25282),
            .I(N__25270));
    LocalMux I__5405 (
            .O(N__25279),
            .I(\c0.data_in_field_61 ));
    Odrv4 I__5404 (
            .O(N__25276),
            .I(\c0.data_in_field_61 ));
    Odrv12 I__5403 (
            .O(N__25273),
            .I(\c0.data_in_field_61 ));
    LocalMux I__5402 (
            .O(N__25270),
            .I(\c0.data_in_field_61 ));
    CascadeMux I__5401 (
            .O(N__25261),
            .I(\c0.n5875_cascade_ ));
    InMux I__5400 (
            .O(N__25258),
            .I(N__25255));
    LocalMux I__5399 (
            .O(N__25255),
            .I(N__25252));
    Span4Mux_v I__5398 (
            .O(N__25252),
            .I(N__25246));
    InMux I__5397 (
            .O(N__25251),
            .I(N__25243));
    InMux I__5396 (
            .O(N__25250),
            .I(N__25240));
    InMux I__5395 (
            .O(N__25249),
            .I(N__25237));
    Span4Mux_h I__5394 (
            .O(N__25246),
            .I(N__25234));
    LocalMux I__5393 (
            .O(N__25243),
            .I(N__25231));
    LocalMux I__5392 (
            .O(N__25240),
            .I(N__25228));
    LocalMux I__5391 (
            .O(N__25237),
            .I(\c0.data_in_field_37 ));
    Odrv4 I__5390 (
            .O(N__25234),
            .I(\c0.data_in_field_37 ));
    Odrv12 I__5389 (
            .O(N__25231),
            .I(\c0.data_in_field_37 ));
    Odrv4 I__5388 (
            .O(N__25228),
            .I(\c0.data_in_field_37 ));
    InMux I__5387 (
            .O(N__25219),
            .I(N__25216));
    LocalMux I__5386 (
            .O(N__25216),
            .I(N__25213));
    Span4Mux_h I__5385 (
            .O(N__25213),
            .I(N__25210));
    Sp12to4 I__5384 (
            .O(N__25210),
            .I(N__25207));
    Span12Mux_s4_v I__5383 (
            .O(N__25207),
            .I(N__25204));
    Odrv12 I__5382 (
            .O(N__25204),
            .I(\c0.n5396 ));
    InMux I__5381 (
            .O(N__25201),
            .I(N__25197));
    CascadeMux I__5380 (
            .O(N__25200),
            .I(N__25193));
    LocalMux I__5379 (
            .O(N__25197),
            .I(N__25189));
    CascadeMux I__5378 (
            .O(N__25196),
            .I(N__25186));
    InMux I__5377 (
            .O(N__25193),
            .I(N__25182));
    InMux I__5376 (
            .O(N__25192),
            .I(N__25179));
    Span4Mux_v I__5375 (
            .O(N__25189),
            .I(N__25176));
    InMux I__5374 (
            .O(N__25186),
            .I(N__25171));
    InMux I__5373 (
            .O(N__25185),
            .I(N__25171));
    LocalMux I__5372 (
            .O(N__25182),
            .I(\c0.data_in_field_53 ));
    LocalMux I__5371 (
            .O(N__25179),
            .I(\c0.data_in_field_53 ));
    Odrv4 I__5370 (
            .O(N__25176),
            .I(\c0.data_in_field_53 ));
    LocalMux I__5369 (
            .O(N__25171),
            .I(\c0.data_in_field_53 ));
    InMux I__5368 (
            .O(N__25162),
            .I(N__25157));
    InMux I__5367 (
            .O(N__25161),
            .I(N__25154));
    InMux I__5366 (
            .O(N__25160),
            .I(N__25151));
    LocalMux I__5365 (
            .O(N__25157),
            .I(N__25147));
    LocalMux I__5364 (
            .O(N__25154),
            .I(N__25144));
    LocalMux I__5363 (
            .O(N__25151),
            .I(N__25140));
    InMux I__5362 (
            .O(N__25150),
            .I(N__25137));
    Span4Mux_v I__5361 (
            .O(N__25147),
            .I(N__25132));
    Span4Mux_h I__5360 (
            .O(N__25144),
            .I(N__25132));
    InMux I__5359 (
            .O(N__25143),
            .I(N__25129));
    Span4Mux_h I__5358 (
            .O(N__25140),
            .I(N__25126));
    LocalMux I__5357 (
            .O(N__25137),
            .I(\c0.data_in_field_88 ));
    Odrv4 I__5356 (
            .O(N__25132),
            .I(\c0.data_in_field_88 ));
    LocalMux I__5355 (
            .O(N__25129),
            .I(\c0.data_in_field_88 ));
    Odrv4 I__5354 (
            .O(N__25126),
            .I(\c0.data_in_field_88 ));
    InMux I__5353 (
            .O(N__25117),
            .I(N__25114));
    LocalMux I__5352 (
            .O(N__25114),
            .I(N__25111));
    Span4Mux_v I__5351 (
            .O(N__25111),
            .I(N__25108));
    Span4Mux_h I__5350 (
            .O(N__25108),
            .I(N__25101));
    InMux I__5349 (
            .O(N__25107),
            .I(N__25096));
    InMux I__5348 (
            .O(N__25106),
            .I(N__25096));
    InMux I__5347 (
            .O(N__25105),
            .I(N__25091));
    InMux I__5346 (
            .O(N__25104),
            .I(N__25091));
    Odrv4 I__5345 (
            .O(N__25101),
            .I(\c0.data_in_field_124 ));
    LocalMux I__5344 (
            .O(N__25096),
            .I(\c0.data_in_field_124 ));
    LocalMux I__5343 (
            .O(N__25091),
            .I(\c0.data_in_field_124 ));
    InMux I__5342 (
            .O(N__25084),
            .I(N__25081));
    LocalMux I__5341 (
            .O(N__25081),
            .I(N__25077));
    CascadeMux I__5340 (
            .O(N__25080),
            .I(N__25074));
    Span4Mux_h I__5339 (
            .O(N__25077),
            .I(N__25071));
    InMux I__5338 (
            .O(N__25074),
            .I(N__25068));
    Odrv4 I__5337 (
            .O(N__25071),
            .I(\c0.n1944 ));
    LocalMux I__5336 (
            .O(N__25068),
            .I(\c0.n1944 ));
    CascadeMux I__5335 (
            .O(N__25063),
            .I(\c0.n1944_cascade_ ));
    CascadeMux I__5334 (
            .O(N__25060),
            .I(\c0.n20_cascade_ ));
    InMux I__5333 (
            .O(N__25057),
            .I(N__25053));
    InMux I__5332 (
            .O(N__25056),
            .I(N__25049));
    LocalMux I__5331 (
            .O(N__25053),
            .I(N__25046));
    InMux I__5330 (
            .O(N__25052),
            .I(N__25043));
    LocalMux I__5329 (
            .O(N__25049),
            .I(N__25040));
    Span12Mux_s2_h I__5328 (
            .O(N__25046),
            .I(N__25033));
    LocalMux I__5327 (
            .O(N__25043),
            .I(N__25033));
    Span4Mux_v I__5326 (
            .O(N__25040),
            .I(N__25030));
    InMux I__5325 (
            .O(N__25039),
            .I(N__25025));
    InMux I__5324 (
            .O(N__25038),
            .I(N__25025));
    Odrv12 I__5323 (
            .O(N__25033),
            .I(\c0.data_in_field_43 ));
    Odrv4 I__5322 (
            .O(N__25030),
            .I(\c0.data_in_field_43 ));
    LocalMux I__5321 (
            .O(N__25025),
            .I(\c0.data_in_field_43 ));
    InMux I__5320 (
            .O(N__25018),
            .I(N__25015));
    LocalMux I__5319 (
            .O(N__25015),
            .I(N__25012));
    Odrv12 I__5318 (
            .O(N__25012),
            .I(\c0.n24 ));
    InMux I__5317 (
            .O(N__25009),
            .I(N__25005));
    CascadeMux I__5316 (
            .O(N__25008),
            .I(N__25000));
    LocalMux I__5315 (
            .O(N__25005),
            .I(N__24997));
    InMux I__5314 (
            .O(N__25004),
            .I(N__24994));
    InMux I__5313 (
            .O(N__25003),
            .I(N__24991));
    InMux I__5312 (
            .O(N__25000),
            .I(N__24988));
    Span4Mux_h I__5311 (
            .O(N__24997),
            .I(N__24983));
    LocalMux I__5310 (
            .O(N__24994),
            .I(N__24983));
    LocalMux I__5309 (
            .O(N__24991),
            .I(N__24980));
    LocalMux I__5308 (
            .O(N__24988),
            .I(\c0.data_in_field_139 ));
    Odrv4 I__5307 (
            .O(N__24983),
            .I(\c0.data_in_field_139 ));
    Odrv12 I__5306 (
            .O(N__24980),
            .I(\c0.data_in_field_139 ));
    CascadeMux I__5305 (
            .O(N__24973),
            .I(\c0.n1947_cascade_ ));
    InMux I__5304 (
            .O(N__24970),
            .I(N__24967));
    LocalMux I__5303 (
            .O(N__24967),
            .I(\c0.n10 ));
    CascadeMux I__5302 (
            .O(N__24964),
            .I(N__24961));
    InMux I__5301 (
            .O(N__24961),
            .I(N__24957));
    CascadeMux I__5300 (
            .O(N__24960),
            .I(N__24953));
    LocalMux I__5299 (
            .O(N__24957),
            .I(N__24950));
    InMux I__5298 (
            .O(N__24956),
            .I(N__24947));
    InMux I__5297 (
            .O(N__24953),
            .I(N__24944));
    Span4Mux_v I__5296 (
            .O(N__24950),
            .I(N__24939));
    LocalMux I__5295 (
            .O(N__24947),
            .I(N__24939));
    LocalMux I__5294 (
            .O(N__24944),
            .I(N__24936));
    Span4Mux_h I__5293 (
            .O(N__24939),
            .I(N__24933));
    Span12Mux_s9_h I__5292 (
            .O(N__24936),
            .I(N__24928));
    Span4Mux_h I__5291 (
            .O(N__24933),
            .I(N__24925));
    InMux I__5290 (
            .O(N__24932),
            .I(N__24920));
    InMux I__5289 (
            .O(N__24931),
            .I(N__24920));
    Odrv12 I__5288 (
            .O(N__24928),
            .I(\c0.data_in_field_51 ));
    Odrv4 I__5287 (
            .O(N__24925),
            .I(\c0.data_in_field_51 ));
    LocalMux I__5286 (
            .O(N__24920),
            .I(\c0.data_in_field_51 ));
    InMux I__5285 (
            .O(N__24913),
            .I(N__24910));
    LocalMux I__5284 (
            .O(N__24910),
            .I(N__24906));
    InMux I__5283 (
            .O(N__24909),
            .I(N__24903));
    Odrv12 I__5282 (
            .O(N__24906),
            .I(\c0.n1922 ));
    LocalMux I__5281 (
            .O(N__24903),
            .I(\c0.n1922 ));
    InMux I__5280 (
            .O(N__24898),
            .I(N__24895));
    LocalMux I__5279 (
            .O(N__24895),
            .I(N__24891));
    InMux I__5278 (
            .O(N__24894),
            .I(N__24888));
    Span4Mux_h I__5277 (
            .O(N__24891),
            .I(N__24880));
    LocalMux I__5276 (
            .O(N__24888),
            .I(N__24880));
    InMux I__5275 (
            .O(N__24887),
            .I(N__24877));
    InMux I__5274 (
            .O(N__24886),
            .I(N__24872));
    InMux I__5273 (
            .O(N__24885),
            .I(N__24872));
    Odrv4 I__5272 (
            .O(N__24880),
            .I(\c0.data_in_field_75 ));
    LocalMux I__5271 (
            .O(N__24877),
            .I(\c0.data_in_field_75 ));
    LocalMux I__5270 (
            .O(N__24872),
            .I(\c0.data_in_field_75 ));
    InMux I__5269 (
            .O(N__24865),
            .I(N__24862));
    LocalMux I__5268 (
            .O(N__24862),
            .I(N__24859));
    Span4Mux_h I__5267 (
            .O(N__24859),
            .I(N__24856));
    Odrv4 I__5266 (
            .O(N__24856),
            .I(\c0.n5474 ));
    InMux I__5265 (
            .O(N__24853),
            .I(N__24850));
    LocalMux I__5264 (
            .O(N__24850),
            .I(N__24847));
    Span12Mux_s9_h I__5263 (
            .O(N__24847),
            .I(N__24844));
    Odrv12 I__5262 (
            .O(N__24844),
            .I(\c0.n26_adj_1884 ));
    InMux I__5261 (
            .O(N__24841),
            .I(N__24837));
    InMux I__5260 (
            .O(N__24840),
            .I(N__24833));
    LocalMux I__5259 (
            .O(N__24837),
            .I(N__24830));
    CascadeMux I__5258 (
            .O(N__24836),
            .I(N__24825));
    LocalMux I__5257 (
            .O(N__24833),
            .I(N__24822));
    Span4Mux_h I__5256 (
            .O(N__24830),
            .I(N__24819));
    InMux I__5255 (
            .O(N__24829),
            .I(N__24816));
    InMux I__5254 (
            .O(N__24828),
            .I(N__24813));
    InMux I__5253 (
            .O(N__24825),
            .I(N__24810));
    Span4Mux_v I__5252 (
            .O(N__24822),
            .I(N__24805));
    Span4Mux_h I__5251 (
            .O(N__24819),
            .I(N__24805));
    LocalMux I__5250 (
            .O(N__24816),
            .I(N__24802));
    LocalMux I__5249 (
            .O(N__24813),
            .I(\c0.data_in_field_98 ));
    LocalMux I__5248 (
            .O(N__24810),
            .I(\c0.data_in_field_98 ));
    Odrv4 I__5247 (
            .O(N__24805),
            .I(\c0.data_in_field_98 ));
    Odrv4 I__5246 (
            .O(N__24802),
            .I(\c0.data_in_field_98 ));
    CascadeMux I__5245 (
            .O(N__24793),
            .I(N__24790));
    InMux I__5244 (
            .O(N__24790),
            .I(N__24786));
    InMux I__5243 (
            .O(N__24789),
            .I(N__24783));
    LocalMux I__5242 (
            .O(N__24786),
            .I(N__24780));
    LocalMux I__5241 (
            .O(N__24783),
            .I(N__24776));
    Span4Mux_v I__5240 (
            .O(N__24780),
            .I(N__24773));
    InMux I__5239 (
            .O(N__24779),
            .I(N__24770));
    Span4Mux_v I__5238 (
            .O(N__24776),
            .I(N__24767));
    Span4Mux_h I__5237 (
            .O(N__24773),
            .I(N__24764));
    LocalMux I__5236 (
            .O(N__24770),
            .I(data_in_12_7));
    Odrv4 I__5235 (
            .O(N__24767),
            .I(data_in_12_7));
    Odrv4 I__5234 (
            .O(N__24764),
            .I(data_in_12_7));
    CascadeMux I__5233 (
            .O(N__24757),
            .I(N__24753));
    InMux I__5232 (
            .O(N__24756),
            .I(N__24750));
    InMux I__5231 (
            .O(N__24753),
            .I(N__24747));
    LocalMux I__5230 (
            .O(N__24750),
            .I(N__24744));
    LocalMux I__5229 (
            .O(N__24747),
            .I(N__24741));
    Span4Mux_v I__5228 (
            .O(N__24744),
            .I(N__24736));
    Span4Mux_v I__5227 (
            .O(N__24741),
            .I(N__24733));
    CascadeMux I__5226 (
            .O(N__24740),
            .I(N__24730));
    InMux I__5225 (
            .O(N__24739),
            .I(N__24727));
    Span4Mux_h I__5224 (
            .O(N__24736),
            .I(N__24724));
    Sp12to4 I__5223 (
            .O(N__24733),
            .I(N__24721));
    InMux I__5222 (
            .O(N__24730),
            .I(N__24718));
    LocalMux I__5221 (
            .O(N__24727),
            .I(\c0.data_in_field_103 ));
    Odrv4 I__5220 (
            .O(N__24724),
            .I(\c0.data_in_field_103 ));
    Odrv12 I__5219 (
            .O(N__24721),
            .I(\c0.data_in_field_103 ));
    LocalMux I__5218 (
            .O(N__24718),
            .I(\c0.data_in_field_103 ));
    InMux I__5217 (
            .O(N__24709),
            .I(N__24706));
    LocalMux I__5216 (
            .O(N__24706),
            .I(N__24703));
    Span4Mux_v I__5215 (
            .O(N__24703),
            .I(N__24700));
    Span4Mux_h I__5214 (
            .O(N__24700),
            .I(N__24694));
    InMux I__5213 (
            .O(N__24699),
            .I(N__24687));
    InMux I__5212 (
            .O(N__24698),
            .I(N__24687));
    InMux I__5211 (
            .O(N__24697),
            .I(N__24687));
    Odrv4 I__5210 (
            .O(N__24694),
            .I(\c0.data_in_field_28 ));
    LocalMux I__5209 (
            .O(N__24687),
            .I(\c0.data_in_field_28 ));
    InMux I__5208 (
            .O(N__24682),
            .I(N__24679));
    LocalMux I__5207 (
            .O(N__24679),
            .I(N__24676));
    Span4Mux_h I__5206 (
            .O(N__24676),
            .I(N__24672));
    InMux I__5205 (
            .O(N__24675),
            .I(N__24669));
    Span4Mux_v I__5204 (
            .O(N__24672),
            .I(N__24665));
    LocalMux I__5203 (
            .O(N__24669),
            .I(N__24662));
    InMux I__5202 (
            .O(N__24668),
            .I(N__24658));
    Span4Mux_h I__5201 (
            .O(N__24665),
            .I(N__24655));
    Span4Mux_v I__5200 (
            .O(N__24662),
            .I(N__24652));
    InMux I__5199 (
            .O(N__24661),
            .I(N__24649));
    LocalMux I__5198 (
            .O(N__24658),
            .I(\c0.data_in_field_20 ));
    Odrv4 I__5197 (
            .O(N__24655),
            .I(\c0.data_in_field_20 ));
    Odrv4 I__5196 (
            .O(N__24652),
            .I(\c0.data_in_field_20 ));
    LocalMux I__5195 (
            .O(N__24649),
            .I(\c0.data_in_field_20 ));
    InMux I__5194 (
            .O(N__24640),
            .I(N__24636));
    InMux I__5193 (
            .O(N__24639),
            .I(N__24632));
    LocalMux I__5192 (
            .O(N__24636),
            .I(N__24629));
    InMux I__5191 (
            .O(N__24635),
            .I(N__24626));
    LocalMux I__5190 (
            .O(N__24632),
            .I(N__24623));
    Span4Mux_v I__5189 (
            .O(N__24629),
            .I(N__24618));
    LocalMux I__5188 (
            .O(N__24626),
            .I(N__24618));
    Span4Mux_v I__5187 (
            .O(N__24623),
            .I(N__24613));
    Span4Mux_h I__5186 (
            .O(N__24618),
            .I(N__24610));
    InMux I__5185 (
            .O(N__24617),
            .I(N__24605));
    InMux I__5184 (
            .O(N__24616),
            .I(N__24605));
    Odrv4 I__5183 (
            .O(N__24613),
            .I(\c0.data_in_field_12 ));
    Odrv4 I__5182 (
            .O(N__24610),
            .I(\c0.data_in_field_12 ));
    LocalMux I__5181 (
            .O(N__24605),
            .I(\c0.data_in_field_12 ));
    CascadeMux I__5180 (
            .O(N__24598),
            .I(\c0.n5851_cascade_ ));
    CascadeMux I__5179 (
            .O(N__24595),
            .I(N__24592));
    InMux I__5178 (
            .O(N__24592),
            .I(N__24589));
    LocalMux I__5177 (
            .O(N__24589),
            .I(N__24586));
    Span4Mux_h I__5176 (
            .O(N__24586),
            .I(N__24583));
    Odrv4 I__5175 (
            .O(N__24583),
            .I(\c0.n5408 ));
    InMux I__5174 (
            .O(N__24580),
            .I(N__24576));
    InMux I__5173 (
            .O(N__24579),
            .I(N__24573));
    LocalMux I__5172 (
            .O(N__24576),
            .I(N__24570));
    LocalMux I__5171 (
            .O(N__24573),
            .I(N__24567));
    Span4Mux_h I__5170 (
            .O(N__24570),
            .I(N__24564));
    Span4Mux_h I__5169 (
            .O(N__24567),
            .I(N__24561));
    Span4Mux_h I__5168 (
            .O(N__24564),
            .I(N__24558));
    Span4Mux_v I__5167 (
            .O(N__24561),
            .I(N__24555));
    Odrv4 I__5166 (
            .O(N__24558),
            .I(\c0.n5267 ));
    Odrv4 I__5165 (
            .O(N__24555),
            .I(\c0.n5267 ));
    CascadeMux I__5164 (
            .O(N__24550),
            .I(N__24547));
    InMux I__5163 (
            .O(N__24547),
            .I(N__24544));
    LocalMux I__5162 (
            .O(N__24544),
            .I(N__24541));
    Span4Mux_h I__5161 (
            .O(N__24541),
            .I(N__24538));
    Odrv4 I__5160 (
            .O(N__24538),
            .I(\c0.n5905 ));
    InMux I__5159 (
            .O(N__24535),
            .I(N__24532));
    LocalMux I__5158 (
            .O(N__24532),
            .I(\c0.n2074 ));
    CascadeMux I__5157 (
            .O(N__24529),
            .I(N__24525));
    InMux I__5156 (
            .O(N__24528),
            .I(N__24521));
    InMux I__5155 (
            .O(N__24525),
            .I(N__24518));
    CascadeMux I__5154 (
            .O(N__24524),
            .I(N__24515));
    LocalMux I__5153 (
            .O(N__24521),
            .I(N__24512));
    LocalMux I__5152 (
            .O(N__24518),
            .I(N__24509));
    InMux I__5151 (
            .O(N__24515),
            .I(N__24506));
    Span4Mux_v I__5150 (
            .O(N__24512),
            .I(N__24500));
    Span4Mux_v I__5149 (
            .O(N__24509),
            .I(N__24500));
    LocalMux I__5148 (
            .O(N__24506),
            .I(N__24497));
    InMux I__5147 (
            .O(N__24505),
            .I(N__24494));
    Sp12to4 I__5146 (
            .O(N__24500),
            .I(N__24489));
    Span12Mux_h I__5145 (
            .O(N__24497),
            .I(N__24489));
    LocalMux I__5144 (
            .O(N__24494),
            .I(data_in_19_5));
    Odrv12 I__5143 (
            .O(N__24489),
            .I(data_in_19_5));
    InMux I__5142 (
            .O(N__24484),
            .I(N__24481));
    LocalMux I__5141 (
            .O(N__24481),
            .I(N__24478));
    Odrv12 I__5140 (
            .O(N__24478),
            .I(\c0.n22_adj_1914 ));
    InMux I__5139 (
            .O(N__24475),
            .I(N__24471));
    InMux I__5138 (
            .O(N__24474),
            .I(N__24468));
    LocalMux I__5137 (
            .O(N__24471),
            .I(N__24465));
    LocalMux I__5136 (
            .O(N__24468),
            .I(N__24462));
    Span4Mux_h I__5135 (
            .O(N__24465),
            .I(N__24458));
    Span4Mux_s2_v I__5134 (
            .O(N__24462),
            .I(N__24455));
    InMux I__5133 (
            .O(N__24461),
            .I(N__24452));
    Span4Mux_h I__5132 (
            .O(N__24458),
            .I(N__24447));
    Span4Mux_h I__5131 (
            .O(N__24455),
            .I(N__24447));
    LocalMux I__5130 (
            .O(N__24452),
            .I(data_in_16_5));
    Odrv4 I__5129 (
            .O(N__24447),
            .I(data_in_16_5));
    CascadeMux I__5128 (
            .O(N__24442),
            .I(N__24439));
    InMux I__5127 (
            .O(N__24439),
            .I(N__24436));
    LocalMux I__5126 (
            .O(N__24436),
            .I(N__24431));
    InMux I__5125 (
            .O(N__24435),
            .I(N__24428));
    CascadeMux I__5124 (
            .O(N__24434),
            .I(N__24425));
    Span4Mux_h I__5123 (
            .O(N__24431),
            .I(N__24420));
    LocalMux I__5122 (
            .O(N__24428),
            .I(N__24420));
    InMux I__5121 (
            .O(N__24425),
            .I(N__24417));
    Span4Mux_h I__5120 (
            .O(N__24420),
            .I(N__24413));
    LocalMux I__5119 (
            .O(N__24417),
            .I(N__24410));
    InMux I__5118 (
            .O(N__24416),
            .I(N__24407));
    Span4Mux_v I__5117 (
            .O(N__24413),
            .I(N__24404));
    Span12Mux_s5_h I__5116 (
            .O(N__24410),
            .I(N__24401));
    LocalMux I__5115 (
            .O(N__24407),
            .I(data_in_19_2));
    Odrv4 I__5114 (
            .O(N__24404),
            .I(data_in_19_2));
    Odrv12 I__5113 (
            .O(N__24401),
            .I(data_in_19_2));
    CascadeMux I__5112 (
            .O(N__24394),
            .I(N__24391));
    InMux I__5111 (
            .O(N__24391),
            .I(N__24388));
    LocalMux I__5110 (
            .O(N__24388),
            .I(N__24385));
    Odrv4 I__5109 (
            .O(N__24385),
            .I(\c0.n5779 ));
    InMux I__5108 (
            .O(N__24382),
            .I(N__24376));
    InMux I__5107 (
            .O(N__24381),
            .I(N__24376));
    LocalMux I__5106 (
            .O(N__24376),
            .I(N__24372));
    InMux I__5105 (
            .O(N__24375),
            .I(N__24369));
    Odrv4 I__5104 (
            .O(N__24372),
            .I(data_in_13_0));
    LocalMux I__5103 (
            .O(N__24369),
            .I(data_in_13_0));
    InMux I__5102 (
            .O(N__24364),
            .I(N__24358));
    InMux I__5101 (
            .O(N__24363),
            .I(N__24358));
    LocalMux I__5100 (
            .O(N__24358),
            .I(N__24355));
    Span4Mux_h I__5099 (
            .O(N__24355),
            .I(N__24352));
    Span4Mux_h I__5098 (
            .O(N__24352),
            .I(N__24348));
    InMux I__5097 (
            .O(N__24351),
            .I(N__24345));
    Odrv4 I__5096 (
            .O(N__24348),
            .I(data_in_14_0));
    LocalMux I__5095 (
            .O(N__24345),
            .I(data_in_14_0));
    InMux I__5094 (
            .O(N__24340),
            .I(N__24337));
    LocalMux I__5093 (
            .O(N__24337),
            .I(N__24334));
    Span4Mux_h I__5092 (
            .O(N__24334),
            .I(N__24331));
    Odrv4 I__5091 (
            .O(N__24331),
            .I(\c0.n1929 ));
    InMux I__5090 (
            .O(N__24328),
            .I(N__24324));
    CascadeMux I__5089 (
            .O(N__24327),
            .I(N__24320));
    LocalMux I__5088 (
            .O(N__24324),
            .I(N__24317));
    CascadeMux I__5087 (
            .O(N__24323),
            .I(N__24313));
    InMux I__5086 (
            .O(N__24320),
            .I(N__24310));
    Span4Mux_v I__5085 (
            .O(N__24317),
            .I(N__24307));
    InMux I__5084 (
            .O(N__24316),
            .I(N__24304));
    InMux I__5083 (
            .O(N__24313),
            .I(N__24301));
    LocalMux I__5082 (
            .O(N__24310),
            .I(N__24298));
    Span4Mux_h I__5081 (
            .O(N__24307),
            .I(N__24293));
    LocalMux I__5080 (
            .O(N__24304),
            .I(N__24293));
    LocalMux I__5079 (
            .O(N__24301),
            .I(\c0.data_in_field_112 ));
    Odrv4 I__5078 (
            .O(N__24298),
            .I(\c0.data_in_field_112 ));
    Odrv4 I__5077 (
            .O(N__24293),
            .I(\c0.data_in_field_112 ));
    CascadeMux I__5076 (
            .O(N__24286),
            .I(\c0.n1929_cascade_ ));
    CascadeMux I__5075 (
            .O(N__24283),
            .I(\c0.n10_adj_1870_cascade_ ));
    InMux I__5074 (
            .O(N__24280),
            .I(N__24276));
    CascadeMux I__5073 (
            .O(N__24279),
            .I(N__24273));
    LocalMux I__5072 (
            .O(N__24276),
            .I(N__24270));
    InMux I__5071 (
            .O(N__24273),
            .I(N__24267));
    Span4Mux_v I__5070 (
            .O(N__24270),
            .I(N__24264));
    LocalMux I__5069 (
            .O(N__24267),
            .I(N__24261));
    Span4Mux_h I__5068 (
            .O(N__24264),
            .I(N__24258));
    Span4Mux_v I__5067 (
            .O(N__24261),
            .I(N__24255));
    Odrv4 I__5066 (
            .O(N__24258),
            .I(\c0.n5204 ));
    Odrv4 I__5065 (
            .O(N__24255),
            .I(\c0.n5204 ));
    InMux I__5064 (
            .O(N__24250),
            .I(N__24247));
    LocalMux I__5063 (
            .O(N__24247),
            .I(N__24243));
    InMux I__5062 (
            .O(N__24246),
            .I(N__24240));
    Span4Mux_s2_v I__5061 (
            .O(N__24243),
            .I(N__24235));
    LocalMux I__5060 (
            .O(N__24240),
            .I(N__24235));
    Span4Mux_h I__5059 (
            .O(N__24235),
            .I(N__24231));
    InMux I__5058 (
            .O(N__24234),
            .I(N__24228));
    Odrv4 I__5057 (
            .O(N__24231),
            .I(data_in_7_5));
    LocalMux I__5056 (
            .O(N__24228),
            .I(data_in_7_5));
    CascadeMux I__5055 (
            .O(N__24223),
            .I(N__24219));
    InMux I__5054 (
            .O(N__24222),
            .I(N__24216));
    InMux I__5053 (
            .O(N__24219),
            .I(N__24213));
    LocalMux I__5052 (
            .O(N__24216),
            .I(N__24208));
    LocalMux I__5051 (
            .O(N__24213),
            .I(N__24205));
    InMux I__5050 (
            .O(N__24212),
            .I(N__24202));
    InMux I__5049 (
            .O(N__24211),
            .I(N__24199));
    Span12Mux_s2_v I__5048 (
            .O(N__24208),
            .I(N__24196));
    Span4Mux_v I__5047 (
            .O(N__24205),
            .I(N__24193));
    LocalMux I__5046 (
            .O(N__24202),
            .I(data_in_18_6));
    LocalMux I__5045 (
            .O(N__24199),
            .I(data_in_18_6));
    Odrv12 I__5044 (
            .O(N__24196),
            .I(data_in_18_6));
    Odrv4 I__5043 (
            .O(N__24193),
            .I(data_in_18_6));
    CascadeMux I__5042 (
            .O(N__24184),
            .I(N__24180));
    InMux I__5041 (
            .O(N__24183),
            .I(N__24177));
    InMux I__5040 (
            .O(N__24180),
            .I(N__24174));
    LocalMux I__5039 (
            .O(N__24177),
            .I(N__24171));
    LocalMux I__5038 (
            .O(N__24174),
            .I(N__24167));
    Span4Mux_h I__5037 (
            .O(N__24171),
            .I(N__24164));
    InMux I__5036 (
            .O(N__24170),
            .I(N__24161));
    Odrv4 I__5035 (
            .O(N__24167),
            .I(data_in_17_6));
    Odrv4 I__5034 (
            .O(N__24164),
            .I(data_in_17_6));
    LocalMux I__5033 (
            .O(N__24161),
            .I(data_in_17_6));
    InMux I__5032 (
            .O(N__24154),
            .I(N__24151));
    LocalMux I__5031 (
            .O(N__24151),
            .I(N__24147));
    InMux I__5030 (
            .O(N__24150),
            .I(N__24143));
    Span4Mux_v I__5029 (
            .O(N__24147),
            .I(N__24140));
    InMux I__5028 (
            .O(N__24146),
            .I(N__24136));
    LocalMux I__5027 (
            .O(N__24143),
            .I(N__24133));
    Sp12to4 I__5026 (
            .O(N__24140),
            .I(N__24130));
    InMux I__5025 (
            .O(N__24139),
            .I(N__24127));
    LocalMux I__5024 (
            .O(N__24136),
            .I(data_in_1_5));
    Odrv12 I__5023 (
            .O(N__24133),
            .I(data_in_1_5));
    Odrv12 I__5022 (
            .O(N__24130),
            .I(data_in_1_5));
    LocalMux I__5021 (
            .O(N__24127),
            .I(data_in_1_5));
    CascadeMux I__5020 (
            .O(N__24118),
            .I(N__24115));
    InMux I__5019 (
            .O(N__24115),
            .I(N__24111));
    InMux I__5018 (
            .O(N__24114),
            .I(N__24108));
    LocalMux I__5017 (
            .O(N__24111),
            .I(N__24105));
    LocalMux I__5016 (
            .O(N__24108),
            .I(N__24102));
    Span4Mux_v I__5015 (
            .O(N__24105),
            .I(N__24098));
    Span4Mux_h I__5014 (
            .O(N__24102),
            .I(N__24095));
    InMux I__5013 (
            .O(N__24101),
            .I(N__24092));
    Odrv4 I__5012 (
            .O(N__24098),
            .I(data_in_7_7));
    Odrv4 I__5011 (
            .O(N__24095),
            .I(data_in_7_7));
    LocalMux I__5010 (
            .O(N__24092),
            .I(data_in_7_7));
    InMux I__5009 (
            .O(N__24085),
            .I(N__24082));
    LocalMux I__5008 (
            .O(N__24082),
            .I(N__24078));
    InMux I__5007 (
            .O(N__24081),
            .I(N__24075));
    Span4Mux_v I__5006 (
            .O(N__24078),
            .I(N__24072));
    LocalMux I__5005 (
            .O(N__24075),
            .I(N__24069));
    Sp12to4 I__5004 (
            .O(N__24072),
            .I(N__24062));
    Span12Mux_v I__5003 (
            .O(N__24069),
            .I(N__24062));
    InMux I__5002 (
            .O(N__24068),
            .I(N__24057));
    InMux I__5001 (
            .O(N__24067),
            .I(N__24057));
    Odrv12 I__5000 (
            .O(N__24062),
            .I(\c0.data_in_field_121 ));
    LocalMux I__4999 (
            .O(N__24057),
            .I(\c0.data_in_field_121 ));
    InMux I__4998 (
            .O(N__24052),
            .I(N__24049));
    LocalMux I__4997 (
            .O(N__24049),
            .I(N__24044));
    InMux I__4996 (
            .O(N__24048),
            .I(N__24040));
    InMux I__4995 (
            .O(N__24047),
            .I(N__24037));
    Span4Mux_h I__4994 (
            .O(N__24044),
            .I(N__24034));
    InMux I__4993 (
            .O(N__24043),
            .I(N__24031));
    LocalMux I__4992 (
            .O(N__24040),
            .I(N__24026));
    LocalMux I__4991 (
            .O(N__24037),
            .I(N__24026));
    Odrv4 I__4990 (
            .O(N__24034),
            .I(data_in_3_7));
    LocalMux I__4989 (
            .O(N__24031),
            .I(data_in_3_7));
    Odrv4 I__4988 (
            .O(N__24026),
            .I(data_in_3_7));
    CascadeMux I__4987 (
            .O(N__24019),
            .I(N__24016));
    InMux I__4986 (
            .O(N__24016),
            .I(N__24012));
    InMux I__4985 (
            .O(N__24015),
            .I(N__24009));
    LocalMux I__4984 (
            .O(N__24012),
            .I(N__24004));
    LocalMux I__4983 (
            .O(N__24009),
            .I(N__24004));
    Span4Mux_s3_v I__4982 (
            .O(N__24004),
            .I(N__24000));
    InMux I__4981 (
            .O(N__24003),
            .I(N__23997));
    Span4Mux_v I__4980 (
            .O(N__24000),
            .I(N__23994));
    LocalMux I__4979 (
            .O(N__23997),
            .I(N__23991));
    Odrv4 I__4978 (
            .O(N__23994),
            .I(data_in_17_5));
    Odrv4 I__4977 (
            .O(N__23991),
            .I(data_in_17_5));
    CascadeMux I__4976 (
            .O(N__23986),
            .I(N__23983));
    InMux I__4975 (
            .O(N__23983),
            .I(N__23980));
    LocalMux I__4974 (
            .O(N__23980),
            .I(N__23976));
    InMux I__4973 (
            .O(N__23979),
            .I(N__23973));
    Span4Mux_h I__4972 (
            .O(N__23976),
            .I(N__23969));
    LocalMux I__4971 (
            .O(N__23973),
            .I(N__23966));
    InMux I__4970 (
            .O(N__23972),
            .I(N__23963));
    Odrv4 I__4969 (
            .O(N__23969),
            .I(data_in_7_1));
    Odrv4 I__4968 (
            .O(N__23966),
            .I(data_in_7_1));
    LocalMux I__4967 (
            .O(N__23963),
            .I(data_in_7_1));
    InMux I__4966 (
            .O(N__23956),
            .I(N__23953));
    LocalMux I__4965 (
            .O(N__23953),
            .I(N__23950));
    Span4Mux_s2_v I__4964 (
            .O(N__23950),
            .I(N__23945));
    InMux I__4963 (
            .O(N__23949),
            .I(N__23940));
    InMux I__4962 (
            .O(N__23948),
            .I(N__23940));
    Span4Mux_h I__4961 (
            .O(N__23945),
            .I(N__23937));
    LocalMux I__4960 (
            .O(N__23940),
            .I(data_in_6_1));
    Odrv4 I__4959 (
            .O(N__23937),
            .I(data_in_6_1));
    InMux I__4958 (
            .O(N__23932),
            .I(N__23929));
    LocalMux I__4957 (
            .O(N__23929),
            .I(N__23925));
    InMux I__4956 (
            .O(N__23928),
            .I(N__23922));
    Span4Mux_h I__4955 (
            .O(N__23925),
            .I(N__23915));
    LocalMux I__4954 (
            .O(N__23922),
            .I(N__23915));
    InMux I__4953 (
            .O(N__23921),
            .I(N__23912));
    InMux I__4952 (
            .O(N__23920),
            .I(N__23908));
    Span4Mux_v I__4951 (
            .O(N__23915),
            .I(N__23903));
    LocalMux I__4950 (
            .O(N__23912),
            .I(N__23903));
    InMux I__4949 (
            .O(N__23911),
            .I(N__23900));
    LocalMux I__4948 (
            .O(N__23908),
            .I(\c0.data_in_field_141 ));
    Odrv4 I__4947 (
            .O(N__23903),
            .I(\c0.data_in_field_141 ));
    LocalMux I__4946 (
            .O(N__23900),
            .I(\c0.data_in_field_141 ));
    InMux I__4945 (
            .O(N__23893),
            .I(N__23888));
    InMux I__4944 (
            .O(N__23892),
            .I(N__23885));
    InMux I__4943 (
            .O(N__23891),
            .I(N__23882));
    LocalMux I__4942 (
            .O(N__23888),
            .I(N__23879));
    LocalMux I__4941 (
            .O(N__23885),
            .I(N__23876));
    LocalMux I__4940 (
            .O(N__23882),
            .I(N__23873));
    Span4Mux_h I__4939 (
            .O(N__23879),
            .I(N__23868));
    Span4Mux_s2_v I__4938 (
            .O(N__23876),
            .I(N__23868));
    Span4Mux_v I__4937 (
            .O(N__23873),
            .I(N__23865));
    Span4Mux_h I__4936 (
            .O(N__23868),
            .I(N__23861));
    Span4Mux_v I__4935 (
            .O(N__23865),
            .I(N__23858));
    InMux I__4934 (
            .O(N__23864),
            .I(N__23855));
    Span4Mux_v I__4933 (
            .O(N__23861),
            .I(N__23852));
    Odrv4 I__4932 (
            .O(N__23858),
            .I(data_in_1_6));
    LocalMux I__4931 (
            .O(N__23855),
            .I(data_in_1_6));
    Odrv4 I__4930 (
            .O(N__23852),
            .I(data_in_1_6));
    InMux I__4929 (
            .O(N__23845),
            .I(N__23841));
    InMux I__4928 (
            .O(N__23844),
            .I(N__23838));
    LocalMux I__4927 (
            .O(N__23841),
            .I(N__23835));
    LocalMux I__4926 (
            .O(N__23838),
            .I(N__23832));
    Span4Mux_h I__4925 (
            .O(N__23835),
            .I(N__23829));
    Span4Mux_v I__4924 (
            .O(N__23832),
            .I(N__23825));
    Span4Mux_s0_v I__4923 (
            .O(N__23829),
            .I(N__23822));
    InMux I__4922 (
            .O(N__23828),
            .I(N__23819));
    Odrv4 I__4921 (
            .O(N__23825),
            .I(data_in_9_7));
    Odrv4 I__4920 (
            .O(N__23822),
            .I(data_in_9_7));
    LocalMux I__4919 (
            .O(N__23819),
            .I(data_in_9_7));
    CascadeMux I__4918 (
            .O(N__23812),
            .I(N__23809));
    InMux I__4917 (
            .O(N__23809),
            .I(N__23806));
    LocalMux I__4916 (
            .O(N__23806),
            .I(N__23803));
    Span12Mux_v I__4915 (
            .O(N__23803),
            .I(N__23798));
    InMux I__4914 (
            .O(N__23802),
            .I(N__23793));
    InMux I__4913 (
            .O(N__23801),
            .I(N__23793));
    Odrv12 I__4912 (
            .O(N__23798),
            .I(data_in_6_7));
    LocalMux I__4911 (
            .O(N__23793),
            .I(data_in_6_7));
    InMux I__4910 (
            .O(N__23788),
            .I(N__23784));
    InMux I__4909 (
            .O(N__23787),
            .I(N__23781));
    LocalMux I__4908 (
            .O(N__23784),
            .I(N__23778));
    LocalMux I__4907 (
            .O(N__23781),
            .I(N__23775));
    Span4Mux_h I__4906 (
            .O(N__23778),
            .I(N__23768));
    Span4Mux_h I__4905 (
            .O(N__23775),
            .I(N__23768));
    InMux I__4904 (
            .O(N__23774),
            .I(N__23763));
    InMux I__4903 (
            .O(N__23773),
            .I(N__23763));
    Odrv4 I__4902 (
            .O(N__23768),
            .I(data_in_3_1));
    LocalMux I__4901 (
            .O(N__23763),
            .I(data_in_3_1));
    InMux I__4900 (
            .O(N__23758),
            .I(N__23754));
    InMux I__4899 (
            .O(N__23757),
            .I(N__23751));
    LocalMux I__4898 (
            .O(N__23754),
            .I(N__23747));
    LocalMux I__4897 (
            .O(N__23751),
            .I(N__23744));
    InMux I__4896 (
            .O(N__23750),
            .I(N__23741));
    Span4Mux_v I__4895 (
            .O(N__23747),
            .I(N__23736));
    Span4Mux_h I__4894 (
            .O(N__23744),
            .I(N__23731));
    LocalMux I__4893 (
            .O(N__23741),
            .I(N__23731));
    CascadeMux I__4892 (
            .O(N__23740),
            .I(N__23728));
    InMux I__4891 (
            .O(N__23739),
            .I(N__23725));
    Span4Mux_h I__4890 (
            .O(N__23736),
            .I(N__23722));
    Span4Mux_v I__4889 (
            .O(N__23731),
            .I(N__23719));
    InMux I__4888 (
            .O(N__23728),
            .I(N__23716));
    LocalMux I__4887 (
            .O(N__23725),
            .I(\c0.data_in_field_21 ));
    Odrv4 I__4886 (
            .O(N__23722),
            .I(\c0.data_in_field_21 ));
    Odrv4 I__4885 (
            .O(N__23719),
            .I(\c0.data_in_field_21 ));
    LocalMux I__4884 (
            .O(N__23716),
            .I(\c0.data_in_field_21 ));
    CascadeMux I__4883 (
            .O(N__23707),
            .I(N__23704));
    InMux I__4882 (
            .O(N__23704),
            .I(N__23701));
    LocalMux I__4881 (
            .O(N__23701),
            .I(N__23698));
    Span12Mux_s8_h I__4880 (
            .O(N__23698),
            .I(N__23695));
    Odrv12 I__4879 (
            .O(N__23695),
            .I(\c0.n5881 ));
    InMux I__4878 (
            .O(N__23692),
            .I(N__23688));
    InMux I__4877 (
            .O(N__23691),
            .I(N__23685));
    LocalMux I__4876 (
            .O(N__23688),
            .I(N__23682));
    LocalMux I__4875 (
            .O(N__23685),
            .I(N__23679));
    Span4Mux_v I__4874 (
            .O(N__23682),
            .I(N__23676));
    Span4Mux_h I__4873 (
            .O(N__23679),
            .I(N__23673));
    Span4Mux_s2_v I__4872 (
            .O(N__23676),
            .I(N__23669));
    Span4Mux_h I__4871 (
            .O(N__23673),
            .I(N__23666));
    InMux I__4870 (
            .O(N__23672),
            .I(N__23663));
    Odrv4 I__4869 (
            .O(N__23669),
            .I(data_in_15_6));
    Odrv4 I__4868 (
            .O(N__23666),
            .I(data_in_15_6));
    LocalMux I__4867 (
            .O(N__23663),
            .I(data_in_15_6));
    CascadeMux I__4866 (
            .O(N__23656),
            .I(N__23653));
    InMux I__4865 (
            .O(N__23653),
            .I(N__23648));
    InMux I__4864 (
            .O(N__23652),
            .I(N__23643));
    InMux I__4863 (
            .O(N__23651),
            .I(N__23643));
    LocalMux I__4862 (
            .O(N__23648),
            .I(\c0.data_in_field_29 ));
    LocalMux I__4861 (
            .O(N__23643),
            .I(\c0.data_in_field_29 ));
    InMux I__4860 (
            .O(N__23638),
            .I(N__23635));
    LocalMux I__4859 (
            .O(N__23635),
            .I(N__23632));
    Span4Mux_h I__4858 (
            .O(N__23632),
            .I(N__23629));
    Span4Mux_h I__4857 (
            .O(N__23629),
            .I(N__23626));
    Odrv4 I__4856 (
            .O(N__23626),
            .I(\c0.n2046 ));
    InMux I__4855 (
            .O(N__23623),
            .I(N__23620));
    LocalMux I__4854 (
            .O(N__23620),
            .I(N__23615));
    InMux I__4853 (
            .O(N__23619),
            .I(N__23612));
    InMux I__4852 (
            .O(N__23618),
            .I(N__23609));
    Span4Mux_h I__4851 (
            .O(N__23615),
            .I(N__23604));
    LocalMux I__4850 (
            .O(N__23612),
            .I(N__23604));
    LocalMux I__4849 (
            .O(N__23609),
            .I(N__23601));
    Span4Mux_h I__4848 (
            .O(N__23604),
            .I(N__23597));
    Span4Mux_h I__4847 (
            .O(N__23601),
            .I(N__23594));
    InMux I__4846 (
            .O(N__23600),
            .I(N__23591));
    Span4Mux_h I__4845 (
            .O(N__23597),
            .I(N__23588));
    Span4Mux_h I__4844 (
            .O(N__23594),
            .I(N__23585));
    LocalMux I__4843 (
            .O(N__23591),
            .I(\c0.data_in_field_85 ));
    Odrv4 I__4842 (
            .O(N__23588),
            .I(\c0.data_in_field_85 ));
    Odrv4 I__4841 (
            .O(N__23585),
            .I(\c0.data_in_field_85 ));
    CascadeMux I__4840 (
            .O(N__23578),
            .I(\c0.n2046_cascade_ ));
    InMux I__4839 (
            .O(N__23575),
            .I(N__23572));
    LocalMux I__4838 (
            .O(N__23572),
            .I(N__23568));
    InMux I__4837 (
            .O(N__23571),
            .I(N__23565));
    Span4Mux_h I__4836 (
            .O(N__23568),
            .I(N__23562));
    LocalMux I__4835 (
            .O(N__23565),
            .I(N__23559));
    Odrv4 I__4834 (
            .O(N__23562),
            .I(\c0.n5108 ));
    Odrv12 I__4833 (
            .O(N__23559),
            .I(\c0.n5108 ));
    InMux I__4832 (
            .O(N__23554),
            .I(N__23550));
    InMux I__4831 (
            .O(N__23553),
            .I(N__23547));
    LocalMux I__4830 (
            .O(N__23550),
            .I(N__23543));
    LocalMux I__4829 (
            .O(N__23547),
            .I(N__23540));
    InMux I__4828 (
            .O(N__23546),
            .I(N__23536));
    Span4Mux_h I__4827 (
            .O(N__23543),
            .I(N__23532));
    Span4Mux_v I__4826 (
            .O(N__23540),
            .I(N__23529));
    InMux I__4825 (
            .O(N__23539),
            .I(N__23526));
    LocalMux I__4824 (
            .O(N__23536),
            .I(N__23523));
    InMux I__4823 (
            .O(N__23535),
            .I(N__23520));
    Span4Mux_h I__4822 (
            .O(N__23532),
            .I(N__23517));
    Span4Mux_h I__4821 (
            .O(N__23529),
            .I(N__23512));
    LocalMux I__4820 (
            .O(N__23526),
            .I(N__23512));
    Span4Mux_v I__4819 (
            .O(N__23523),
            .I(N__23509));
    LocalMux I__4818 (
            .O(N__23520),
            .I(\c0.data_in_field_89 ));
    Odrv4 I__4817 (
            .O(N__23517),
            .I(\c0.data_in_field_89 ));
    Odrv4 I__4816 (
            .O(N__23512),
            .I(\c0.data_in_field_89 ));
    Odrv4 I__4815 (
            .O(N__23509),
            .I(\c0.data_in_field_89 ));
    InMux I__4814 (
            .O(N__23500),
            .I(N__23496));
    InMux I__4813 (
            .O(N__23499),
            .I(N__23493));
    LocalMux I__4812 (
            .O(N__23496),
            .I(N__23488));
    LocalMux I__4811 (
            .O(N__23493),
            .I(N__23485));
    InMux I__4810 (
            .O(N__23492),
            .I(N__23482));
    InMux I__4809 (
            .O(N__23491),
            .I(N__23479));
    Span4Mux_v I__4808 (
            .O(N__23488),
            .I(N__23472));
    Span4Mux_h I__4807 (
            .O(N__23485),
            .I(N__23472));
    LocalMux I__4806 (
            .O(N__23482),
            .I(N__23472));
    LocalMux I__4805 (
            .O(N__23479),
            .I(N__23469));
    Span4Mux_h I__4804 (
            .O(N__23472),
            .I(N__23464));
    Span4Mux_v I__4803 (
            .O(N__23469),
            .I(N__23461));
    InMux I__4802 (
            .O(N__23468),
            .I(N__23456));
    InMux I__4801 (
            .O(N__23467),
            .I(N__23456));
    Odrv4 I__4800 (
            .O(N__23464),
            .I(\c0.data_in_field_120 ));
    Odrv4 I__4799 (
            .O(N__23461),
            .I(\c0.data_in_field_120 ));
    LocalMux I__4798 (
            .O(N__23456),
            .I(\c0.data_in_field_120 ));
    InMux I__4797 (
            .O(N__23449),
            .I(N__23446));
    LocalMux I__4796 (
            .O(N__23446),
            .I(N__23443));
    Span4Mux_h I__4795 (
            .O(N__23443),
            .I(N__23440));
    Odrv4 I__4794 (
            .O(N__23440),
            .I(\c0.n23_adj_1925 ));
    CascadeMux I__4793 (
            .O(N__23437),
            .I(N__23433));
    InMux I__4792 (
            .O(N__23436),
            .I(N__23429));
    InMux I__4791 (
            .O(N__23433),
            .I(N__23426));
    InMux I__4790 (
            .O(N__23432),
            .I(N__23423));
    LocalMux I__4789 (
            .O(N__23429),
            .I(N__23419));
    LocalMux I__4788 (
            .O(N__23426),
            .I(N__23416));
    LocalMux I__4787 (
            .O(N__23423),
            .I(N__23413));
    InMux I__4786 (
            .O(N__23422),
            .I(N__23410));
    Span12Mux_h I__4785 (
            .O(N__23419),
            .I(N__23407));
    Span4Mux_h I__4784 (
            .O(N__23416),
            .I(N__23404));
    Span4Mux_h I__4783 (
            .O(N__23413),
            .I(N__23401));
    LocalMux I__4782 (
            .O(N__23410),
            .I(\c0.data_in_field_83 ));
    Odrv12 I__4781 (
            .O(N__23407),
            .I(\c0.data_in_field_83 ));
    Odrv4 I__4780 (
            .O(N__23404),
            .I(\c0.data_in_field_83 ));
    Odrv4 I__4779 (
            .O(N__23401),
            .I(\c0.data_in_field_83 ));
    InMux I__4778 (
            .O(N__23392),
            .I(N__23389));
    LocalMux I__4777 (
            .O(N__23389),
            .I(N__23386));
    Span4Mux_v I__4776 (
            .O(N__23386),
            .I(N__23383));
    Odrv4 I__4775 (
            .O(N__23383),
            .I(\c0.n5797 ));
    InMux I__4774 (
            .O(N__23380),
            .I(N__23376));
    InMux I__4773 (
            .O(N__23379),
            .I(N__23373));
    LocalMux I__4772 (
            .O(N__23376),
            .I(N__23369));
    LocalMux I__4771 (
            .O(N__23373),
            .I(N__23366));
    InMux I__4770 (
            .O(N__23372),
            .I(N__23363));
    Span4Mux_v I__4769 (
            .O(N__23369),
            .I(N__23358));
    Span4Mux_h I__4768 (
            .O(N__23366),
            .I(N__23358));
    LocalMux I__4767 (
            .O(N__23363),
            .I(N__23355));
    Span4Mux_h I__4766 (
            .O(N__23358),
            .I(N__23350));
    Span4Mux_h I__4765 (
            .O(N__23355),
            .I(N__23347));
    InMux I__4764 (
            .O(N__23354),
            .I(N__23342));
    InMux I__4763 (
            .O(N__23353),
            .I(N__23342));
    Odrv4 I__4762 (
            .O(N__23350),
            .I(\c0.data_in_field_19 ));
    Odrv4 I__4761 (
            .O(N__23347),
            .I(\c0.data_in_field_19 ));
    LocalMux I__4760 (
            .O(N__23342),
            .I(\c0.data_in_field_19 ));
    InMux I__4759 (
            .O(N__23335),
            .I(N__23332));
    LocalMux I__4758 (
            .O(N__23332),
            .I(N__23329));
    Span4Mux_h I__4757 (
            .O(N__23329),
            .I(N__23326));
    Odrv4 I__4756 (
            .O(N__23326),
            .I(\c0.n23 ));
    CascadeMux I__4755 (
            .O(N__23323),
            .I(N__23320));
    InMux I__4754 (
            .O(N__23320),
            .I(N__23316));
    InMux I__4753 (
            .O(N__23319),
            .I(N__23313));
    LocalMux I__4752 (
            .O(N__23316),
            .I(N__23309));
    LocalMux I__4751 (
            .O(N__23313),
            .I(N__23306));
    InMux I__4750 (
            .O(N__23312),
            .I(N__23302));
    Span4Mux_v I__4749 (
            .O(N__23309),
            .I(N__23299));
    Span4Mux_h I__4748 (
            .O(N__23306),
            .I(N__23296));
    InMux I__4747 (
            .O(N__23305),
            .I(N__23293));
    LocalMux I__4746 (
            .O(N__23302),
            .I(N__23290));
    Span4Mux_h I__4745 (
            .O(N__23299),
            .I(N__23287));
    Span4Mux_h I__4744 (
            .O(N__23296),
            .I(N__23284));
    LocalMux I__4743 (
            .O(N__23293),
            .I(data_in_3_3));
    Odrv12 I__4742 (
            .O(N__23290),
            .I(data_in_3_3));
    Odrv4 I__4741 (
            .O(N__23287),
            .I(data_in_3_3));
    Odrv4 I__4740 (
            .O(N__23284),
            .I(data_in_3_3));
    InMux I__4739 (
            .O(N__23275),
            .I(N__23272));
    LocalMux I__4738 (
            .O(N__23272),
            .I(N__23269));
    Span4Mux_s2_v I__4737 (
            .O(N__23269),
            .I(N__23266));
    Span4Mux_h I__4736 (
            .O(N__23266),
            .I(N__23263));
    Odrv4 I__4735 (
            .O(N__23263),
            .I(\c0.n25_adj_1960 ));
    CascadeMux I__4734 (
            .O(N__23260),
            .I(N__23257));
    InMux I__4733 (
            .O(N__23257),
            .I(N__23252));
    InMux I__4732 (
            .O(N__23256),
            .I(N__23249));
    InMux I__4731 (
            .O(N__23255),
            .I(N__23245));
    LocalMux I__4730 (
            .O(N__23252),
            .I(N__23240));
    LocalMux I__4729 (
            .O(N__23249),
            .I(N__23240));
    InMux I__4728 (
            .O(N__23248),
            .I(N__23236));
    LocalMux I__4727 (
            .O(N__23245),
            .I(N__23233));
    Span4Mux_v I__4726 (
            .O(N__23240),
            .I(N__23230));
    InMux I__4725 (
            .O(N__23239),
            .I(N__23227));
    LocalMux I__4724 (
            .O(N__23236),
            .I(N__23222));
    Span4Mux_h I__4723 (
            .O(N__23233),
            .I(N__23222));
    Odrv4 I__4722 (
            .O(N__23230),
            .I(\c0.data_in_field_67 ));
    LocalMux I__4721 (
            .O(N__23227),
            .I(\c0.data_in_field_67 ));
    Odrv4 I__4720 (
            .O(N__23222),
            .I(\c0.data_in_field_67 ));
    InMux I__4719 (
            .O(N__23215),
            .I(N__23212));
    LocalMux I__4718 (
            .O(N__23212),
            .I(N__23208));
    InMux I__4717 (
            .O(N__23211),
            .I(N__23205));
    Span4Mux_h I__4716 (
            .O(N__23208),
            .I(N__23202));
    LocalMux I__4715 (
            .O(N__23205),
            .I(N__23199));
    Span4Mux_v I__4714 (
            .O(N__23202),
            .I(N__23194));
    Span4Mux_v I__4713 (
            .O(N__23199),
            .I(N__23194));
    Odrv4 I__4712 (
            .O(N__23194),
            .I(\c0.n5093 ));
    InMux I__4711 (
            .O(N__23191),
            .I(N__23188));
    LocalMux I__4710 (
            .O(N__23188),
            .I(N__23185));
    Span4Mux_h I__4709 (
            .O(N__23185),
            .I(N__23182));
    Odrv4 I__4708 (
            .O(N__23182),
            .I(\c0.n5162 ));
    InMux I__4707 (
            .O(N__23179),
            .I(N__23176));
    LocalMux I__4706 (
            .O(N__23176),
            .I(N__23172));
    InMux I__4705 (
            .O(N__23175),
            .I(N__23169));
    Odrv12 I__4704 (
            .O(N__23172),
            .I(\c0.n5213 ));
    LocalMux I__4703 (
            .O(N__23169),
            .I(\c0.n5213 ));
    CascadeMux I__4702 (
            .O(N__23164),
            .I(\c0.n5099_cascade_ ));
    InMux I__4701 (
            .O(N__23161),
            .I(N__23158));
    LocalMux I__4700 (
            .O(N__23158),
            .I(N__23155));
    Span4Mux_h I__4699 (
            .O(N__23155),
            .I(N__23152));
    Odrv4 I__4698 (
            .O(N__23152),
            .I(\c0.n19 ));
    InMux I__4697 (
            .O(N__23149),
            .I(N__23145));
    CascadeMux I__4696 (
            .O(N__23148),
            .I(N__23142));
    LocalMux I__4695 (
            .O(N__23145),
            .I(N__23139));
    InMux I__4694 (
            .O(N__23142),
            .I(N__23135));
    Span4Mux_h I__4693 (
            .O(N__23139),
            .I(N__23132));
    InMux I__4692 (
            .O(N__23138),
            .I(N__23129));
    LocalMux I__4691 (
            .O(N__23135),
            .I(\c0.data_in_field_104 ));
    Odrv4 I__4690 (
            .O(N__23132),
            .I(\c0.data_in_field_104 ));
    LocalMux I__4689 (
            .O(N__23129),
            .I(\c0.data_in_field_104 ));
    InMux I__4688 (
            .O(N__23122),
            .I(N__23119));
    LocalMux I__4687 (
            .O(N__23119),
            .I(N__23116));
    Span4Mux_v I__4686 (
            .O(N__23116),
            .I(N__23113));
    Span4Mux_h I__4685 (
            .O(N__23113),
            .I(N__23108));
    InMux I__4684 (
            .O(N__23112),
            .I(N__23103));
    InMux I__4683 (
            .O(N__23111),
            .I(N__23103));
    Odrv4 I__4682 (
            .O(N__23108),
            .I(data_in_0_6));
    LocalMux I__4681 (
            .O(N__23103),
            .I(data_in_0_6));
    CascadeMux I__4680 (
            .O(N__23098),
            .I(N__23095));
    InMux I__4679 (
            .O(N__23095),
            .I(N__23090));
    InMux I__4678 (
            .O(N__23094),
            .I(N__23085));
    InMux I__4677 (
            .O(N__23093),
            .I(N__23085));
    LocalMux I__4676 (
            .O(N__23090),
            .I(data_in_12_0));
    LocalMux I__4675 (
            .O(N__23085),
            .I(data_in_12_0));
    InMux I__4674 (
            .O(N__23080),
            .I(N__23077));
    LocalMux I__4673 (
            .O(N__23077),
            .I(N__23074));
    Span4Mux_h I__4672 (
            .O(N__23074),
            .I(N__23071));
    Odrv4 I__4671 (
            .O(N__23071),
            .I(\c0.n13 ));
    InMux I__4670 (
            .O(N__23068),
            .I(N__23064));
    InMux I__4669 (
            .O(N__23067),
            .I(N__23061));
    LocalMux I__4668 (
            .O(N__23064),
            .I(N__23058));
    LocalMux I__4667 (
            .O(N__23061),
            .I(N__23055));
    Span4Mux_v I__4666 (
            .O(N__23058),
            .I(N__23051));
    Span4Mux_v I__4665 (
            .O(N__23055),
            .I(N__23048));
    CascadeMux I__4664 (
            .O(N__23054),
            .I(N__23044));
    Span4Mux_h I__4663 (
            .O(N__23051),
            .I(N__23041));
    Span4Mux_h I__4662 (
            .O(N__23048),
            .I(N__23038));
    InMux I__4661 (
            .O(N__23047),
            .I(N__23033));
    InMux I__4660 (
            .O(N__23044),
            .I(N__23033));
    Odrv4 I__4659 (
            .O(N__23041),
            .I(\c0.data_in_field_117 ));
    Odrv4 I__4658 (
            .O(N__23038),
            .I(\c0.data_in_field_117 ));
    LocalMux I__4657 (
            .O(N__23033),
            .I(\c0.data_in_field_117 ));
    CascadeMux I__4656 (
            .O(N__23026),
            .I(\c0.n2074_cascade_ ));
    CascadeMux I__4655 (
            .O(N__23023),
            .I(N__23020));
    InMux I__4654 (
            .O(N__23020),
            .I(N__23017));
    LocalMux I__4653 (
            .O(N__23017),
            .I(N__23014));
    Span4Mux_h I__4652 (
            .O(N__23014),
            .I(N__23011));
    Odrv4 I__4651 (
            .O(N__23011),
            .I(\c0.n10_adj_1888 ));
    InMux I__4650 (
            .O(N__23008),
            .I(N__23004));
    InMux I__4649 (
            .O(N__23007),
            .I(N__23001));
    LocalMux I__4648 (
            .O(N__23004),
            .I(N__22998));
    LocalMux I__4647 (
            .O(N__23001),
            .I(N__22992));
    Span4Mux_h I__4646 (
            .O(N__22998),
            .I(N__22989));
    InMux I__4645 (
            .O(N__22997),
            .I(N__22982));
    InMux I__4644 (
            .O(N__22996),
            .I(N__22982));
    InMux I__4643 (
            .O(N__22995),
            .I(N__22982));
    Odrv4 I__4642 (
            .O(N__22992),
            .I(\c0.data_in_field_95 ));
    Odrv4 I__4641 (
            .O(N__22989),
            .I(\c0.data_in_field_95 ));
    LocalMux I__4640 (
            .O(N__22982),
            .I(\c0.data_in_field_95 ));
    InMux I__4639 (
            .O(N__22975),
            .I(N__22972));
    LocalMux I__4638 (
            .O(N__22972),
            .I(N__22968));
    CascadeMux I__4637 (
            .O(N__22971),
            .I(N__22965));
    Span4Mux_h I__4636 (
            .O(N__22968),
            .I(N__22962));
    InMux I__4635 (
            .O(N__22965),
            .I(N__22959));
    Odrv4 I__4634 (
            .O(N__22962),
            .I(\c0.n1851 ));
    LocalMux I__4633 (
            .O(N__22959),
            .I(\c0.n1851 ));
    InMux I__4632 (
            .O(N__22954),
            .I(N__22951));
    LocalMux I__4631 (
            .O(N__22951),
            .I(N__22947));
    InMux I__4630 (
            .O(N__22950),
            .I(N__22943));
    Span4Mux_h I__4629 (
            .O(N__22947),
            .I(N__22940));
    InMux I__4628 (
            .O(N__22946),
            .I(N__22937));
    LocalMux I__4627 (
            .O(N__22943),
            .I(N__22933));
    Sp12to4 I__4626 (
            .O(N__22940),
            .I(N__22928));
    LocalMux I__4625 (
            .O(N__22937),
            .I(N__22928));
    CascadeMux I__4624 (
            .O(N__22936),
            .I(N__22922));
    Span4Mux_v I__4623 (
            .O(N__22933),
            .I(N__22919));
    Span12Mux_s7_v I__4622 (
            .O(N__22928),
            .I(N__22916));
    InMux I__4621 (
            .O(N__22927),
            .I(N__22911));
    InMux I__4620 (
            .O(N__22926),
            .I(N__22911));
    InMux I__4619 (
            .O(N__22925),
            .I(N__22906));
    InMux I__4618 (
            .O(N__22922),
            .I(N__22906));
    Odrv4 I__4617 (
            .O(N__22919),
            .I(\c0.data_in_field_96 ));
    Odrv12 I__4616 (
            .O(N__22916),
            .I(\c0.data_in_field_96 ));
    LocalMux I__4615 (
            .O(N__22911),
            .I(\c0.data_in_field_96 ));
    LocalMux I__4614 (
            .O(N__22906),
            .I(\c0.data_in_field_96 ));
    InMux I__4613 (
            .O(N__22897),
            .I(N__22894));
    LocalMux I__4612 (
            .O(N__22894),
            .I(N__22891));
    Odrv12 I__4611 (
            .O(N__22891),
            .I(\c0.n5099 ));
    CascadeMux I__4610 (
            .O(N__22888),
            .I(\c0.n5447_cascade_ ));
    CascadeMux I__4609 (
            .O(N__22885),
            .I(\c0.n5755_cascade_ ));
    InMux I__4608 (
            .O(N__22882),
            .I(N__22879));
    LocalMux I__4607 (
            .O(N__22879),
            .I(N__22876));
    Span12Mux_s9_v I__4606 (
            .O(N__22876),
            .I(N__22873));
    Odrv12 I__4605 (
            .O(N__22873),
            .I(\c0.n5758 ));
    InMux I__4604 (
            .O(N__22870),
            .I(N__22866));
    InMux I__4603 (
            .O(N__22869),
            .I(N__22861));
    LocalMux I__4602 (
            .O(N__22866),
            .I(N__22858));
    InMux I__4601 (
            .O(N__22865),
            .I(N__22855));
    InMux I__4600 (
            .O(N__22864),
            .I(N__22852));
    LocalMux I__4599 (
            .O(N__22861),
            .I(N__22849));
    Span12Mux_s5_h I__4598 (
            .O(N__22858),
            .I(N__22846));
    LocalMux I__4597 (
            .O(N__22855),
            .I(N__22843));
    LocalMux I__4596 (
            .O(N__22852),
            .I(\c0.data_in_field_54 ));
    Odrv12 I__4595 (
            .O(N__22849),
            .I(\c0.data_in_field_54 ));
    Odrv12 I__4594 (
            .O(N__22846),
            .I(\c0.data_in_field_54 ));
    Odrv4 I__4593 (
            .O(N__22843),
            .I(\c0.data_in_field_54 ));
    InMux I__4592 (
            .O(N__22834),
            .I(N__22831));
    LocalMux I__4591 (
            .O(N__22831),
            .I(N__22827));
    InMux I__4590 (
            .O(N__22830),
            .I(N__22824));
    Span4Mux_v I__4589 (
            .O(N__22827),
            .I(N__22818));
    LocalMux I__4588 (
            .O(N__22824),
            .I(N__22815));
    InMux I__4587 (
            .O(N__22823),
            .I(N__22812));
    InMux I__4586 (
            .O(N__22822),
            .I(N__22807));
    InMux I__4585 (
            .O(N__22821),
            .I(N__22807));
    Span4Mux_h I__4584 (
            .O(N__22818),
            .I(N__22800));
    Span4Mux_v I__4583 (
            .O(N__22815),
            .I(N__22800));
    LocalMux I__4582 (
            .O(N__22812),
            .I(N__22800));
    LocalMux I__4581 (
            .O(N__22807),
            .I(\c0.data_in_field_10 ));
    Odrv4 I__4580 (
            .O(N__22800),
            .I(\c0.data_in_field_10 ));
    InMux I__4579 (
            .O(N__22795),
            .I(N__22792));
    LocalMux I__4578 (
            .O(N__22792),
            .I(\c0.n5438 ));
    InMux I__4577 (
            .O(N__22789),
            .I(N__22786));
    LocalMux I__4576 (
            .O(N__22786),
            .I(N__22782));
    InMux I__4575 (
            .O(N__22785),
            .I(N__22779));
    Span4Mux_h I__4574 (
            .O(N__22782),
            .I(N__22773));
    LocalMux I__4573 (
            .O(N__22779),
            .I(N__22773));
    InMux I__4572 (
            .O(N__22778),
            .I(N__22770));
    Span4Mux_v I__4571 (
            .O(N__22773),
            .I(N__22763));
    LocalMux I__4570 (
            .O(N__22770),
            .I(N__22763));
    InMux I__4569 (
            .O(N__22769),
            .I(N__22758));
    InMux I__4568 (
            .O(N__22768),
            .I(N__22758));
    Span4Mux_h I__4567 (
            .O(N__22763),
            .I(N__22755));
    LocalMux I__4566 (
            .O(N__22758),
            .I(\c0.data_in_field_82 ));
    Odrv4 I__4565 (
            .O(N__22755),
            .I(\c0.data_in_field_82 ));
    CascadeMux I__4564 (
            .O(N__22750),
            .I(\c0.n5767_cascade_ ));
    InMux I__4563 (
            .O(N__22747),
            .I(N__22744));
    LocalMux I__4562 (
            .O(N__22744),
            .I(\c0.n5444 ));
    InMux I__4561 (
            .O(N__22741),
            .I(N__22738));
    LocalMux I__4560 (
            .O(N__22738),
            .I(\c0.n5761 ));
    CascadeMux I__4559 (
            .O(N__22735),
            .I(N__22731));
    InMux I__4558 (
            .O(N__22734),
            .I(N__22728));
    InMux I__4557 (
            .O(N__22731),
            .I(N__22725));
    LocalMux I__4556 (
            .O(N__22728),
            .I(N__22722));
    LocalMux I__4555 (
            .O(N__22725),
            .I(N__22718));
    Span4Mux_h I__4554 (
            .O(N__22722),
            .I(N__22715));
    InMux I__4553 (
            .O(N__22721),
            .I(N__22712));
    Odrv12 I__4552 (
            .O(N__22718),
            .I(data_in_11_7));
    Odrv4 I__4551 (
            .O(N__22715),
            .I(data_in_11_7));
    LocalMux I__4550 (
            .O(N__22712),
            .I(data_in_11_7));
    CascadeMux I__4549 (
            .O(N__22705),
            .I(N__22702));
    InMux I__4548 (
            .O(N__22702),
            .I(N__22699));
    LocalMux I__4547 (
            .O(N__22699),
            .I(N__22696));
    Span4Mux_h I__4546 (
            .O(N__22696),
            .I(N__22691));
    InMux I__4545 (
            .O(N__22695),
            .I(N__22688));
    InMux I__4544 (
            .O(N__22694),
            .I(N__22685));
    Odrv4 I__4543 (
            .O(N__22691),
            .I(data_in_10_7));
    LocalMux I__4542 (
            .O(N__22688),
            .I(data_in_10_7));
    LocalMux I__4541 (
            .O(N__22685),
            .I(data_in_10_7));
    CascadeMux I__4540 (
            .O(N__22678),
            .I(N__22675));
    InMux I__4539 (
            .O(N__22675),
            .I(N__22672));
    LocalMux I__4538 (
            .O(N__22672),
            .I(N__22667));
    InMux I__4537 (
            .O(N__22671),
            .I(N__22664));
    InMux I__4536 (
            .O(N__22670),
            .I(N__22660));
    Span4Mux_v I__4535 (
            .O(N__22667),
            .I(N__22655));
    LocalMux I__4534 (
            .O(N__22664),
            .I(N__22655));
    InMux I__4533 (
            .O(N__22663),
            .I(N__22652));
    LocalMux I__4532 (
            .O(N__22660),
            .I(data_in_2_7));
    Odrv4 I__4531 (
            .O(N__22655),
            .I(data_in_2_7));
    LocalMux I__4530 (
            .O(N__22652),
            .I(data_in_2_7));
    InMux I__4529 (
            .O(N__22645),
            .I(N__22642));
    LocalMux I__4528 (
            .O(N__22642),
            .I(\c0.n27_adj_1956 ));
    CascadeMux I__4527 (
            .O(N__22639),
            .I(N__22636));
    InMux I__4526 (
            .O(N__22636),
            .I(N__22633));
    LocalMux I__4525 (
            .O(N__22633),
            .I(N__22630));
    Odrv4 I__4524 (
            .O(N__22630),
            .I(\c0.n26_adj_1958 ));
    InMux I__4523 (
            .O(N__22627),
            .I(N__22624));
    LocalMux I__4522 (
            .O(N__22624),
            .I(N__22619));
    CascadeMux I__4521 (
            .O(N__22623),
            .I(N__22616));
    InMux I__4520 (
            .O(N__22622),
            .I(N__22613));
    Span4Mux_s1_h I__4519 (
            .O(N__22619),
            .I(N__22610));
    InMux I__4518 (
            .O(N__22616),
            .I(N__22607));
    LocalMux I__4517 (
            .O(N__22613),
            .I(N__22604));
    Span4Mux_h I__4516 (
            .O(N__22610),
            .I(N__22598));
    LocalMux I__4515 (
            .O(N__22607),
            .I(N__22598));
    Span4Mux_h I__4514 (
            .O(N__22604),
            .I(N__22594));
    InMux I__4513 (
            .O(N__22603),
            .I(N__22591));
    Sp12to4 I__4512 (
            .O(N__22598),
            .I(N__22588));
    InMux I__4511 (
            .O(N__22597),
            .I(N__22585));
    Span4Mux_v I__4510 (
            .O(N__22594),
            .I(N__22582));
    LocalMux I__4509 (
            .O(N__22591),
            .I(\c0.data_in_field_135 ));
    Odrv12 I__4508 (
            .O(N__22588),
            .I(\c0.data_in_field_135 ));
    LocalMux I__4507 (
            .O(N__22585),
            .I(\c0.data_in_field_135 ));
    Odrv4 I__4506 (
            .O(N__22582),
            .I(\c0.data_in_field_135 ));
    InMux I__4505 (
            .O(N__22573),
            .I(N__22568));
    CascadeMux I__4504 (
            .O(N__22572),
            .I(N__22564));
    InMux I__4503 (
            .O(N__22571),
            .I(N__22561));
    LocalMux I__4502 (
            .O(N__22568),
            .I(N__22558));
    InMux I__4501 (
            .O(N__22567),
            .I(N__22555));
    InMux I__4500 (
            .O(N__22564),
            .I(N__22552));
    LocalMux I__4499 (
            .O(N__22561),
            .I(N__22549));
    Span4Mux_v I__4498 (
            .O(N__22558),
            .I(N__22546));
    LocalMux I__4497 (
            .O(N__22555),
            .I(N__22541));
    LocalMux I__4496 (
            .O(N__22552),
            .I(N__22541));
    Odrv4 I__4495 (
            .O(N__22549),
            .I(\c0.data_in_field_113 ));
    Odrv4 I__4494 (
            .O(N__22546),
            .I(\c0.data_in_field_113 ));
    Odrv4 I__4493 (
            .O(N__22541),
            .I(\c0.data_in_field_113 ));
    InMux I__4492 (
            .O(N__22534),
            .I(N__22530));
    InMux I__4491 (
            .O(N__22533),
            .I(N__22527));
    LocalMux I__4490 (
            .O(N__22530),
            .I(\c0.n1772 ));
    LocalMux I__4489 (
            .O(N__22527),
            .I(\c0.n1772 ));
    InMux I__4488 (
            .O(N__22522),
            .I(N__22519));
    LocalMux I__4487 (
            .O(N__22519),
            .I(N__22516));
    Span4Mux_v I__4486 (
            .O(N__22516),
            .I(N__22513));
    Span4Mux_v I__4485 (
            .O(N__22513),
            .I(N__22510));
    Odrv4 I__4484 (
            .O(N__22510),
            .I(\c0.n5144 ));
    CascadeMux I__4483 (
            .O(N__22507),
            .I(\c0.n5144_cascade_ ));
    InMux I__4482 (
            .O(N__22504),
            .I(N__22501));
    LocalMux I__4481 (
            .O(N__22501),
            .I(\c0.n31 ));
    CascadeMux I__4480 (
            .O(N__22498),
            .I(N__22494));
    InMux I__4479 (
            .O(N__22497),
            .I(N__22491));
    InMux I__4478 (
            .O(N__22494),
            .I(N__22488));
    LocalMux I__4477 (
            .O(N__22491),
            .I(N__22485));
    LocalMux I__4476 (
            .O(N__22488),
            .I(N__22481));
    Span4Mux_h I__4475 (
            .O(N__22485),
            .I(N__22478));
    InMux I__4474 (
            .O(N__22484),
            .I(N__22475));
    Odrv12 I__4473 (
            .O(N__22481),
            .I(data_in_8_5));
    Odrv4 I__4472 (
            .O(N__22478),
            .I(data_in_8_5));
    LocalMux I__4471 (
            .O(N__22475),
            .I(data_in_8_5));
    InMux I__4470 (
            .O(N__22468),
            .I(N__22465));
    LocalMux I__4469 (
            .O(N__22465),
            .I(N__22461));
    InMux I__4468 (
            .O(N__22464),
            .I(N__22458));
    Span4Mux_v I__4467 (
            .O(N__22461),
            .I(N__22454));
    LocalMux I__4466 (
            .O(N__22458),
            .I(N__22451));
    InMux I__4465 (
            .O(N__22457),
            .I(N__22448));
    Odrv4 I__4464 (
            .O(N__22454),
            .I(data_in_8_7));
    Odrv4 I__4463 (
            .O(N__22451),
            .I(data_in_8_7));
    LocalMux I__4462 (
            .O(N__22448),
            .I(data_in_8_7));
    InMux I__4461 (
            .O(N__22441),
            .I(N__22438));
    LocalMux I__4460 (
            .O(N__22438),
            .I(N__22434));
    InMux I__4459 (
            .O(N__22437),
            .I(N__22431));
    Span4Mux_h I__4458 (
            .O(N__22434),
            .I(N__22426));
    LocalMux I__4457 (
            .O(N__22431),
            .I(N__22426));
    Odrv4 I__4456 (
            .O(N__22426),
            .I(\c0.n5249 ));
    InMux I__4455 (
            .O(N__22423),
            .I(N__22420));
    LocalMux I__4454 (
            .O(N__22420),
            .I(N__22417));
    Span4Mux_v I__4453 (
            .O(N__22417),
            .I(N__22413));
    CascadeMux I__4452 (
            .O(N__22416),
            .I(N__22410));
    Span4Mux_s0_v I__4451 (
            .O(N__22413),
            .I(N__22407));
    InMux I__4450 (
            .O(N__22410),
            .I(N__22404));
    Odrv4 I__4449 (
            .O(N__22407),
            .I(rx_data_2));
    LocalMux I__4448 (
            .O(N__22404),
            .I(rx_data_2));
    CascadeMux I__4447 (
            .O(N__22399),
            .I(N__22396));
    InMux I__4446 (
            .O(N__22396),
            .I(N__22393));
    LocalMux I__4445 (
            .O(N__22393),
            .I(N__22390));
    Span4Mux_v I__4444 (
            .O(N__22390),
            .I(N__22386));
    InMux I__4443 (
            .O(N__22389),
            .I(N__22383));
    Span4Mux_h I__4442 (
            .O(N__22386),
            .I(N__22380));
    LocalMux I__4441 (
            .O(N__22383),
            .I(\c0.n5255 ));
    Odrv4 I__4440 (
            .O(N__22380),
            .I(\c0.n5255 ));
    InMux I__4439 (
            .O(N__22375),
            .I(N__22372));
    LocalMux I__4438 (
            .O(N__22372),
            .I(N__22368));
    InMux I__4437 (
            .O(N__22371),
            .I(N__22365));
    Span4Mux_s3_h I__4436 (
            .O(N__22368),
            .I(N__22358));
    LocalMux I__4435 (
            .O(N__22365),
            .I(N__22358));
    InMux I__4434 (
            .O(N__22364),
            .I(N__22355));
    InMux I__4433 (
            .O(N__22363),
            .I(N__22352));
    Span4Mux_v I__4432 (
            .O(N__22358),
            .I(N__22347));
    LocalMux I__4431 (
            .O(N__22355),
            .I(N__22347));
    LocalMux I__4430 (
            .O(N__22352),
            .I(data_in_1_3));
    Odrv4 I__4429 (
            .O(N__22347),
            .I(data_in_1_3));
    InMux I__4428 (
            .O(N__22342),
            .I(N__22339));
    LocalMux I__4427 (
            .O(N__22339),
            .I(N__22336));
    Odrv4 I__4426 (
            .O(N__22336),
            .I(\c0.n28_adj_1954 ));
    InMux I__4425 (
            .O(N__22333),
            .I(N__22330));
    LocalMux I__4424 (
            .O(N__22330),
            .I(N__22327));
    Odrv12 I__4423 (
            .O(N__22327),
            .I(\c0.n26_adj_1955 ));
    CascadeMux I__4422 (
            .O(N__22324),
            .I(\c0.n25_adj_1957_cascade_ ));
    InMux I__4421 (
            .O(N__22321),
            .I(N__22318));
    LocalMux I__4420 (
            .O(N__22318),
            .I(\c0.n4465 ));
    InMux I__4419 (
            .O(N__22315),
            .I(N__22312));
    LocalMux I__4418 (
            .O(N__22312),
            .I(N__22309));
    Span4Mux_h I__4417 (
            .O(N__22309),
            .I(N__22304));
    InMux I__4416 (
            .O(N__22308),
            .I(N__22300));
    InMux I__4415 (
            .O(N__22307),
            .I(N__22297));
    Span4Mux_v I__4414 (
            .O(N__22304),
            .I(N__22294));
    InMux I__4413 (
            .O(N__22303),
            .I(N__22291));
    LocalMux I__4412 (
            .O(N__22300),
            .I(\c0.data_in_field_17 ));
    LocalMux I__4411 (
            .O(N__22297),
            .I(\c0.data_in_field_17 ));
    Odrv4 I__4410 (
            .O(N__22294),
            .I(\c0.data_in_field_17 ));
    LocalMux I__4409 (
            .O(N__22291),
            .I(\c0.data_in_field_17 ));
    CascadeMux I__4408 (
            .O(N__22282),
            .I(N__22278));
    InMux I__4407 (
            .O(N__22281),
            .I(N__22273));
    InMux I__4406 (
            .O(N__22278),
            .I(N__22273));
    LocalMux I__4405 (
            .O(N__22273),
            .I(N__22269));
    InMux I__4404 (
            .O(N__22272),
            .I(N__22266));
    Span4Mux_h I__4403 (
            .O(N__22269),
            .I(N__22262));
    LocalMux I__4402 (
            .O(N__22266),
            .I(N__22259));
    InMux I__4401 (
            .O(N__22265),
            .I(N__22256));
    Span4Mux_v I__4400 (
            .O(N__22262),
            .I(N__22253));
    Odrv4 I__4399 (
            .O(N__22259),
            .I(data_in_1_4));
    LocalMux I__4398 (
            .O(N__22256),
            .I(data_in_1_4));
    Odrv4 I__4397 (
            .O(N__22253),
            .I(data_in_1_4));
    InMux I__4396 (
            .O(N__22246),
            .I(N__22242));
    InMux I__4395 (
            .O(N__22245),
            .I(N__22239));
    LocalMux I__4394 (
            .O(N__22242),
            .I(N__22235));
    LocalMux I__4393 (
            .O(N__22239),
            .I(N__22232));
    InMux I__4392 (
            .O(N__22238),
            .I(N__22228));
    Span4Mux_v I__4391 (
            .O(N__22235),
            .I(N__22225));
    Span4Mux_h I__4390 (
            .O(N__22232),
            .I(N__22222));
    InMux I__4389 (
            .O(N__22231),
            .I(N__22219));
    LocalMux I__4388 (
            .O(N__22228),
            .I(\c0.data_in_field_22 ));
    Odrv4 I__4387 (
            .O(N__22225),
            .I(\c0.data_in_field_22 ));
    Odrv4 I__4386 (
            .O(N__22222),
            .I(\c0.data_in_field_22 ));
    LocalMux I__4385 (
            .O(N__22219),
            .I(\c0.data_in_field_22 ));
    CascadeMux I__4384 (
            .O(N__22210),
            .I(\c0.n2005_cascade_ ));
    CascadeMux I__4383 (
            .O(N__22207),
            .I(\c0.n10_adj_1873_cascade_ ));
    InMux I__4382 (
            .O(N__22204),
            .I(N__22201));
    LocalMux I__4381 (
            .O(N__22201),
            .I(\c0.n1825 ));
    InMux I__4380 (
            .O(N__22198),
            .I(N__22195));
    LocalMux I__4379 (
            .O(N__22195),
            .I(N__22190));
    InMux I__4378 (
            .O(N__22194),
            .I(N__22184));
    InMux I__4377 (
            .O(N__22193),
            .I(N__22184));
    Span4Mux_v I__4376 (
            .O(N__22190),
            .I(N__22181));
    InMux I__4375 (
            .O(N__22189),
            .I(N__22178));
    LocalMux I__4374 (
            .O(N__22184),
            .I(\c0.data_in_field_55 ));
    Odrv4 I__4373 (
            .O(N__22181),
            .I(\c0.data_in_field_55 ));
    LocalMux I__4372 (
            .O(N__22178),
            .I(\c0.data_in_field_55 ));
    InMux I__4371 (
            .O(N__22171),
            .I(N__22168));
    LocalMux I__4370 (
            .O(N__22168),
            .I(\c0.n13_adj_1951 ));
    InMux I__4369 (
            .O(N__22165),
            .I(N__22162));
    LocalMux I__4368 (
            .O(N__22162),
            .I(N__22157));
    InMux I__4367 (
            .O(N__22161),
            .I(N__22154));
    InMux I__4366 (
            .O(N__22160),
            .I(N__22151));
    Span4Mux_h I__4365 (
            .O(N__22157),
            .I(N__22146));
    LocalMux I__4364 (
            .O(N__22154),
            .I(N__22146));
    LocalMux I__4363 (
            .O(N__22151),
            .I(N__22142));
    Span4Mux_v I__4362 (
            .O(N__22146),
            .I(N__22138));
    InMux I__4361 (
            .O(N__22145),
            .I(N__22135));
    Span4Mux_v I__4360 (
            .O(N__22142),
            .I(N__22132));
    InMux I__4359 (
            .O(N__22141),
            .I(N__22129));
    Span4Mux_s2_v I__4358 (
            .O(N__22138),
            .I(N__22126));
    LocalMux I__4357 (
            .O(N__22135),
            .I(\c0.data_in_field_23 ));
    Odrv4 I__4356 (
            .O(N__22132),
            .I(\c0.data_in_field_23 ));
    LocalMux I__4355 (
            .O(N__22129),
            .I(\c0.data_in_field_23 ));
    Odrv4 I__4354 (
            .O(N__22126),
            .I(\c0.data_in_field_23 ));
    CascadeMux I__4353 (
            .O(N__22117),
            .I(N__22114));
    InMux I__4352 (
            .O(N__22114),
            .I(N__22111));
    LocalMux I__4351 (
            .O(N__22111),
            .I(N__22108));
    Span4Mux_v I__4350 (
            .O(N__22108),
            .I(N__22105));
    Odrv4 I__4349 (
            .O(N__22105),
            .I(\c0.n6107 ));
    InMux I__4348 (
            .O(N__22102),
            .I(N__22099));
    LocalMux I__4347 (
            .O(N__22099),
            .I(N__22096));
    Span4Mux_v I__4346 (
            .O(N__22096),
            .I(N__22093));
    Odrv4 I__4345 (
            .O(N__22093),
            .I(\c0.n18_adj_1891 ));
    InMux I__4344 (
            .O(N__22090),
            .I(N__22086));
    InMux I__4343 (
            .O(N__22089),
            .I(N__22083));
    LocalMux I__4342 (
            .O(N__22086),
            .I(\c0.n1978 ));
    LocalMux I__4341 (
            .O(N__22083),
            .I(\c0.n1978 ));
    InMux I__4340 (
            .O(N__22078),
            .I(N__22074));
    InMux I__4339 (
            .O(N__22077),
            .I(N__22071));
    LocalMux I__4338 (
            .O(N__22074),
            .I(N__22068));
    LocalMux I__4337 (
            .O(N__22071),
            .I(\c0.n5261 ));
    Odrv4 I__4336 (
            .O(N__22068),
            .I(\c0.n5261 ));
    CascadeMux I__4335 (
            .O(N__22063),
            .I(\c0.n5689_cascade_ ));
    InMux I__4334 (
            .O(N__22060),
            .I(N__22057));
    LocalMux I__4333 (
            .O(N__22057),
            .I(N__22054));
    Sp12to4 I__4332 (
            .O(N__22054),
            .I(N__22051));
    Span12Mux_v I__4331 (
            .O(N__22051),
            .I(N__22048));
    Odrv12 I__4330 (
            .O(N__22048),
            .I(\c0.n5366 ));
    InMux I__4329 (
            .O(N__22045),
            .I(N__22042));
    LocalMux I__4328 (
            .O(N__22042),
            .I(N__22039));
    Span4Mux_h I__4327 (
            .O(N__22039),
            .I(N__22036));
    Odrv4 I__4326 (
            .O(N__22036),
            .I(\c0.n14_adj_1967 ));
    InMux I__4325 (
            .O(N__22033),
            .I(N__22030));
    LocalMux I__4324 (
            .O(N__22030),
            .I(\c0.n5276 ));
    InMux I__4323 (
            .O(N__22027),
            .I(N__22024));
    LocalMux I__4322 (
            .O(N__22024),
            .I(N__22020));
    InMux I__4321 (
            .O(N__22023),
            .I(N__22017));
    Odrv4 I__4320 (
            .O(N__22020),
            .I(\c0.n5201 ));
    LocalMux I__4319 (
            .O(N__22017),
            .I(\c0.n5201 ));
    CascadeMux I__4318 (
            .O(N__22012),
            .I(\c0.n5276_cascade_ ));
    InMux I__4317 (
            .O(N__22009),
            .I(N__22006));
    LocalMux I__4316 (
            .O(N__22006),
            .I(N__22003));
    Span4Mux_v I__4315 (
            .O(N__22003),
            .I(N__22000));
    Odrv4 I__4314 (
            .O(N__22000),
            .I(\c0.n37 ));
    InMux I__4313 (
            .O(N__21997),
            .I(N__21994));
    LocalMux I__4312 (
            .O(N__21994),
            .I(N__21989));
    InMux I__4311 (
            .O(N__21993),
            .I(N__21986));
    CascadeMux I__4310 (
            .O(N__21992),
            .I(N__21983));
    Span4Mux_v I__4309 (
            .O(N__21989),
            .I(N__21980));
    LocalMux I__4308 (
            .O(N__21986),
            .I(N__21977));
    InMux I__4307 (
            .O(N__21983),
            .I(N__21973));
    Span4Mux_h I__4306 (
            .O(N__21980),
            .I(N__21970));
    Span4Mux_h I__4305 (
            .O(N__21977),
            .I(N__21967));
    InMux I__4304 (
            .O(N__21976),
            .I(N__21964));
    LocalMux I__4303 (
            .O(N__21973),
            .I(\c0.data_in_field_36 ));
    Odrv4 I__4302 (
            .O(N__21970),
            .I(\c0.data_in_field_36 ));
    Odrv4 I__4301 (
            .O(N__21967),
            .I(\c0.data_in_field_36 ));
    LocalMux I__4300 (
            .O(N__21964),
            .I(\c0.data_in_field_36 ));
    InMux I__4299 (
            .O(N__21955),
            .I(N__21951));
    CascadeMux I__4298 (
            .O(N__21954),
            .I(N__21948));
    LocalMux I__4297 (
            .O(N__21951),
            .I(N__21943));
    InMux I__4296 (
            .O(N__21948),
            .I(N__21940));
    InMux I__4295 (
            .O(N__21947),
            .I(N__21935));
    InMux I__4294 (
            .O(N__21946),
            .I(N__21935));
    Span4Mux_h I__4293 (
            .O(N__21943),
            .I(N__21932));
    LocalMux I__4292 (
            .O(N__21940),
            .I(\c0.data_in_field_105 ));
    LocalMux I__4291 (
            .O(N__21935),
            .I(\c0.data_in_field_105 ));
    Odrv4 I__4290 (
            .O(N__21932),
            .I(\c0.data_in_field_105 ));
    CascadeMux I__4289 (
            .O(N__21925),
            .I(\c0.n2095_cascade_ ));
    InMux I__4288 (
            .O(N__21922),
            .I(N__21919));
    LocalMux I__4287 (
            .O(N__21919),
            .I(N__21915));
    InMux I__4286 (
            .O(N__21918),
            .I(N__21912));
    Span4Mux_h I__4285 (
            .O(N__21915),
            .I(N__21909));
    LocalMux I__4284 (
            .O(N__21912),
            .I(N__21906));
    Odrv4 I__4283 (
            .O(N__21909),
            .I(\c0.n1821 ));
    Odrv12 I__4282 (
            .O(N__21906),
            .I(\c0.n1821 ));
    InMux I__4281 (
            .O(N__21901),
            .I(N__21898));
    LocalMux I__4280 (
            .O(N__21898),
            .I(\c0.n34_adj_1896 ));
    InMux I__4279 (
            .O(N__21895),
            .I(N__21891));
    InMux I__4278 (
            .O(N__21894),
            .I(N__21888));
    LocalMux I__4277 (
            .O(N__21891),
            .I(N__21883));
    LocalMux I__4276 (
            .O(N__21888),
            .I(N__21883));
    Span4Mux_v I__4275 (
            .O(N__21883),
            .I(N__21879));
    InMux I__4274 (
            .O(N__21882),
            .I(N__21876));
    Span4Mux_h I__4273 (
            .O(N__21879),
            .I(N__21871));
    LocalMux I__4272 (
            .O(N__21876),
            .I(N__21868));
    InMux I__4271 (
            .O(N__21875),
            .I(N__21863));
    InMux I__4270 (
            .O(N__21874),
            .I(N__21863));
    Odrv4 I__4269 (
            .O(N__21871),
            .I(\c0.data_in_field_11 ));
    Odrv4 I__4268 (
            .O(N__21868),
            .I(\c0.data_in_field_11 ));
    LocalMux I__4267 (
            .O(N__21863),
            .I(\c0.data_in_field_11 ));
    CascadeMux I__4266 (
            .O(N__21856),
            .I(\c0.n5821_cascade_ ));
    InMux I__4265 (
            .O(N__21853),
            .I(N__21850));
    LocalMux I__4264 (
            .O(N__21850),
            .I(N__21847));
    Span4Mux_s3_h I__4263 (
            .O(N__21847),
            .I(N__21844));
    Span4Mux_h I__4262 (
            .O(N__21844),
            .I(N__21841));
    Odrv4 I__4261 (
            .O(N__21841),
            .I(\c0.n5423 ));
    InMux I__4260 (
            .O(N__21838),
            .I(N__21829));
    InMux I__4259 (
            .O(N__21837),
            .I(N__21829));
    InMux I__4258 (
            .O(N__21836),
            .I(N__21829));
    LocalMux I__4257 (
            .O(N__21829),
            .I(\c0.data_in_field_27 ));
    InMux I__4256 (
            .O(N__21826),
            .I(N__21823));
    LocalMux I__4255 (
            .O(N__21823),
            .I(N__21820));
    Span4Mux_h I__4254 (
            .O(N__21820),
            .I(N__21817));
    Odrv4 I__4253 (
            .O(N__21817),
            .I(\c0.n2080 ));
    CascadeMux I__4252 (
            .O(N__21814),
            .I(\c0.n2080_cascade_ ));
    InMux I__4251 (
            .O(N__21811),
            .I(N__21805));
    InMux I__4250 (
            .O(N__21810),
            .I(N__21805));
    LocalMux I__4249 (
            .O(N__21805),
            .I(\c0.n5243 ));
    CascadeMux I__4248 (
            .O(N__21802),
            .I(N__21799));
    InMux I__4247 (
            .O(N__21799),
            .I(N__21796));
    LocalMux I__4246 (
            .O(N__21796),
            .I(N__21793));
    Span4Mux_v I__4245 (
            .O(N__21793),
            .I(N__21790));
    Span4Mux_h I__4244 (
            .O(N__21790),
            .I(N__21787));
    Span4Mux_s2_h I__4243 (
            .O(N__21787),
            .I(N__21784));
    Odrv4 I__4242 (
            .O(N__21784),
            .I(\c0.n16_adj_1922 ));
    InMux I__4241 (
            .O(N__21781),
            .I(N__21778));
    LocalMux I__4240 (
            .O(N__21778),
            .I(\c0.n25_adj_1926 ));
    InMux I__4239 (
            .O(N__21775),
            .I(N__21772));
    LocalMux I__4238 (
            .O(N__21772),
            .I(N__21769));
    Span4Mux_s3_h I__4237 (
            .O(N__21769),
            .I(N__21766));
    Odrv4 I__4236 (
            .O(N__21766),
            .I(\c0.n5429 ));
    InMux I__4235 (
            .O(N__21763),
            .I(N__21760));
    LocalMux I__4234 (
            .O(N__21760),
            .I(N__21757));
    Span4Mux_v I__4233 (
            .O(N__21757),
            .I(N__21754));
    Odrv4 I__4232 (
            .O(N__21754),
            .I(\c0.n5791 ));
    InMux I__4231 (
            .O(N__21751),
            .I(N__21748));
    LocalMux I__4230 (
            .O(N__21748),
            .I(N__21745));
    Odrv12 I__4229 (
            .O(N__21745),
            .I(\c0.n5432 ));
    InMux I__4228 (
            .O(N__21742),
            .I(N__21739));
    LocalMux I__4227 (
            .O(N__21739),
            .I(N__21736));
    Span4Mux_h I__4226 (
            .O(N__21736),
            .I(N__21730));
    InMux I__4225 (
            .O(N__21735),
            .I(N__21727));
    InMux I__4224 (
            .O(N__21734),
            .I(N__21722));
    InMux I__4223 (
            .O(N__21733),
            .I(N__21722));
    Odrv4 I__4222 (
            .O(N__21730),
            .I(\c0.data_in_field_30 ));
    LocalMux I__4221 (
            .O(N__21727),
            .I(\c0.data_in_field_30 ));
    LocalMux I__4220 (
            .O(N__21722),
            .I(\c0.data_in_field_30 ));
    InMux I__4219 (
            .O(N__21715),
            .I(N__21712));
    LocalMux I__4218 (
            .O(N__21712),
            .I(N__21708));
    InMux I__4217 (
            .O(N__21711),
            .I(N__21704));
    Span4Mux_v I__4216 (
            .O(N__21708),
            .I(N__21701));
    InMux I__4215 (
            .O(N__21707),
            .I(N__21698));
    LocalMux I__4214 (
            .O(N__21704),
            .I(N__21695));
    Span4Mux_h I__4213 (
            .O(N__21701),
            .I(N__21692));
    LocalMux I__4212 (
            .O(N__21698),
            .I(N__21687));
    Span4Mux_v I__4211 (
            .O(N__21695),
            .I(N__21687));
    Odrv4 I__4210 (
            .O(N__21692),
            .I(\c0.data_in_field_13 ));
    Odrv4 I__4209 (
            .O(N__21687),
            .I(\c0.data_in_field_13 ));
    InMux I__4208 (
            .O(N__21682),
            .I(N__21679));
    LocalMux I__4207 (
            .O(N__21679),
            .I(N__21676));
    Span4Mux_s3_h I__4206 (
            .O(N__21676),
            .I(N__21673));
    Span4Mux_h I__4205 (
            .O(N__21673),
            .I(N__21670));
    Odrv4 I__4204 (
            .O(N__21670),
            .I(\c0.n5393 ));
    CascadeMux I__4203 (
            .O(N__21667),
            .I(N__21664));
    InMux I__4202 (
            .O(N__21664),
            .I(N__21660));
    InMux I__4201 (
            .O(N__21663),
            .I(N__21657));
    LocalMux I__4200 (
            .O(N__21660),
            .I(N__21652));
    LocalMux I__4199 (
            .O(N__21657),
            .I(N__21652));
    Span4Mux_v I__4198 (
            .O(N__21652),
            .I(N__21649));
    Span4Mux_h I__4197 (
            .O(N__21649),
            .I(N__21645));
    InMux I__4196 (
            .O(N__21648),
            .I(N__21642));
    Odrv4 I__4195 (
            .O(N__21645),
            .I(data_in_14_7));
    LocalMux I__4194 (
            .O(N__21642),
            .I(data_in_14_7));
    InMux I__4193 (
            .O(N__21637),
            .I(N__21634));
    LocalMux I__4192 (
            .O(N__21634),
            .I(\c0.n10_adj_1898 ));
    InMux I__4191 (
            .O(N__21631),
            .I(N__21628));
    LocalMux I__4190 (
            .O(N__21628),
            .I(N__21625));
    Span4Mux_s2_h I__4189 (
            .O(N__21625),
            .I(N__21621));
    InMux I__4188 (
            .O(N__21624),
            .I(N__21618));
    Span4Mux_h I__4187 (
            .O(N__21621),
            .I(N__21613));
    LocalMux I__4186 (
            .O(N__21618),
            .I(N__21610));
    InMux I__4185 (
            .O(N__21617),
            .I(N__21605));
    InMux I__4184 (
            .O(N__21616),
            .I(N__21605));
    Odrv4 I__4183 (
            .O(N__21613),
            .I(\c0.data_in_field_69 ));
    Odrv4 I__4182 (
            .O(N__21610),
            .I(\c0.data_in_field_69 ));
    LocalMux I__4181 (
            .O(N__21605),
            .I(\c0.data_in_field_69 ));
    InMux I__4180 (
            .O(N__21598),
            .I(N__21595));
    LocalMux I__4179 (
            .O(N__21595),
            .I(\c0.n5159 ));
    InMux I__4178 (
            .O(N__21592),
            .I(N__21589));
    LocalMux I__4177 (
            .O(N__21589),
            .I(N__21585));
    InMux I__4176 (
            .O(N__21588),
            .I(N__21582));
    Span4Mux_v I__4175 (
            .O(N__21585),
            .I(N__21574));
    LocalMux I__4174 (
            .O(N__21582),
            .I(N__21574));
    InMux I__4173 (
            .O(N__21581),
            .I(N__21569));
    InMux I__4172 (
            .O(N__21580),
            .I(N__21569));
    InMux I__4171 (
            .O(N__21579),
            .I(N__21566));
    Span4Mux_h I__4170 (
            .O(N__21574),
            .I(N__21563));
    LocalMux I__4169 (
            .O(N__21569),
            .I(\c0.data_in_field_99 ));
    LocalMux I__4168 (
            .O(N__21566),
            .I(\c0.data_in_field_99 ));
    Odrv4 I__4167 (
            .O(N__21563),
            .I(\c0.data_in_field_99 ));
    CascadeMux I__4166 (
            .O(N__21556),
            .I(\c0.n5159_cascade_ ));
    CascadeMux I__4165 (
            .O(N__21553),
            .I(\c0.n5683_cascade_ ));
    InMux I__4164 (
            .O(N__21550),
            .I(N__21547));
    LocalMux I__4163 (
            .O(N__21547),
            .I(\c0.n5695 ));
    CascadeMux I__4162 (
            .O(N__21544),
            .I(\c0.n5480_cascade_ ));
    InMux I__4161 (
            .O(N__21541),
            .I(N__21538));
    LocalMux I__4160 (
            .O(N__21538),
            .I(\c0.n5483 ));
    CascadeMux I__4159 (
            .O(N__21535),
            .I(\c0.n5677_cascade_ ));
    InMux I__4158 (
            .O(N__21532),
            .I(N__21529));
    LocalMux I__4157 (
            .O(N__21529),
            .I(N__21526));
    Odrv12 I__4156 (
            .O(N__21526),
            .I(\c0.n5680 ));
    InMux I__4155 (
            .O(N__21523),
            .I(N__21518));
    InMux I__4154 (
            .O(N__21522),
            .I(N__21514));
    InMux I__4153 (
            .O(N__21521),
            .I(N__21511));
    LocalMux I__4152 (
            .O(N__21518),
            .I(N__21508));
    InMux I__4151 (
            .O(N__21517),
            .I(N__21505));
    LocalMux I__4150 (
            .O(N__21514),
            .I(data_in_18_5));
    LocalMux I__4149 (
            .O(N__21511),
            .I(data_in_18_5));
    Odrv12 I__4148 (
            .O(N__21508),
            .I(data_in_18_5));
    LocalMux I__4147 (
            .O(N__21505),
            .I(data_in_18_5));
    InMux I__4146 (
            .O(N__21496),
            .I(N__21493));
    LocalMux I__4145 (
            .O(N__21493),
            .I(\c0.n24_adj_1895 ));
    InMux I__4144 (
            .O(N__21490),
            .I(N__21487));
    LocalMux I__4143 (
            .O(N__21487),
            .I(N__21484));
    Span4Mux_v I__4142 (
            .O(N__21484),
            .I(N__21481));
    Span4Mux_v I__4141 (
            .O(N__21481),
            .I(N__21477));
    CascadeMux I__4140 (
            .O(N__21480),
            .I(N__21474));
    Span4Mux_h I__4139 (
            .O(N__21477),
            .I(N__21471));
    InMux I__4138 (
            .O(N__21474),
            .I(N__21468));
    Odrv4 I__4137 (
            .O(N__21471),
            .I(rx_data_0));
    LocalMux I__4136 (
            .O(N__21468),
            .I(rx_data_0));
    InMux I__4135 (
            .O(N__21463),
            .I(N__21459));
    InMux I__4134 (
            .O(N__21462),
            .I(N__21456));
    LocalMux I__4133 (
            .O(N__21459),
            .I(N__21453));
    LocalMux I__4132 (
            .O(N__21456),
            .I(N__21450));
    Span4Mux_h I__4131 (
            .O(N__21453),
            .I(N__21447));
    Span12Mux_s7_v I__4130 (
            .O(N__21450),
            .I(N__21442));
    Span4Mux_v I__4129 (
            .O(N__21447),
            .I(N__21439));
    InMux I__4128 (
            .O(N__21446),
            .I(N__21434));
    InMux I__4127 (
            .O(N__21445),
            .I(N__21434));
    Odrv12 I__4126 (
            .O(N__21442),
            .I(data_in_19_0));
    Odrv4 I__4125 (
            .O(N__21439),
            .I(data_in_19_0));
    LocalMux I__4124 (
            .O(N__21434),
            .I(data_in_19_0));
    InMux I__4123 (
            .O(N__21427),
            .I(N__21424));
    LocalMux I__4122 (
            .O(N__21424),
            .I(N__21421));
    Odrv4 I__4121 (
            .O(N__21421),
            .I(\c0.n3567 ));
    InMux I__4120 (
            .O(N__21418),
            .I(N__21409));
    InMux I__4119 (
            .O(N__21417),
            .I(N__21404));
    InMux I__4118 (
            .O(N__21416),
            .I(N__21401));
    InMux I__4117 (
            .O(N__21415),
            .I(N__21398));
    InMux I__4116 (
            .O(N__21414),
            .I(N__21395));
    InMux I__4115 (
            .O(N__21413),
            .I(N__21392));
    InMux I__4114 (
            .O(N__21412),
            .I(N__21389));
    LocalMux I__4113 (
            .O(N__21409),
            .I(N__21386));
    InMux I__4112 (
            .O(N__21408),
            .I(N__21381));
    InMux I__4111 (
            .O(N__21407),
            .I(N__21381));
    LocalMux I__4110 (
            .O(N__21404),
            .I(N__21376));
    LocalMux I__4109 (
            .O(N__21401),
            .I(N__21367));
    LocalMux I__4108 (
            .O(N__21398),
            .I(N__21367));
    LocalMux I__4107 (
            .O(N__21395),
            .I(N__21367));
    LocalMux I__4106 (
            .O(N__21392),
            .I(N__21367));
    LocalMux I__4105 (
            .O(N__21389),
            .I(N__21364));
    Span4Mux_v I__4104 (
            .O(N__21386),
            .I(N__21361));
    LocalMux I__4103 (
            .O(N__21381),
            .I(N__21358));
    InMux I__4102 (
            .O(N__21380),
            .I(N__21353));
    InMux I__4101 (
            .O(N__21379),
            .I(N__21353));
    Span4Mux_v I__4100 (
            .O(N__21376),
            .I(N__21346));
    Span4Mux_v I__4099 (
            .O(N__21367),
            .I(N__21346));
    Span4Mux_h I__4098 (
            .O(N__21364),
            .I(N__21346));
    Span4Mux_h I__4097 (
            .O(N__21361),
            .I(N__21340));
    Span4Mux_v I__4096 (
            .O(N__21358),
            .I(N__21340));
    LocalMux I__4095 (
            .O(N__21353),
            .I(N__21335));
    Span4Mux_h I__4094 (
            .O(N__21346),
            .I(N__21335));
    InMux I__4093 (
            .O(N__21345),
            .I(N__21332));
    Odrv4 I__4092 (
            .O(N__21340),
            .I(\c0.byte_transmit_counter_3 ));
    Odrv4 I__4091 (
            .O(N__21335),
            .I(\c0.byte_transmit_counter_3 ));
    LocalMux I__4090 (
            .O(N__21332),
            .I(\c0.byte_transmit_counter_3 ));
    CascadeMux I__4089 (
            .O(N__21325),
            .I(\c0.n5523_cascade_ ));
    InMux I__4088 (
            .O(N__21322),
            .I(N__21315));
    InMux I__4087 (
            .O(N__21321),
            .I(N__21309));
    InMux I__4086 (
            .O(N__21320),
            .I(N__21306));
    InMux I__4085 (
            .O(N__21319),
            .I(N__21303));
    InMux I__4084 (
            .O(N__21318),
            .I(N__21300));
    LocalMux I__4083 (
            .O(N__21315),
            .I(N__21297));
    InMux I__4082 (
            .O(N__21314),
            .I(N__21294));
    InMux I__4081 (
            .O(N__21313),
            .I(N__21289));
    InMux I__4080 (
            .O(N__21312),
            .I(N__21289));
    LocalMux I__4079 (
            .O(N__21309),
            .I(N__21283));
    LocalMux I__4078 (
            .O(N__21306),
            .I(N__21283));
    LocalMux I__4077 (
            .O(N__21303),
            .I(N__21280));
    LocalMux I__4076 (
            .O(N__21300),
            .I(N__21275));
    Span4Mux_v I__4075 (
            .O(N__21297),
            .I(N__21275));
    LocalMux I__4074 (
            .O(N__21294),
            .I(N__21270));
    LocalMux I__4073 (
            .O(N__21289),
            .I(N__21270));
    InMux I__4072 (
            .O(N__21288),
            .I(N__21267));
    Span4Mux_v I__4071 (
            .O(N__21283),
            .I(N__21262));
    Span4Mux_h I__4070 (
            .O(N__21280),
            .I(N__21262));
    Span4Mux_h I__4069 (
            .O(N__21275),
            .I(N__21258));
    Span4Mux_v I__4068 (
            .O(N__21270),
            .I(N__21255));
    LocalMux I__4067 (
            .O(N__21267),
            .I(N__21250));
    Span4Mux_h I__4066 (
            .O(N__21262),
            .I(N__21250));
    InMux I__4065 (
            .O(N__21261),
            .I(N__21247));
    Odrv4 I__4064 (
            .O(N__21258),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__4063 (
            .O(N__21255),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__4062 (
            .O(N__21250),
            .I(\c0.byte_transmit_counter_2 ));
    LocalMux I__4061 (
            .O(N__21247),
            .I(\c0.byte_transmit_counter_2 ));
    CascadeMux I__4060 (
            .O(N__21238),
            .I(N__21235));
    InMux I__4059 (
            .O(N__21235),
            .I(N__21232));
    LocalMux I__4058 (
            .O(N__21232),
            .I(N__21227));
    InMux I__4057 (
            .O(N__21231),
            .I(N__21224));
    InMux I__4056 (
            .O(N__21230),
            .I(N__21221));
    Span4Mux_v I__4055 (
            .O(N__21227),
            .I(N__21218));
    LocalMux I__4054 (
            .O(N__21224),
            .I(N__21215));
    LocalMux I__4053 (
            .O(N__21221),
            .I(N__21212));
    Odrv4 I__4052 (
            .O(N__21218),
            .I(\c0.n1236 ));
    Odrv4 I__4051 (
            .O(N__21215),
            .I(\c0.n1236 ));
    Odrv4 I__4050 (
            .O(N__21212),
            .I(\c0.n1236 ));
    InMux I__4049 (
            .O(N__21205),
            .I(N__21202));
    LocalMux I__4048 (
            .O(N__21202),
            .I(\c0.n5515 ));
    CascadeMux I__4047 (
            .O(N__21199),
            .I(\c0.n5513_cascade_ ));
    InMux I__4046 (
            .O(N__21196),
            .I(N__21192));
    InMux I__4045 (
            .O(N__21195),
            .I(N__21183));
    LocalMux I__4044 (
            .O(N__21192),
            .I(N__21180));
    InMux I__4043 (
            .O(N__21191),
            .I(N__21177));
    InMux I__4042 (
            .O(N__21190),
            .I(N__21174));
    InMux I__4041 (
            .O(N__21189),
            .I(N__21169));
    InMux I__4040 (
            .O(N__21188),
            .I(N__21169));
    InMux I__4039 (
            .O(N__21187),
            .I(N__21166));
    InMux I__4038 (
            .O(N__21186),
            .I(N__21163));
    LocalMux I__4037 (
            .O(N__21183),
            .I(N__21160));
    Span4Mux_h I__4036 (
            .O(N__21180),
            .I(N__21149));
    LocalMux I__4035 (
            .O(N__21177),
            .I(N__21149));
    LocalMux I__4034 (
            .O(N__21174),
            .I(N__21149));
    LocalMux I__4033 (
            .O(N__21169),
            .I(N__21149));
    LocalMux I__4032 (
            .O(N__21166),
            .I(N__21149));
    LocalMux I__4031 (
            .O(N__21163),
            .I(N__21143));
    Span4Mux_h I__4030 (
            .O(N__21160),
            .I(N__21143));
    Span4Mux_v I__4029 (
            .O(N__21149),
            .I(N__21140));
    InMux I__4028 (
            .O(N__21148),
            .I(N__21137));
    Odrv4 I__4027 (
            .O(N__21143),
            .I(\c0.byte_transmit_counter_4 ));
    Odrv4 I__4026 (
            .O(N__21140),
            .I(\c0.byte_transmit_counter_4 ));
    LocalMux I__4025 (
            .O(N__21137),
            .I(\c0.byte_transmit_counter_4 ));
    InMux I__4024 (
            .O(N__21130),
            .I(N__21127));
    LocalMux I__4023 (
            .O(N__21127),
            .I(tx_data_6_N_keep));
    InMux I__4022 (
            .O(N__21124),
            .I(N__21120));
    InMux I__4021 (
            .O(N__21123),
            .I(N__21116));
    LocalMux I__4020 (
            .O(N__21120),
            .I(N__21113));
    InMux I__4019 (
            .O(N__21119),
            .I(N__21110));
    LocalMux I__4018 (
            .O(N__21116),
            .I(N__21105));
    Span4Mux_v I__4017 (
            .O(N__21113),
            .I(N__21100));
    LocalMux I__4016 (
            .O(N__21110),
            .I(N__21100));
    InMux I__4015 (
            .O(N__21109),
            .I(N__21097));
    InMux I__4014 (
            .O(N__21108),
            .I(N__21094));
    Span4Mux_v I__4013 (
            .O(N__21105),
            .I(N__21091));
    Span4Mux_h I__4012 (
            .O(N__21100),
            .I(N__21088));
    LocalMux I__4011 (
            .O(N__21097),
            .I(data_out_10_5));
    LocalMux I__4010 (
            .O(N__21094),
            .I(data_out_10_5));
    Odrv4 I__4009 (
            .O(N__21091),
            .I(data_out_10_5));
    Odrv4 I__4008 (
            .O(N__21088),
            .I(data_out_10_5));
    InMux I__4007 (
            .O(N__21079),
            .I(N__21072));
    InMux I__4006 (
            .O(N__21078),
            .I(N__21069));
    InMux I__4005 (
            .O(N__21077),
            .I(N__21066));
    InMux I__4004 (
            .O(N__21076),
            .I(N__21063));
    InMux I__4003 (
            .O(N__21075),
            .I(N__21060));
    LocalMux I__4002 (
            .O(N__21072),
            .I(N__21056));
    LocalMux I__4001 (
            .O(N__21069),
            .I(N__21053));
    LocalMux I__4000 (
            .O(N__21066),
            .I(N__21050));
    LocalMux I__3999 (
            .O(N__21063),
            .I(N__21045));
    LocalMux I__3998 (
            .O(N__21060),
            .I(N__21045));
    InMux I__3997 (
            .O(N__21059),
            .I(N__21041));
    Span4Mux_v I__3996 (
            .O(N__21056),
            .I(N__21038));
    Span4Mux_h I__3995 (
            .O(N__21053),
            .I(N__21035));
    Span4Mux_v I__3994 (
            .O(N__21050),
            .I(N__21030));
    Span4Mux_h I__3993 (
            .O(N__21045),
            .I(N__21030));
    InMux I__3992 (
            .O(N__21044),
            .I(N__21027));
    LocalMux I__3991 (
            .O(N__21041),
            .I(data_out_10_1));
    Odrv4 I__3990 (
            .O(N__21038),
            .I(data_out_10_1));
    Odrv4 I__3989 (
            .O(N__21035),
            .I(data_out_10_1));
    Odrv4 I__3988 (
            .O(N__21030),
            .I(data_out_10_1));
    LocalMux I__3987 (
            .O(N__21027),
            .I(data_out_10_1));
    InMux I__3986 (
            .O(N__21016),
            .I(N__21013));
    LocalMux I__3985 (
            .O(N__21013),
            .I(N__21009));
    InMux I__3984 (
            .O(N__21012),
            .I(N__21003));
    Span4Mux_v I__3983 (
            .O(N__21009),
            .I(N__21000));
    InMux I__3982 (
            .O(N__21008),
            .I(N__20995));
    InMux I__3981 (
            .O(N__21007),
            .I(N__20995));
    InMux I__3980 (
            .O(N__21006),
            .I(N__20992));
    LocalMux I__3979 (
            .O(N__21003),
            .I(data_out_10_3));
    Odrv4 I__3978 (
            .O(N__21000),
            .I(data_out_10_3));
    LocalMux I__3977 (
            .O(N__20995),
            .I(data_out_10_3));
    LocalMux I__3976 (
            .O(N__20992),
            .I(data_out_10_3));
    CascadeMux I__3975 (
            .O(N__20983),
            .I(N__20980));
    InMux I__3974 (
            .O(N__20980),
            .I(N__20976));
    InMux I__3973 (
            .O(N__20979),
            .I(N__20973));
    LocalMux I__3972 (
            .O(N__20976),
            .I(N__20970));
    LocalMux I__3971 (
            .O(N__20973),
            .I(N__20967));
    Span4Mux_v I__3970 (
            .O(N__20970),
            .I(N__20962));
    Span4Mux_s3_h I__3969 (
            .O(N__20967),
            .I(N__20962));
    Span4Mux_v I__3968 (
            .O(N__20962),
            .I(N__20959));
    Odrv4 I__3967 (
            .O(N__20959),
            .I(n5132));
    CascadeMux I__3966 (
            .O(N__20956),
            .I(\c0.n5839_cascade_ ));
    CascadeMux I__3965 (
            .O(N__20953),
            .I(\c0.n5833_cascade_ ));
    CascadeMux I__3964 (
            .O(N__20950),
            .I(\c0.n5417_cascade_ ));
    InMux I__3963 (
            .O(N__20947),
            .I(N__20944));
    LocalMux I__3962 (
            .O(N__20944),
            .I(\c0.n5414 ));
    InMux I__3961 (
            .O(N__20941),
            .I(N__20938));
    LocalMux I__3960 (
            .O(N__20938),
            .I(\c0.n5827 ));
    InMux I__3959 (
            .O(N__20935),
            .I(N__20927));
    InMux I__3958 (
            .O(N__20934),
            .I(N__20922));
    InMux I__3957 (
            .O(N__20933),
            .I(N__20922));
    InMux I__3956 (
            .O(N__20932),
            .I(N__20917));
    InMux I__3955 (
            .O(N__20931),
            .I(N__20917));
    CascadeMux I__3954 (
            .O(N__20930),
            .I(N__20912));
    LocalMux I__3953 (
            .O(N__20927),
            .I(N__20908));
    LocalMux I__3952 (
            .O(N__20922),
            .I(N__20903));
    LocalMux I__3951 (
            .O(N__20917),
            .I(N__20903));
    InMux I__3950 (
            .O(N__20916),
            .I(N__20900));
    CascadeMux I__3949 (
            .O(N__20915),
            .I(N__20895));
    InMux I__3948 (
            .O(N__20912),
            .I(N__20892));
    InMux I__3947 (
            .O(N__20911),
            .I(N__20889));
    Sp12to4 I__3946 (
            .O(N__20908),
            .I(N__20882));
    Sp12to4 I__3945 (
            .O(N__20903),
            .I(N__20882));
    LocalMux I__3944 (
            .O(N__20900),
            .I(N__20882));
    InMux I__3943 (
            .O(N__20899),
            .I(N__20877));
    InMux I__3942 (
            .O(N__20898),
            .I(N__20877));
    InMux I__3941 (
            .O(N__20895),
            .I(N__20874));
    LocalMux I__3940 (
            .O(N__20892),
            .I(r_Rx_Data));
    LocalMux I__3939 (
            .O(N__20889),
            .I(r_Rx_Data));
    Odrv12 I__3938 (
            .O(N__20882),
            .I(r_Rx_Data));
    LocalMux I__3937 (
            .O(N__20877),
            .I(r_Rx_Data));
    LocalMux I__3936 (
            .O(N__20874),
            .I(r_Rx_Data));
    CascadeMux I__3935 (
            .O(N__20863),
            .I(N__20860));
    InMux I__3934 (
            .O(N__20860),
            .I(N__20854));
    InMux I__3933 (
            .O(N__20859),
            .I(N__20854));
    LocalMux I__3932 (
            .O(N__20854),
            .I(N__20851));
    Span4Mux_v I__3931 (
            .O(N__20851),
            .I(N__20847));
    InMux I__3930 (
            .O(N__20850),
            .I(N__20844));
    Odrv4 I__3929 (
            .O(N__20847),
            .I(n1714));
    LocalMux I__3928 (
            .O(N__20844),
            .I(n1714));
    InMux I__3927 (
            .O(N__20839),
            .I(N__20836));
    LocalMux I__3926 (
            .O(N__20836),
            .I(N__20832));
    InMux I__3925 (
            .O(N__20835),
            .I(N__20829));
    Odrv4 I__3924 (
            .O(N__20832),
            .I(n3342));
    LocalMux I__3923 (
            .O(N__20829),
            .I(n3342));
    CascadeMux I__3922 (
            .O(N__20824),
            .I(N__20821));
    InMux I__3921 (
            .O(N__20821),
            .I(N__20815));
    InMux I__3920 (
            .O(N__20820),
            .I(N__20815));
    LocalMux I__3919 (
            .O(N__20815),
            .I(rx_data_7));
    InMux I__3918 (
            .O(N__20812),
            .I(N__20808));
    InMux I__3917 (
            .O(N__20811),
            .I(N__20805));
    LocalMux I__3916 (
            .O(N__20808),
            .I(N__20802));
    LocalMux I__3915 (
            .O(N__20805),
            .I(N__20799));
    Span4Mux_h I__3914 (
            .O(N__20802),
            .I(N__20793));
    Span4Mux_s1_v I__3913 (
            .O(N__20799),
            .I(N__20793));
    InMux I__3912 (
            .O(N__20798),
            .I(N__20790));
    Odrv4 I__3911 (
            .O(N__20793),
            .I(data_in_17_1));
    LocalMux I__3910 (
            .O(N__20790),
            .I(data_in_17_1));
    InMux I__3909 (
            .O(N__20785),
            .I(N__20781));
    InMux I__3908 (
            .O(N__20784),
            .I(N__20778));
    LocalMux I__3907 (
            .O(N__20781),
            .I(N__20775));
    LocalMux I__3906 (
            .O(N__20778),
            .I(data_out_19_6));
    Odrv4 I__3905 (
            .O(N__20775),
            .I(data_out_19_6));
    CascadeMux I__3904 (
            .O(N__20770),
            .I(N__20767));
    InMux I__3903 (
            .O(N__20767),
            .I(N__20764));
    LocalMux I__3902 (
            .O(N__20764),
            .I(N__20760));
    InMux I__3901 (
            .O(N__20763),
            .I(N__20757));
    Span4Mux_h I__3900 (
            .O(N__20760),
            .I(N__20754));
    LocalMux I__3899 (
            .O(N__20757),
            .I(data_out_18_6));
    Odrv4 I__3898 (
            .O(N__20754),
            .I(data_out_18_6));
    InMux I__3897 (
            .O(N__20749),
            .I(N__20745));
    InMux I__3896 (
            .O(N__20748),
            .I(N__20740));
    LocalMux I__3895 (
            .O(N__20745),
            .I(N__20736));
    InMux I__3894 (
            .O(N__20744),
            .I(N__20731));
    InMux I__3893 (
            .O(N__20743),
            .I(N__20731));
    LocalMux I__3892 (
            .O(N__20740),
            .I(N__20727));
    InMux I__3891 (
            .O(N__20739),
            .I(N__20724));
    Span4Mux_v I__3890 (
            .O(N__20736),
            .I(N__20719));
    LocalMux I__3889 (
            .O(N__20731),
            .I(N__20719));
    InMux I__3888 (
            .O(N__20730),
            .I(N__20715));
    Span4Mux_v I__3887 (
            .O(N__20727),
            .I(N__20712));
    LocalMux I__3886 (
            .O(N__20724),
            .I(N__20709));
    Span4Mux_h I__3885 (
            .O(N__20719),
            .I(N__20706));
    InMux I__3884 (
            .O(N__20718),
            .I(N__20703));
    LocalMux I__3883 (
            .O(N__20715),
            .I(data_out_11_5));
    Odrv4 I__3882 (
            .O(N__20712),
            .I(data_out_11_5));
    Odrv4 I__3881 (
            .O(N__20709),
            .I(data_out_11_5));
    Odrv4 I__3880 (
            .O(N__20706),
            .I(data_out_11_5));
    LocalMux I__3879 (
            .O(N__20703),
            .I(data_out_11_5));
    InMux I__3878 (
            .O(N__20692),
            .I(N__20689));
    LocalMux I__3877 (
            .O(N__20689),
            .I(N__20686));
    Odrv4 I__3876 (
            .O(N__20686),
            .I(n5176));
    InMux I__3875 (
            .O(N__20683),
            .I(N__20680));
    LocalMux I__3874 (
            .O(N__20680),
            .I(N__20674));
    InMux I__3873 (
            .O(N__20679),
            .I(N__20671));
    InMux I__3872 (
            .O(N__20678),
            .I(N__20668));
    InMux I__3871 (
            .O(N__20677),
            .I(N__20665));
    Span4Mux_v I__3870 (
            .O(N__20674),
            .I(N__20658));
    LocalMux I__3869 (
            .O(N__20671),
            .I(N__20658));
    LocalMux I__3868 (
            .O(N__20668),
            .I(N__20658));
    LocalMux I__3867 (
            .O(N__20665),
            .I(N__20655));
    Span4Mux_h I__3866 (
            .O(N__20658),
            .I(N__20652));
    Odrv4 I__3865 (
            .O(N__20655),
            .I(\c0.n1590 ));
    Odrv4 I__3864 (
            .O(N__20652),
            .I(\c0.n1590 ));
    InMux I__3863 (
            .O(N__20647),
            .I(N__20644));
    LocalMux I__3862 (
            .O(N__20644),
            .I(N__20635));
    InMux I__3861 (
            .O(N__20643),
            .I(N__20632));
    InMux I__3860 (
            .O(N__20642),
            .I(N__20627));
    InMux I__3859 (
            .O(N__20641),
            .I(N__20627));
    CascadeMux I__3858 (
            .O(N__20640),
            .I(N__20624));
    InMux I__3857 (
            .O(N__20639),
            .I(N__20621));
    InMux I__3856 (
            .O(N__20638),
            .I(N__20618));
    Span4Mux_v I__3855 (
            .O(N__20635),
            .I(N__20611));
    LocalMux I__3854 (
            .O(N__20632),
            .I(N__20611));
    LocalMux I__3853 (
            .O(N__20627),
            .I(N__20611));
    InMux I__3852 (
            .O(N__20624),
            .I(N__20607));
    LocalMux I__3851 (
            .O(N__20621),
            .I(N__20604));
    LocalMux I__3850 (
            .O(N__20618),
            .I(N__20599));
    Span4Mux_h I__3849 (
            .O(N__20611),
            .I(N__20599));
    InMux I__3848 (
            .O(N__20610),
            .I(N__20596));
    LocalMux I__3847 (
            .O(N__20607),
            .I(data_out_11_6));
    Odrv4 I__3846 (
            .O(N__20604),
            .I(data_out_11_6));
    Odrv4 I__3845 (
            .O(N__20599),
            .I(data_out_11_6));
    LocalMux I__3844 (
            .O(N__20596),
            .I(data_out_11_6));
    InMux I__3843 (
            .O(N__20587),
            .I(N__20576));
    InMux I__3842 (
            .O(N__20586),
            .I(N__20573));
    InMux I__3841 (
            .O(N__20585),
            .I(N__20568));
    InMux I__3840 (
            .O(N__20584),
            .I(N__20565));
    InMux I__3839 (
            .O(N__20583),
            .I(N__20562));
    InMux I__3838 (
            .O(N__20582),
            .I(N__20557));
    InMux I__3837 (
            .O(N__20581),
            .I(N__20557));
    InMux I__3836 (
            .O(N__20580),
            .I(N__20554));
    InMux I__3835 (
            .O(N__20579),
            .I(N__20551));
    LocalMux I__3834 (
            .O(N__20576),
            .I(N__20548));
    LocalMux I__3833 (
            .O(N__20573),
            .I(N__20545));
    InMux I__3832 (
            .O(N__20572),
            .I(N__20540));
    InMux I__3831 (
            .O(N__20571),
            .I(N__20540));
    LocalMux I__3830 (
            .O(N__20568),
            .I(N__20531));
    LocalMux I__3829 (
            .O(N__20565),
            .I(N__20531));
    LocalMux I__3828 (
            .O(N__20562),
            .I(N__20531));
    LocalMux I__3827 (
            .O(N__20557),
            .I(N__20531));
    LocalMux I__3826 (
            .O(N__20554),
            .I(N__20525));
    LocalMux I__3825 (
            .O(N__20551),
            .I(N__20525));
    Span4Mux_v I__3824 (
            .O(N__20548),
            .I(N__20518));
    Span4Mux_v I__3823 (
            .O(N__20545),
            .I(N__20518));
    LocalMux I__3822 (
            .O(N__20540),
            .I(N__20518));
    Span4Mux_v I__3821 (
            .O(N__20531),
            .I(N__20515));
    InMux I__3820 (
            .O(N__20530),
            .I(N__20512));
    Span4Mux_v I__3819 (
            .O(N__20525),
            .I(N__20505));
    Span4Mux_h I__3818 (
            .O(N__20518),
            .I(N__20502));
    Sp12to4 I__3817 (
            .O(N__20515),
            .I(N__20497));
    LocalMux I__3816 (
            .O(N__20512),
            .I(N__20497));
    InMux I__3815 (
            .O(N__20511),
            .I(N__20490));
    InMux I__3814 (
            .O(N__20510),
            .I(N__20490));
    InMux I__3813 (
            .O(N__20509),
            .I(N__20490));
    InMux I__3812 (
            .O(N__20508),
            .I(N__20487));
    Odrv4 I__3811 (
            .O(N__20505),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__3810 (
            .O(N__20502),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv12 I__3809 (
            .O(N__20497),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__3808 (
            .O(N__20490),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__3807 (
            .O(N__20487),
            .I(\c0.byte_transmit_counter_1 ));
    CascadeMux I__3806 (
            .O(N__20476),
            .I(N__20472));
    InMux I__3805 (
            .O(N__20475),
            .I(N__20463));
    InMux I__3804 (
            .O(N__20472),
            .I(N__20463));
    InMux I__3803 (
            .O(N__20471),
            .I(N__20460));
    InMux I__3802 (
            .O(N__20470),
            .I(N__20456));
    CascadeMux I__3801 (
            .O(N__20469),
            .I(N__20453));
    InMux I__3800 (
            .O(N__20468),
            .I(N__20450));
    LocalMux I__3799 (
            .O(N__20463),
            .I(N__20447));
    LocalMux I__3798 (
            .O(N__20460),
            .I(N__20444));
    InMux I__3797 (
            .O(N__20459),
            .I(N__20441));
    LocalMux I__3796 (
            .O(N__20456),
            .I(N__20438));
    InMux I__3795 (
            .O(N__20453),
            .I(N__20435));
    LocalMux I__3794 (
            .O(N__20450),
            .I(N__20432));
    Span4Mux_h I__3793 (
            .O(N__20447),
            .I(N__20427));
    Span4Mux_v I__3792 (
            .O(N__20444),
            .I(N__20427));
    LocalMux I__3791 (
            .O(N__20441),
            .I(data_out_10_6));
    Odrv12 I__3790 (
            .O(N__20438),
            .I(data_out_10_6));
    LocalMux I__3789 (
            .O(N__20435),
            .I(data_out_10_6));
    Odrv4 I__3788 (
            .O(N__20432),
            .I(data_out_10_6));
    Odrv4 I__3787 (
            .O(N__20427),
            .I(data_out_10_6));
    InMux I__3786 (
            .O(N__20416),
            .I(N__20400));
    InMux I__3785 (
            .O(N__20415),
            .I(N__20397));
    InMux I__3784 (
            .O(N__20414),
            .I(N__20394));
    InMux I__3783 (
            .O(N__20413),
            .I(N__20388));
    InMux I__3782 (
            .O(N__20412),
            .I(N__20385));
    InMux I__3781 (
            .O(N__20411),
            .I(N__20380));
    InMux I__3780 (
            .O(N__20410),
            .I(N__20380));
    InMux I__3779 (
            .O(N__20409),
            .I(N__20373));
    InMux I__3778 (
            .O(N__20408),
            .I(N__20373));
    InMux I__3777 (
            .O(N__20407),
            .I(N__20373));
    InMux I__3776 (
            .O(N__20406),
            .I(N__20368));
    InMux I__3775 (
            .O(N__20405),
            .I(N__20368));
    InMux I__3774 (
            .O(N__20404),
            .I(N__20363));
    InMux I__3773 (
            .O(N__20403),
            .I(N__20363));
    LocalMux I__3772 (
            .O(N__20400),
            .I(N__20356));
    LocalMux I__3771 (
            .O(N__20397),
            .I(N__20356));
    LocalMux I__3770 (
            .O(N__20394),
            .I(N__20356));
    InMux I__3769 (
            .O(N__20393),
            .I(N__20351));
    InMux I__3768 (
            .O(N__20392),
            .I(N__20348));
    InMux I__3767 (
            .O(N__20391),
            .I(N__20345));
    LocalMux I__3766 (
            .O(N__20388),
            .I(N__20334));
    LocalMux I__3765 (
            .O(N__20385),
            .I(N__20334));
    LocalMux I__3764 (
            .O(N__20380),
            .I(N__20334));
    LocalMux I__3763 (
            .O(N__20373),
            .I(N__20334));
    LocalMux I__3762 (
            .O(N__20368),
            .I(N__20334));
    LocalMux I__3761 (
            .O(N__20363),
            .I(N__20329));
    Span4Mux_v I__3760 (
            .O(N__20356),
            .I(N__20329));
    InMux I__3759 (
            .O(N__20355),
            .I(N__20326));
    CascadeMux I__3758 (
            .O(N__20354),
            .I(N__20321));
    LocalMux I__3757 (
            .O(N__20351),
            .I(N__20318));
    LocalMux I__3756 (
            .O(N__20348),
            .I(N__20315));
    LocalMux I__3755 (
            .O(N__20345),
            .I(N__20310));
    Span4Mux_v I__3754 (
            .O(N__20334),
            .I(N__20310));
    Sp12to4 I__3753 (
            .O(N__20329),
            .I(N__20305));
    LocalMux I__3752 (
            .O(N__20326),
            .I(N__20305));
    InMux I__3751 (
            .O(N__20325),
            .I(N__20300));
    InMux I__3750 (
            .O(N__20324),
            .I(N__20300));
    InMux I__3749 (
            .O(N__20321),
            .I(N__20297));
    Odrv4 I__3748 (
            .O(N__20318),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__3747 (
            .O(N__20315),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__3746 (
            .O(N__20310),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv12 I__3745 (
            .O(N__20305),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__3744 (
            .O(N__20300),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__3743 (
            .O(N__20297),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__3742 (
            .O(N__20284),
            .I(N__20281));
    LocalMux I__3741 (
            .O(N__20281),
            .I(N__20278));
    Span4Mux_v I__3740 (
            .O(N__20278),
            .I(N__20275));
    Odrv4 I__3739 (
            .O(N__20275),
            .I(\c0.n6_adj_1877 ));
    InMux I__3738 (
            .O(N__20272),
            .I(N__20269));
    LocalMux I__3737 (
            .O(N__20269),
            .I(N__20266));
    Span4Mux_v I__3736 (
            .O(N__20266),
            .I(N__20260));
    InMux I__3735 (
            .O(N__20265),
            .I(N__20253));
    InMux I__3734 (
            .O(N__20264),
            .I(N__20253));
    InMux I__3733 (
            .O(N__20263),
            .I(N__20253));
    Odrv4 I__3732 (
            .O(N__20260),
            .I(\c0.data_in_field_31 ));
    LocalMux I__3731 (
            .O(N__20253),
            .I(\c0.data_in_field_31 ));
    InMux I__3730 (
            .O(N__20248),
            .I(N__20245));
    LocalMux I__3729 (
            .O(N__20245),
            .I(\c0.n28_adj_1886 ));
    CascadeMux I__3728 (
            .O(N__20242),
            .I(N__20239));
    InMux I__3727 (
            .O(N__20239),
            .I(N__20236));
    LocalMux I__3726 (
            .O(N__20236),
            .I(N__20233));
    Span4Mux_h I__3725 (
            .O(N__20233),
            .I(N__20230));
    Odrv4 I__3724 (
            .O(N__20230),
            .I(\c0.n5222 ));
    InMux I__3723 (
            .O(N__20227),
            .I(N__20224));
    LocalMux I__3722 (
            .O(N__20224),
            .I(N__20221));
    Odrv4 I__3721 (
            .O(N__20221),
            .I(\c0.n34 ));
    InMux I__3720 (
            .O(N__20218),
            .I(N__20214));
    InMux I__3719 (
            .O(N__20217),
            .I(N__20211));
    LocalMux I__3718 (
            .O(N__20214),
            .I(N__20208));
    LocalMux I__3717 (
            .O(N__20211),
            .I(N__20204));
    Sp12to4 I__3716 (
            .O(N__20208),
            .I(N__20201));
    InMux I__3715 (
            .O(N__20207),
            .I(N__20198));
    Odrv4 I__3714 (
            .O(N__20204),
            .I(data_in_15_5));
    Odrv12 I__3713 (
            .O(N__20201),
            .I(data_in_15_5));
    LocalMux I__3712 (
            .O(N__20198),
            .I(data_in_15_5));
    CascadeMux I__3711 (
            .O(N__20191),
            .I(\c0.n1686_cascade_ ));
    InMux I__3710 (
            .O(N__20188),
            .I(N__20182));
    InMux I__3709 (
            .O(N__20187),
            .I(N__20179));
    InMux I__3708 (
            .O(N__20186),
            .I(N__20176));
    InMux I__3707 (
            .O(N__20185),
            .I(N__20173));
    LocalMux I__3706 (
            .O(N__20182),
            .I(\c0.data_in_field_25 ));
    LocalMux I__3705 (
            .O(N__20179),
            .I(\c0.data_in_field_25 ));
    LocalMux I__3704 (
            .O(N__20176),
            .I(\c0.data_in_field_25 ));
    LocalMux I__3703 (
            .O(N__20173),
            .I(\c0.data_in_field_25 ));
    InMux I__3702 (
            .O(N__20164),
            .I(N__20160));
    InMux I__3701 (
            .O(N__20163),
            .I(N__20156));
    LocalMux I__3700 (
            .O(N__20160),
            .I(N__20153));
    InMux I__3699 (
            .O(N__20159),
            .I(N__20150));
    LocalMux I__3698 (
            .O(N__20156),
            .I(N__20146));
    Span4Mux_v I__3697 (
            .O(N__20153),
            .I(N__20143));
    LocalMux I__3696 (
            .O(N__20150),
            .I(N__20140));
    InMux I__3695 (
            .O(N__20149),
            .I(N__20137));
    Span4Mux_h I__3694 (
            .O(N__20146),
            .I(N__20134));
    Span4Mux_h I__3693 (
            .O(N__20143),
            .I(N__20131));
    Span4Mux_v I__3692 (
            .O(N__20140),
            .I(N__20124));
    LocalMux I__3691 (
            .O(N__20137),
            .I(N__20124));
    Span4Mux_v I__3690 (
            .O(N__20134),
            .I(N__20124));
    Odrv4 I__3689 (
            .O(N__20131),
            .I(data_in_19_7));
    Odrv4 I__3688 (
            .O(N__20124),
            .I(data_in_19_7));
    InMux I__3687 (
            .O(N__20119),
            .I(N__20116));
    LocalMux I__3686 (
            .O(N__20116),
            .I(N__20112));
    CascadeMux I__3685 (
            .O(N__20115),
            .I(N__20109));
    Span4Mux_h I__3684 (
            .O(N__20112),
            .I(N__20106));
    InMux I__3683 (
            .O(N__20109),
            .I(N__20102));
    Span4Mux_v I__3682 (
            .O(N__20106),
            .I(N__20099));
    InMux I__3681 (
            .O(N__20105),
            .I(N__20096));
    LocalMux I__3680 (
            .O(N__20102),
            .I(\c0.data_in_field_7 ));
    Odrv4 I__3679 (
            .O(N__20099),
            .I(\c0.data_in_field_7 ));
    LocalMux I__3678 (
            .O(N__20096),
            .I(\c0.data_in_field_7 ));
    CascadeMux I__3677 (
            .O(N__20089),
            .I(\c0.n5162_cascade_ ));
    InMux I__3676 (
            .O(N__20086),
            .I(N__20081));
    InMux I__3675 (
            .O(N__20085),
            .I(N__20078));
    InMux I__3674 (
            .O(N__20084),
            .I(N__20075));
    LocalMux I__3673 (
            .O(N__20081),
            .I(N__20072));
    LocalMux I__3672 (
            .O(N__20078),
            .I(N__20068));
    LocalMux I__3671 (
            .O(N__20075),
            .I(N__20063));
    Span4Mux_v I__3670 (
            .O(N__20072),
            .I(N__20063));
    InMux I__3669 (
            .O(N__20071),
            .I(N__20060));
    Odrv4 I__3668 (
            .O(N__20068),
            .I(data_in_18_1));
    Odrv4 I__3667 (
            .O(N__20063),
            .I(data_in_18_1));
    LocalMux I__3666 (
            .O(N__20060),
            .I(data_in_18_1));
    CascadeMux I__3665 (
            .O(N__20053),
            .I(\c0.n1825_cascade_ ));
    InMux I__3664 (
            .O(N__20050),
            .I(N__20047));
    LocalMux I__3663 (
            .O(N__20047),
            .I(N__20044));
    Span4Mux_h I__3662 (
            .O(N__20044),
            .I(N__20037));
    InMux I__3661 (
            .O(N__20043),
            .I(N__20034));
    InMux I__3660 (
            .O(N__20042),
            .I(N__20031));
    InMux I__3659 (
            .O(N__20041),
            .I(N__20026));
    InMux I__3658 (
            .O(N__20040),
            .I(N__20026));
    Odrv4 I__3657 (
            .O(N__20037),
            .I(\c0.data_in_field_133 ));
    LocalMux I__3656 (
            .O(N__20034),
            .I(\c0.data_in_field_133 ));
    LocalMux I__3655 (
            .O(N__20031),
            .I(\c0.data_in_field_133 ));
    LocalMux I__3654 (
            .O(N__20026),
            .I(\c0.data_in_field_133 ));
    InMux I__3653 (
            .O(N__20017),
            .I(N__20014));
    LocalMux I__3652 (
            .O(N__20014),
            .I(N__20009));
    InMux I__3651 (
            .O(N__20013),
            .I(N__20006));
    InMux I__3650 (
            .O(N__20012),
            .I(N__20002));
    Span4Mux_h I__3649 (
            .O(N__20009),
            .I(N__19999));
    LocalMux I__3648 (
            .O(N__20006),
            .I(N__19996));
    InMux I__3647 (
            .O(N__20005),
            .I(N__19993));
    LocalMux I__3646 (
            .O(N__20002),
            .I(\c0.data_in_field_73 ));
    Odrv4 I__3645 (
            .O(N__19999),
            .I(\c0.data_in_field_73 ));
    Odrv12 I__3644 (
            .O(N__19996),
            .I(\c0.data_in_field_73 ));
    LocalMux I__3643 (
            .O(N__19993),
            .I(\c0.data_in_field_73 ));
    InMux I__3642 (
            .O(N__19984),
            .I(N__19980));
    CascadeMux I__3641 (
            .O(N__19983),
            .I(N__19976));
    LocalMux I__3640 (
            .O(N__19980),
            .I(N__19973));
    CascadeMux I__3639 (
            .O(N__19979),
            .I(N__19970));
    InMux I__3638 (
            .O(N__19976),
            .I(N__19966));
    Span4Mux_h I__3637 (
            .O(N__19973),
            .I(N__19963));
    InMux I__3636 (
            .O(N__19970),
            .I(N__19958));
    InMux I__3635 (
            .O(N__19969),
            .I(N__19958));
    LocalMux I__3634 (
            .O(N__19966),
            .I(\c0.data_in_field_35 ));
    Odrv4 I__3633 (
            .O(N__19963),
            .I(\c0.data_in_field_35 ));
    LocalMux I__3632 (
            .O(N__19958),
            .I(\c0.data_in_field_35 ));
    InMux I__3631 (
            .O(N__19951),
            .I(N__19948));
    LocalMux I__3630 (
            .O(N__19948),
            .I(N__19945));
    Span4Mux_v I__3629 (
            .O(N__19945),
            .I(N__19942));
    Odrv4 I__3628 (
            .O(N__19942),
            .I(\c0.n18 ));
    InMux I__3627 (
            .O(N__19939),
            .I(N__19936));
    LocalMux I__3626 (
            .O(N__19936),
            .I(N__19932));
    InMux I__3625 (
            .O(N__19935),
            .I(N__19929));
    Span4Mux_s2_h I__3624 (
            .O(N__19932),
            .I(N__19924));
    LocalMux I__3623 (
            .O(N__19929),
            .I(N__19924));
    Span4Mux_h I__3622 (
            .O(N__19924),
            .I(N__19919));
    InMux I__3621 (
            .O(N__19923),
            .I(N__19914));
    InMux I__3620 (
            .O(N__19922),
            .I(N__19914));
    Odrv4 I__3619 (
            .O(N__19919),
            .I(\c0.data_in_field_137 ));
    LocalMux I__3618 (
            .O(N__19914),
            .I(\c0.data_in_field_137 ));
    CascadeMux I__3617 (
            .O(N__19909),
            .I(N__19906));
    InMux I__3616 (
            .O(N__19906),
            .I(N__19900));
    InMux I__3615 (
            .O(N__19905),
            .I(N__19900));
    LocalMux I__3614 (
            .O(N__19900),
            .I(N__19897));
    Span4Mux_h I__3613 (
            .O(N__19897),
            .I(N__19894));
    Odrv4 I__3612 (
            .O(N__19894),
            .I(\c0.n2036 ));
    InMux I__3611 (
            .O(N__19891),
            .I(N__19888));
    LocalMux I__3610 (
            .O(N__19888),
            .I(\c0.n20_adj_1892 ));
    InMux I__3609 (
            .O(N__19885),
            .I(N__19881));
    InMux I__3608 (
            .O(N__19884),
            .I(N__19878));
    LocalMux I__3607 (
            .O(N__19881),
            .I(\c0.n2033 ));
    LocalMux I__3606 (
            .O(N__19878),
            .I(\c0.n2033 ));
    CascadeMux I__3605 (
            .O(N__19873),
            .I(\c0.n10_adj_1963_cascade_ ));
    InMux I__3604 (
            .O(N__19870),
            .I(N__19867));
    LocalMux I__3603 (
            .O(N__19867),
            .I(\c0.n5114 ));
    CascadeMux I__3602 (
            .O(N__19864),
            .I(\c0.n5114_cascade_ ));
    InMux I__3601 (
            .O(N__19861),
            .I(N__19858));
    LocalMux I__3600 (
            .O(N__19858),
            .I(N__19855));
    Odrv4 I__3599 (
            .O(N__19855),
            .I(\c0.n30_adj_1903 ));
    CascadeMux I__3598 (
            .O(N__19852),
            .I(N__19849));
    InMux I__3597 (
            .O(N__19849),
            .I(N__19846));
    LocalMux I__3596 (
            .O(N__19846),
            .I(N__19843));
    Span4Mux_h I__3595 (
            .O(N__19843),
            .I(N__19840));
    Span4Mux_h I__3594 (
            .O(N__19840),
            .I(N__19837));
    Odrv4 I__3593 (
            .O(N__19837),
            .I(\c0.n5743 ));
    InMux I__3592 (
            .O(N__19834),
            .I(N__19831));
    LocalMux I__3591 (
            .O(N__19831),
            .I(N__19827));
    InMux I__3590 (
            .O(N__19830),
            .I(N__19821));
    Span4Mux_s3_v I__3589 (
            .O(N__19827),
            .I(N__19818));
    InMux I__3588 (
            .O(N__19826),
            .I(N__19811));
    InMux I__3587 (
            .O(N__19825),
            .I(N__19811));
    InMux I__3586 (
            .O(N__19824),
            .I(N__19811));
    LocalMux I__3585 (
            .O(N__19821),
            .I(\c0.data_in_field_87 ));
    Odrv4 I__3584 (
            .O(N__19818),
            .I(\c0.data_in_field_87 ));
    LocalMux I__3583 (
            .O(N__19811),
            .I(\c0.data_in_field_87 ));
    CascadeMux I__3582 (
            .O(N__19804),
            .I(N__19801));
    InMux I__3581 (
            .O(N__19801),
            .I(N__19797));
    InMux I__3580 (
            .O(N__19800),
            .I(N__19794));
    LocalMux I__3579 (
            .O(N__19797),
            .I(N__19788));
    LocalMux I__3578 (
            .O(N__19794),
            .I(N__19785));
    InMux I__3577 (
            .O(N__19793),
            .I(N__19782));
    InMux I__3576 (
            .O(N__19792),
            .I(N__19777));
    InMux I__3575 (
            .O(N__19791),
            .I(N__19777));
    Span4Mux_v I__3574 (
            .O(N__19788),
            .I(N__19772));
    Span4Mux_s3_v I__3573 (
            .O(N__19785),
            .I(N__19772));
    LocalMux I__3572 (
            .O(N__19782),
            .I(N__19769));
    LocalMux I__3571 (
            .O(N__19777),
            .I(\c0.data_in_field_57 ));
    Odrv4 I__3570 (
            .O(N__19772),
            .I(\c0.data_in_field_57 ));
    Odrv12 I__3569 (
            .O(N__19769),
            .I(\c0.data_in_field_57 ));
    InMux I__3568 (
            .O(N__19762),
            .I(N__19759));
    LocalMux I__3567 (
            .O(N__19759),
            .I(\c0.n5198 ));
    CascadeMux I__3566 (
            .O(N__19756),
            .I(N__19753));
    InMux I__3565 (
            .O(N__19753),
            .I(N__19750));
    LocalMux I__3564 (
            .O(N__19750),
            .I(N__19747));
    Span4Mux_v I__3563 (
            .O(N__19747),
            .I(N__19743));
    InMux I__3562 (
            .O(N__19746),
            .I(N__19740));
    Span4Mux_h I__3561 (
            .O(N__19743),
            .I(N__19737));
    LocalMux I__3560 (
            .O(N__19740),
            .I(\c0.n1918 ));
    Odrv4 I__3559 (
            .O(N__19737),
            .I(\c0.n1918 ));
    InMux I__3558 (
            .O(N__19732),
            .I(N__19729));
    LocalMux I__3557 (
            .O(N__19729),
            .I(\c0.n18_adj_1910 ));
    CascadeMux I__3556 (
            .O(N__19726),
            .I(\c0.n17_adj_1912_cascade_ ));
    InMux I__3555 (
            .O(N__19723),
            .I(N__19720));
    LocalMux I__3554 (
            .O(N__19720),
            .I(\c0.n12_adj_1911 ));
    InMux I__3553 (
            .O(N__19717),
            .I(N__19714));
    LocalMux I__3552 (
            .O(N__19714),
            .I(\c0.n19_adj_1920 ));
    InMux I__3551 (
            .O(N__19711),
            .I(N__19708));
    LocalMux I__3550 (
            .O(N__19708),
            .I(\c0.n28_adj_1902 ));
    InMux I__3549 (
            .O(N__19705),
            .I(N__19702));
    LocalMux I__3548 (
            .O(N__19702),
            .I(\c0.n32 ));
    CascadeMux I__3547 (
            .O(N__19699),
            .I(\c0.n29_adj_1905_cascade_ ));
    InMux I__3546 (
            .O(N__19696),
            .I(N__19693));
    LocalMux I__3545 (
            .O(N__19693),
            .I(\c0.n31_adj_1904 ));
    InMux I__3544 (
            .O(N__19690),
            .I(N__19687));
    LocalMux I__3543 (
            .O(N__19687),
            .I(N__19684));
    Odrv4 I__3542 (
            .O(N__19684),
            .I(\c0.n5278 ));
    InMux I__3541 (
            .O(N__19681),
            .I(N__19677));
    InMux I__3540 (
            .O(N__19680),
            .I(N__19674));
    LocalMux I__3539 (
            .O(N__19677),
            .I(N__19671));
    LocalMux I__3538 (
            .O(N__19674),
            .I(N__19663));
    Span4Mux_h I__3537 (
            .O(N__19671),
            .I(N__19663));
    InMux I__3536 (
            .O(N__19670),
            .I(N__19660));
    InMux I__3535 (
            .O(N__19669),
            .I(N__19657));
    InMux I__3534 (
            .O(N__19668),
            .I(N__19654));
    Odrv4 I__3533 (
            .O(N__19663),
            .I(\c0.data_in_field_134 ));
    LocalMux I__3532 (
            .O(N__19660),
            .I(\c0.data_in_field_134 ));
    LocalMux I__3531 (
            .O(N__19657),
            .I(\c0.data_in_field_134 ));
    LocalMux I__3530 (
            .O(N__19654),
            .I(\c0.data_in_field_134 ));
    CascadeMux I__3529 (
            .O(N__19645),
            .I(\c0.n12_cascade_ ));
    InMux I__3528 (
            .O(N__19642),
            .I(N__19638));
    InMux I__3527 (
            .O(N__19641),
            .I(N__19635));
    LocalMux I__3526 (
            .O(N__19638),
            .I(\c0.n1880 ));
    LocalMux I__3525 (
            .O(N__19635),
            .I(\c0.n1880 ));
    InMux I__3524 (
            .O(N__19630),
            .I(N__19626));
    InMux I__3523 (
            .O(N__19629),
            .I(N__19623));
    LocalMux I__3522 (
            .O(N__19626),
            .I(N__19620));
    LocalMux I__3521 (
            .O(N__19623),
            .I(N__19615));
    Span4Mux_h I__3520 (
            .O(N__19620),
            .I(N__19615));
    Sp12to4 I__3519 (
            .O(N__19615),
            .I(N__19611));
    InMux I__3518 (
            .O(N__19614),
            .I(N__19608));
    Odrv12 I__3517 (
            .O(N__19611),
            .I(data_in_15_0));
    LocalMux I__3516 (
            .O(N__19608),
            .I(data_in_15_0));
    InMux I__3515 (
            .O(N__19603),
            .I(N__19597));
    InMux I__3514 (
            .O(N__19602),
            .I(N__19597));
    LocalMux I__3513 (
            .O(N__19597),
            .I(N__19594));
    Odrv4 I__3512 (
            .O(N__19594),
            .I(\c0.n5210 ));
    InMux I__3511 (
            .O(N__19591),
            .I(N__19588));
    LocalMux I__3510 (
            .O(N__19588),
            .I(\c0.tx2_transmit_N_1031 ));
    InMux I__3509 (
            .O(N__19585),
            .I(N__19581));
    CascadeMux I__3508 (
            .O(N__19584),
            .I(N__19578));
    LocalMux I__3507 (
            .O(N__19581),
            .I(N__19575));
    InMux I__3506 (
            .O(N__19578),
            .I(N__19572));
    Odrv4 I__3505 (
            .O(N__19575),
            .I(\c0.n1785 ));
    LocalMux I__3504 (
            .O(N__19572),
            .I(\c0.n1785 ));
    InMux I__3503 (
            .O(N__19567),
            .I(N__19564));
    LocalMux I__3502 (
            .O(N__19564),
            .I(\c0.n11 ));
    InMux I__3501 (
            .O(N__19561),
            .I(N__19558));
    LocalMux I__3500 (
            .O(N__19558),
            .I(N__19555));
    Odrv4 I__3499 (
            .O(N__19555),
            .I(\c0.n24_adj_1924 ));
    CascadeMux I__3498 (
            .O(N__19552),
            .I(\c0.n5259_cascade_ ));
    CascadeMux I__3497 (
            .O(N__19549),
            .I(N__19546));
    InMux I__3496 (
            .O(N__19546),
            .I(N__19543));
    LocalMux I__3495 (
            .O(N__19543),
            .I(\c0.n21_adj_1933 ));
    InMux I__3494 (
            .O(N__19540),
            .I(N__19537));
    LocalMux I__3493 (
            .O(N__19537),
            .I(N__19534));
    Odrv4 I__3492 (
            .O(N__19534),
            .I(\c0.n16 ));
    CascadeMux I__3491 (
            .O(N__19531),
            .I(N__19528));
    InMux I__3490 (
            .O(N__19528),
            .I(N__19525));
    LocalMux I__3489 (
            .O(N__19525),
            .I(N__19522));
    Span4Mux_h I__3488 (
            .O(N__19522),
            .I(N__19519));
    Span4Mux_s3_h I__3487 (
            .O(N__19519),
            .I(N__19515));
    InMux I__3486 (
            .O(N__19518),
            .I(N__19512));
    Odrv4 I__3485 (
            .O(N__19515),
            .I(\c0.n1893 ));
    LocalMux I__3484 (
            .O(N__19512),
            .I(\c0.n1893 ));
    InMux I__3483 (
            .O(N__19507),
            .I(N__19504));
    LocalMux I__3482 (
            .O(N__19504),
            .I(N__19500));
    InMux I__3481 (
            .O(N__19503),
            .I(N__19497));
    Span4Mux_h I__3480 (
            .O(N__19500),
            .I(N__19494));
    LocalMux I__3479 (
            .O(N__19497),
            .I(N__19491));
    Odrv4 I__3478 (
            .O(N__19494),
            .I(\c0.n2008 ));
    Odrv4 I__3477 (
            .O(N__19491),
            .I(\c0.n2008 ));
    InMux I__3476 (
            .O(N__19486),
            .I(N__19483));
    LocalMux I__3475 (
            .O(N__19483),
            .I(N__19480));
    Odrv4 I__3474 (
            .O(N__19480),
            .I(\c0.n5225 ));
    CascadeMux I__3473 (
            .O(N__19477),
            .I(\c0.n5198_cascade_ ));
    InMux I__3472 (
            .O(N__19474),
            .I(N__19471));
    LocalMux I__3471 (
            .O(N__19471),
            .I(N__19467));
    InMux I__3470 (
            .O(N__19470),
            .I(N__19464));
    Span4Mux_h I__3469 (
            .O(N__19467),
            .I(N__19461));
    LocalMux I__3468 (
            .O(N__19464),
            .I(N__19458));
    Odrv4 I__3467 (
            .O(N__19461),
            .I(\c0.n6103 ));
    Odrv4 I__3466 (
            .O(N__19458),
            .I(\c0.n6103 ));
    InMux I__3465 (
            .O(N__19453),
            .I(N__19450));
    LocalMux I__3464 (
            .O(N__19450),
            .I(\c0.n28 ));
    CascadeMux I__3463 (
            .O(N__19447),
            .I(N__19444));
    InMux I__3462 (
            .O(N__19444),
            .I(N__19441));
    LocalMux I__3461 (
            .O(N__19441),
            .I(N__19437));
    InMux I__3460 (
            .O(N__19440),
            .I(N__19434));
    Span4Mux_v I__3459 (
            .O(N__19437),
            .I(N__19430));
    LocalMux I__3458 (
            .O(N__19434),
            .I(N__19427));
    InMux I__3457 (
            .O(N__19433),
            .I(N__19424));
    Odrv4 I__3456 (
            .O(N__19430),
            .I(data_in_14_5));
    Odrv12 I__3455 (
            .O(N__19427),
            .I(data_in_14_5));
    LocalMux I__3454 (
            .O(N__19424),
            .I(data_in_14_5));
    CascadeMux I__3453 (
            .O(N__19417),
            .I(N__19414));
    InMux I__3452 (
            .O(N__19414),
            .I(N__19411));
    LocalMux I__3451 (
            .O(N__19411),
            .I(N__19408));
    Span4Mux_h I__3450 (
            .O(N__19408),
            .I(N__19405));
    Odrv4 I__3449 (
            .O(N__19405),
            .I(\c0.n5809 ));
    CascadeMux I__3448 (
            .O(N__19402),
            .I(N__19399));
    InMux I__3447 (
            .O(N__19399),
            .I(N__19396));
    LocalMux I__3446 (
            .O(N__19396),
            .I(N__19393));
    Odrv4 I__3445 (
            .O(N__19393),
            .I(\c0.n5241 ));
    CascadeMux I__3444 (
            .O(N__19390),
            .I(\c0.tx2_transmit_N_1031_cascade_ ));
    InMux I__3443 (
            .O(N__19387),
            .I(N__19384));
    LocalMux I__3442 (
            .O(N__19384),
            .I(N__19381));
    Odrv4 I__3441 (
            .O(N__19381),
            .I(\c0.n38_adj_1934 ));
    InMux I__3440 (
            .O(N__19378),
            .I(N__19375));
    LocalMux I__3439 (
            .O(N__19375),
            .I(\c0.n14_adj_1900 ));
    InMux I__3438 (
            .O(N__19372),
            .I(N__19363));
    InMux I__3437 (
            .O(N__19371),
            .I(N__19363));
    InMux I__3436 (
            .O(N__19370),
            .I(N__19360));
    InMux I__3435 (
            .O(N__19369),
            .I(N__19357));
    InMux I__3434 (
            .O(N__19368),
            .I(N__19354));
    LocalMux I__3433 (
            .O(N__19363),
            .I(N__19351));
    LocalMux I__3432 (
            .O(N__19360),
            .I(N__19346));
    LocalMux I__3431 (
            .O(N__19357),
            .I(N__19346));
    LocalMux I__3430 (
            .O(N__19354),
            .I(N__19343));
    Span4Mux_v I__3429 (
            .O(N__19351),
            .I(N__19337));
    Span4Mux_v I__3428 (
            .O(N__19346),
            .I(N__19332));
    Span4Mux_v I__3427 (
            .O(N__19343),
            .I(N__19332));
    InMux I__3426 (
            .O(N__19342),
            .I(N__19329));
    InMux I__3425 (
            .O(N__19341),
            .I(N__19326));
    InMux I__3424 (
            .O(N__19340),
            .I(N__19323));
    Odrv4 I__3423 (
            .O(N__19337),
            .I(n1442));
    Odrv4 I__3422 (
            .O(N__19332),
            .I(n1442));
    LocalMux I__3421 (
            .O(N__19329),
            .I(n1442));
    LocalMux I__3420 (
            .O(N__19326),
            .I(n1442));
    LocalMux I__3419 (
            .O(N__19323),
            .I(n1442));
    InMux I__3418 (
            .O(N__19312),
            .I(N__19308));
    InMux I__3417 (
            .O(N__19311),
            .I(N__19305));
    LocalMux I__3416 (
            .O(N__19308),
            .I(r_Tx_Data_6));
    LocalMux I__3415 (
            .O(N__19305),
            .I(r_Tx_Data_6));
    InMux I__3414 (
            .O(N__19300),
            .I(N__19293));
    InMux I__3413 (
            .O(N__19299),
            .I(N__19287));
    InMux I__3412 (
            .O(N__19298),
            .I(N__19287));
    InMux I__3411 (
            .O(N__19297),
            .I(N__19284));
    InMux I__3410 (
            .O(N__19296),
            .I(N__19279));
    LocalMux I__3409 (
            .O(N__19293),
            .I(N__19276));
    InMux I__3408 (
            .O(N__19292),
            .I(N__19273));
    LocalMux I__3407 (
            .O(N__19287),
            .I(N__19268));
    LocalMux I__3406 (
            .O(N__19284),
            .I(N__19268));
    InMux I__3405 (
            .O(N__19283),
            .I(N__19265));
    InMux I__3404 (
            .O(N__19282),
            .I(N__19262));
    LocalMux I__3403 (
            .O(N__19279),
            .I(N__19257));
    Span4Mux_v I__3402 (
            .O(N__19276),
            .I(N__19257));
    LocalMux I__3401 (
            .O(N__19273),
            .I(N__19252));
    Span4Mux_h I__3400 (
            .O(N__19268),
            .I(N__19252));
    LocalMux I__3399 (
            .O(N__19265),
            .I(N__19249));
    LocalMux I__3398 (
            .O(N__19262),
            .I(data_out_10_0));
    Odrv4 I__3397 (
            .O(N__19257),
            .I(data_out_10_0));
    Odrv4 I__3396 (
            .O(N__19252),
            .I(data_out_10_0));
    Odrv12 I__3395 (
            .O(N__19249),
            .I(data_out_10_0));
    InMux I__3394 (
            .O(N__19240),
            .I(N__19237));
    LocalMux I__3393 (
            .O(N__19237),
            .I(N__19234));
    Span4Mux_v I__3392 (
            .O(N__19234),
            .I(N__19231));
    Span4Mux_s3_h I__3391 (
            .O(N__19231),
            .I(N__19228));
    Odrv4 I__3390 (
            .O(N__19228),
            .I(n1748));
    InMux I__3389 (
            .O(N__19225),
            .I(N__19217));
    InMux I__3388 (
            .O(N__19224),
            .I(N__19214));
    CascadeMux I__3387 (
            .O(N__19223),
            .I(N__19210));
    InMux I__3386 (
            .O(N__19222),
            .I(N__19202));
    InMux I__3385 (
            .O(N__19221),
            .I(N__19202));
    InMux I__3384 (
            .O(N__19220),
            .I(N__19199));
    LocalMux I__3383 (
            .O(N__19217),
            .I(N__19196));
    LocalMux I__3382 (
            .O(N__19214),
            .I(N__19193));
    InMux I__3381 (
            .O(N__19213),
            .I(N__19188));
    InMux I__3380 (
            .O(N__19210),
            .I(N__19188));
    InMux I__3379 (
            .O(N__19209),
            .I(N__19185));
    InMux I__3378 (
            .O(N__19208),
            .I(N__19182));
    InMux I__3377 (
            .O(N__19207),
            .I(N__19171));
    LocalMux I__3376 (
            .O(N__19202),
            .I(N__19168));
    LocalMux I__3375 (
            .O(N__19199),
            .I(N__19160));
    Span4Mux_h I__3374 (
            .O(N__19196),
            .I(N__19160));
    Span4Mux_h I__3373 (
            .O(N__19193),
            .I(N__19160));
    LocalMux I__3372 (
            .O(N__19188),
            .I(N__19153));
    LocalMux I__3371 (
            .O(N__19185),
            .I(N__19153));
    LocalMux I__3370 (
            .O(N__19182),
            .I(N__19153));
    InMux I__3369 (
            .O(N__19181),
            .I(N__19142));
    InMux I__3368 (
            .O(N__19180),
            .I(N__19142));
    InMux I__3367 (
            .O(N__19179),
            .I(N__19142));
    InMux I__3366 (
            .O(N__19178),
            .I(N__19142));
    InMux I__3365 (
            .O(N__19177),
            .I(N__19142));
    InMux I__3364 (
            .O(N__19176),
            .I(N__19135));
    InMux I__3363 (
            .O(N__19175),
            .I(N__19135));
    InMux I__3362 (
            .O(N__19174),
            .I(N__19135));
    LocalMux I__3361 (
            .O(N__19171),
            .I(N__19132));
    Span4Mux_h I__3360 (
            .O(N__19168),
            .I(N__19129));
    InMux I__3359 (
            .O(N__19167),
            .I(N__19126));
    Span4Mux_v I__3358 (
            .O(N__19160),
            .I(N__19123));
    Span4Mux_h I__3357 (
            .O(N__19153),
            .I(N__19118));
    LocalMux I__3356 (
            .O(N__19142),
            .I(N__19118));
    LocalMux I__3355 (
            .O(N__19135),
            .I(n21_adj_1999));
    Odrv4 I__3354 (
            .O(N__19132),
            .I(n21_adj_1999));
    Odrv4 I__3353 (
            .O(N__19129),
            .I(n21_adj_1999));
    LocalMux I__3352 (
            .O(N__19126),
            .I(n21_adj_1999));
    Odrv4 I__3351 (
            .O(N__19123),
            .I(n21_adj_1999));
    Odrv4 I__3350 (
            .O(N__19118),
            .I(n21_adj_1999));
    CascadeMux I__3349 (
            .O(N__19105),
            .I(N__19102));
    InMux I__3348 (
            .O(N__19102),
            .I(N__19099));
    LocalMux I__3347 (
            .O(N__19099),
            .I(N__19095));
    InMux I__3346 (
            .O(N__19098),
            .I(N__19092));
    Odrv12 I__3345 (
            .O(N__19095),
            .I(data_10));
    LocalMux I__3344 (
            .O(N__19092),
            .I(data_10));
    InMux I__3343 (
            .O(N__19087),
            .I(N__19084));
    LocalMux I__3342 (
            .O(N__19084),
            .I(N__19075));
    InMux I__3341 (
            .O(N__19083),
            .I(N__19072));
    InMux I__3340 (
            .O(N__19082),
            .I(N__19065));
    InMux I__3339 (
            .O(N__19081),
            .I(N__19065));
    InMux I__3338 (
            .O(N__19080),
            .I(N__19065));
    InMux I__3337 (
            .O(N__19079),
            .I(N__19062));
    InMux I__3336 (
            .O(N__19078),
            .I(N__19059));
    Span4Mux_h I__3335 (
            .O(N__19075),
            .I(N__19051));
    LocalMux I__3334 (
            .O(N__19072),
            .I(N__19051));
    LocalMux I__3333 (
            .O(N__19065),
            .I(N__19046));
    LocalMux I__3332 (
            .O(N__19062),
            .I(N__19046));
    LocalMux I__3331 (
            .O(N__19059),
            .I(N__19043));
    InMux I__3330 (
            .O(N__19058),
            .I(N__19040));
    InMux I__3329 (
            .O(N__19057),
            .I(N__19035));
    InMux I__3328 (
            .O(N__19056),
            .I(N__19035));
    Span4Mux_v I__3327 (
            .O(N__19051),
            .I(N__19024));
    Span4Mux_h I__3326 (
            .O(N__19046),
            .I(N__19021));
    Span4Mux_h I__3325 (
            .O(N__19043),
            .I(N__19016));
    LocalMux I__3324 (
            .O(N__19040),
            .I(N__19016));
    LocalMux I__3323 (
            .O(N__19035),
            .I(N__19013));
    InMux I__3322 (
            .O(N__19034),
            .I(N__19008));
    InMux I__3321 (
            .O(N__19033),
            .I(N__19008));
    InMux I__3320 (
            .O(N__19032),
            .I(N__18997));
    InMux I__3319 (
            .O(N__19031),
            .I(N__18997));
    InMux I__3318 (
            .O(N__19030),
            .I(N__18997));
    InMux I__3317 (
            .O(N__19029),
            .I(N__18997));
    InMux I__3316 (
            .O(N__19028),
            .I(N__18997));
    InMux I__3315 (
            .O(N__19027),
            .I(N__18994));
    Odrv4 I__3314 (
            .O(N__19024),
            .I(n4315));
    Odrv4 I__3313 (
            .O(N__19021),
            .I(n4315));
    Odrv4 I__3312 (
            .O(N__19016),
            .I(n4315));
    Odrv4 I__3311 (
            .O(N__19013),
            .I(n4315));
    LocalMux I__3310 (
            .O(N__19008),
            .I(n4315));
    LocalMux I__3309 (
            .O(N__18997),
            .I(n4315));
    LocalMux I__3308 (
            .O(N__18994),
            .I(n4315));
    InMux I__3307 (
            .O(N__18979),
            .I(N__18973));
    InMux I__3306 (
            .O(N__18978),
            .I(N__18968));
    InMux I__3305 (
            .O(N__18977),
            .I(N__18968));
    InMux I__3304 (
            .O(N__18976),
            .I(N__18964));
    LocalMux I__3303 (
            .O(N__18973),
            .I(N__18959));
    LocalMux I__3302 (
            .O(N__18968),
            .I(N__18959));
    InMux I__3301 (
            .O(N__18967),
            .I(N__18956));
    LocalMux I__3300 (
            .O(N__18964),
            .I(N__18951));
    Span4Mux_v I__3299 (
            .O(N__18959),
            .I(N__18946));
    LocalMux I__3298 (
            .O(N__18956),
            .I(N__18946));
    InMux I__3297 (
            .O(N__18955),
            .I(N__18943));
    InMux I__3296 (
            .O(N__18954),
            .I(N__18940));
    Span4Mux_v I__3295 (
            .O(N__18951),
            .I(N__18935));
    Span4Mux_h I__3294 (
            .O(N__18946),
            .I(N__18935));
    LocalMux I__3293 (
            .O(N__18943),
            .I(data_out_10_2));
    LocalMux I__3292 (
            .O(N__18940),
            .I(data_out_10_2));
    Odrv4 I__3291 (
            .O(N__18935),
            .I(data_out_10_2));
    InMux I__3290 (
            .O(N__18928),
            .I(N__18925));
    LocalMux I__3289 (
            .O(N__18925),
            .I(N__18922));
    Span4Mux_h I__3288 (
            .O(N__18922),
            .I(N__18919));
    Odrv4 I__3287 (
            .O(N__18919),
            .I(\c0.n5411 ));
    InMux I__3286 (
            .O(N__18916),
            .I(N__18913));
    LocalMux I__3285 (
            .O(N__18913),
            .I(N__18910));
    Span4Mux_h I__3284 (
            .O(N__18910),
            .I(N__18907));
    Odrv4 I__3283 (
            .O(N__18907),
            .I(\c0.n5830 ));
    CascadeMux I__3282 (
            .O(N__18904),
            .I(N__18901));
    InMux I__3281 (
            .O(N__18901),
            .I(N__18898));
    LocalMux I__3280 (
            .O(N__18898),
            .I(N__18895));
    Span4Mux_h I__3279 (
            .O(N__18895),
            .I(N__18892));
    Odrv4 I__3278 (
            .O(N__18892),
            .I(\c0.n5941 ));
    CascadeMux I__3277 (
            .O(N__18889),
            .I(N__18885));
    InMux I__3276 (
            .O(N__18888),
            .I(N__18882));
    InMux I__3275 (
            .O(N__18885),
            .I(N__18879));
    LocalMux I__3274 (
            .O(N__18882),
            .I(\c0.data_in_frame_19_2 ));
    LocalMux I__3273 (
            .O(N__18879),
            .I(\c0.data_in_frame_19_2 ));
    CascadeMux I__3272 (
            .O(N__18874),
            .I(N__18871));
    InMux I__3271 (
            .O(N__18871),
            .I(N__18865));
    InMux I__3270 (
            .O(N__18870),
            .I(N__18865));
    LocalMux I__3269 (
            .O(N__18865),
            .I(\c0.data_in_frame_18_5 ));
    CascadeMux I__3268 (
            .O(N__18862),
            .I(N__18858));
    InMux I__3267 (
            .O(N__18861),
            .I(N__18853));
    InMux I__3266 (
            .O(N__18858),
            .I(N__18853));
    LocalMux I__3265 (
            .O(N__18853),
            .I(\c0.data_in_frame_19_5 ));
    CascadeMux I__3264 (
            .O(N__18850),
            .I(N__18847));
    InMux I__3263 (
            .O(N__18847),
            .I(N__18844));
    LocalMux I__3262 (
            .O(N__18844),
            .I(N__18840));
    InMux I__3261 (
            .O(N__18843),
            .I(N__18837));
    Odrv4 I__3260 (
            .O(N__18840),
            .I(data_4));
    LocalMux I__3259 (
            .O(N__18837),
            .I(data_4));
    CascadeMux I__3258 (
            .O(N__18832),
            .I(N__18829));
    InMux I__3257 (
            .O(N__18829),
            .I(N__18825));
    InMux I__3256 (
            .O(N__18828),
            .I(N__18822));
    LocalMux I__3255 (
            .O(N__18825),
            .I(data_14));
    LocalMux I__3254 (
            .O(N__18822),
            .I(data_14));
    CascadeMux I__3253 (
            .O(N__18817),
            .I(N__18814));
    InMux I__3252 (
            .O(N__18814),
            .I(N__18810));
    CascadeMux I__3251 (
            .O(N__18813),
            .I(N__18807));
    LocalMux I__3250 (
            .O(N__18810),
            .I(N__18802));
    InMux I__3249 (
            .O(N__18807),
            .I(N__18799));
    InMux I__3248 (
            .O(N__18806),
            .I(N__18796));
    InMux I__3247 (
            .O(N__18805),
            .I(N__18793));
    Span4Mux_h I__3246 (
            .O(N__18802),
            .I(N__18785));
    LocalMux I__3245 (
            .O(N__18799),
            .I(N__18785));
    LocalMux I__3244 (
            .O(N__18796),
            .I(N__18785));
    LocalMux I__3243 (
            .O(N__18793),
            .I(N__18782));
    InMux I__3242 (
            .O(N__18792),
            .I(N__18776));
    Span4Mux_v I__3241 (
            .O(N__18785),
            .I(N__18771));
    Span4Mux_h I__3240 (
            .O(N__18782),
            .I(N__18771));
    InMux I__3239 (
            .O(N__18781),
            .I(N__18768));
    InMux I__3238 (
            .O(N__18780),
            .I(N__18763));
    InMux I__3237 (
            .O(N__18779),
            .I(N__18763));
    LocalMux I__3236 (
            .O(N__18776),
            .I(data_out_11_4));
    Odrv4 I__3235 (
            .O(N__18771),
            .I(data_out_11_4));
    LocalMux I__3234 (
            .O(N__18768),
            .I(data_out_11_4));
    LocalMux I__3233 (
            .O(N__18763),
            .I(data_out_11_4));
    InMux I__3232 (
            .O(N__18754),
            .I(N__18751));
    LocalMux I__3231 (
            .O(N__18751),
            .I(N__18745));
    InMux I__3230 (
            .O(N__18750),
            .I(N__18742));
    CascadeMux I__3229 (
            .O(N__18749),
            .I(N__18739));
    InMux I__3228 (
            .O(N__18748),
            .I(N__18736));
    Span4Mux_s3_h I__3227 (
            .O(N__18745),
            .I(N__18730));
    LocalMux I__3226 (
            .O(N__18742),
            .I(N__18730));
    InMux I__3225 (
            .O(N__18739),
            .I(N__18727));
    LocalMux I__3224 (
            .O(N__18736),
            .I(N__18724));
    InMux I__3223 (
            .O(N__18735),
            .I(N__18721));
    Span4Mux_h I__3222 (
            .O(N__18730),
            .I(N__18718));
    LocalMux I__3221 (
            .O(N__18727),
            .I(data_out_10_4));
    Odrv4 I__3220 (
            .O(N__18724),
            .I(data_out_10_4));
    LocalMux I__3219 (
            .O(N__18721),
            .I(data_out_10_4));
    Odrv4 I__3218 (
            .O(N__18718),
            .I(data_out_10_4));
    CascadeMux I__3217 (
            .O(N__18709),
            .I(\c0.n9_adj_1887_cascade_ ));
    InMux I__3216 (
            .O(N__18706),
            .I(N__18703));
    LocalMux I__3215 (
            .O(N__18703),
            .I(N__18700));
    Odrv12 I__3214 (
            .O(N__18700),
            .I(\c0.n15_adj_1889 ));
    InMux I__3213 (
            .O(N__18697),
            .I(N__18693));
    InMux I__3212 (
            .O(N__18696),
            .I(N__18690));
    LocalMux I__3211 (
            .O(N__18693),
            .I(data_8));
    LocalMux I__3210 (
            .O(N__18690),
            .I(data_8));
    InMux I__3209 (
            .O(N__18685),
            .I(N__18682));
    LocalMux I__3208 (
            .O(N__18682),
            .I(N__18679));
    Span4Mux_v I__3207 (
            .O(N__18679),
            .I(N__18676));
    Odrv4 I__3206 (
            .O(N__18676),
            .I(\c0.n17_adj_1961 ));
    CascadeMux I__3205 (
            .O(N__18673),
            .I(\c0.n1236_cascade_ ));
    InMux I__3204 (
            .O(N__18670),
            .I(N__18667));
    LocalMux I__3203 (
            .O(N__18667),
            .I(\c0.n2247 ));
    InMux I__3202 (
            .O(N__18664),
            .I(N__18661));
    LocalMux I__3201 (
            .O(N__18661),
            .I(N__18658));
    Span4Mux_v I__3200 (
            .O(N__18658),
            .I(N__18654));
    InMux I__3199 (
            .O(N__18657),
            .I(N__18651));
    Odrv4 I__3198 (
            .O(N__18654),
            .I(\c0.n1227 ));
    LocalMux I__3197 (
            .O(N__18651),
            .I(\c0.n1227 ));
    CascadeMux I__3196 (
            .O(N__18646),
            .I(\c0.n5511_cascade_ ));
    CascadeMux I__3195 (
            .O(N__18643),
            .I(tx_data_7_N_keep_cascade_));
    InMux I__3194 (
            .O(N__18640),
            .I(N__18636));
    InMux I__3193 (
            .O(N__18639),
            .I(N__18633));
    LocalMux I__3192 (
            .O(N__18636),
            .I(r_Tx_Data_7));
    LocalMux I__3191 (
            .O(N__18633),
            .I(r_Tx_Data_7));
    CascadeMux I__3190 (
            .O(N__18628),
            .I(N__18625));
    InMux I__3189 (
            .O(N__18625),
            .I(N__18622));
    LocalMux I__3188 (
            .O(N__18622),
            .I(N__18619));
    Span4Mux_h I__3187 (
            .O(N__18619),
            .I(N__18615));
    InMux I__3186 (
            .O(N__18618),
            .I(N__18612));
    Odrv4 I__3185 (
            .O(N__18615),
            .I(data_7));
    LocalMux I__3184 (
            .O(N__18612),
            .I(data_7));
    InMux I__3183 (
            .O(N__18607),
            .I(\c0.n4391 ));
    InMux I__3182 (
            .O(N__18604),
            .I(bfn_6_18_0_));
    CascadeMux I__3181 (
            .O(N__18601),
            .I(N__18598));
    InMux I__3180 (
            .O(N__18598),
            .I(N__18595));
    LocalMux I__3179 (
            .O(N__18595),
            .I(N__18592));
    Span4Mux_v I__3178 (
            .O(N__18592),
            .I(N__18588));
    InMux I__3177 (
            .O(N__18591),
            .I(N__18585));
    Odrv4 I__3176 (
            .O(N__18588),
            .I(data_9));
    LocalMux I__3175 (
            .O(N__18585),
            .I(data_9));
    InMux I__3174 (
            .O(N__18580),
            .I(\c0.n4393 ));
    InMux I__3173 (
            .O(N__18577),
            .I(\c0.n4394 ));
    CascadeMux I__3172 (
            .O(N__18574),
            .I(N__18571));
    InMux I__3171 (
            .O(N__18571),
            .I(N__18568));
    LocalMux I__3170 (
            .O(N__18568),
            .I(N__18564));
    InMux I__3169 (
            .O(N__18567),
            .I(N__18561));
    Odrv12 I__3168 (
            .O(N__18564),
            .I(data_11));
    LocalMux I__3167 (
            .O(N__18561),
            .I(data_11));
    InMux I__3166 (
            .O(N__18556),
            .I(\c0.n4395 ));
    InMux I__3165 (
            .O(N__18553),
            .I(N__18550));
    LocalMux I__3164 (
            .O(N__18550),
            .I(N__18546));
    InMux I__3163 (
            .O(N__18549),
            .I(N__18543));
    Odrv4 I__3162 (
            .O(N__18546),
            .I(data_12));
    LocalMux I__3161 (
            .O(N__18543),
            .I(data_12));
    InMux I__3160 (
            .O(N__18538),
            .I(\c0.n4396 ));
    CascadeMux I__3159 (
            .O(N__18535),
            .I(N__18532));
    InMux I__3158 (
            .O(N__18532),
            .I(N__18529));
    LocalMux I__3157 (
            .O(N__18529),
            .I(N__18525));
    InMux I__3156 (
            .O(N__18528),
            .I(N__18522));
    Odrv4 I__3155 (
            .O(N__18525),
            .I(data_13));
    LocalMux I__3154 (
            .O(N__18522),
            .I(data_13));
    InMux I__3153 (
            .O(N__18517),
            .I(\c0.n4397 ));
    InMux I__3152 (
            .O(N__18514),
            .I(\c0.n4398 ));
    InMux I__3151 (
            .O(N__18511),
            .I(\c0.n4399 ));
    CascadeMux I__3150 (
            .O(N__18508),
            .I(N__18505));
    InMux I__3149 (
            .O(N__18505),
            .I(N__18501));
    InMux I__3148 (
            .O(N__18504),
            .I(N__18498));
    LocalMux I__3147 (
            .O(N__18501),
            .I(N__18495));
    LocalMux I__3146 (
            .O(N__18498),
            .I(data_15));
    Odrv4 I__3145 (
            .O(N__18495),
            .I(data_15));
    CascadeMux I__3144 (
            .O(N__18490),
            .I(N__18487));
    InMux I__3143 (
            .O(N__18487),
            .I(N__18483));
    InMux I__3142 (
            .O(N__18486),
            .I(N__18480));
    LocalMux I__3141 (
            .O(N__18483),
            .I(data_0));
    LocalMux I__3140 (
            .O(N__18480),
            .I(data_0));
    InMux I__3139 (
            .O(N__18475),
            .I(bfn_6_17_0_));
    CascadeMux I__3138 (
            .O(N__18472),
            .I(N__18469));
    InMux I__3137 (
            .O(N__18469),
            .I(N__18466));
    LocalMux I__3136 (
            .O(N__18466),
            .I(N__18463));
    Span4Mux_h I__3135 (
            .O(N__18463),
            .I(N__18459));
    InMux I__3134 (
            .O(N__18462),
            .I(N__18456));
    Odrv4 I__3133 (
            .O(N__18459),
            .I(data_1));
    LocalMux I__3132 (
            .O(N__18456),
            .I(data_1));
    InMux I__3131 (
            .O(N__18451),
            .I(\c0.n4385 ));
    CascadeMux I__3130 (
            .O(N__18448),
            .I(N__18445));
    InMux I__3129 (
            .O(N__18445),
            .I(N__18442));
    LocalMux I__3128 (
            .O(N__18442),
            .I(N__18438));
    InMux I__3127 (
            .O(N__18441),
            .I(N__18435));
    Odrv4 I__3126 (
            .O(N__18438),
            .I(data_2));
    LocalMux I__3125 (
            .O(N__18435),
            .I(data_2));
    InMux I__3124 (
            .O(N__18430),
            .I(\c0.n4386 ));
    InMux I__3123 (
            .O(N__18427),
            .I(N__18424));
    LocalMux I__3122 (
            .O(N__18424),
            .I(N__18420));
    InMux I__3121 (
            .O(N__18423),
            .I(N__18417));
    Odrv12 I__3120 (
            .O(N__18420),
            .I(data_3));
    LocalMux I__3119 (
            .O(N__18417),
            .I(data_3));
    InMux I__3118 (
            .O(N__18412),
            .I(\c0.n4387 ));
    InMux I__3117 (
            .O(N__18409),
            .I(\c0.n4388 ));
    CascadeMux I__3116 (
            .O(N__18406),
            .I(N__18403));
    InMux I__3115 (
            .O(N__18403),
            .I(N__18400));
    LocalMux I__3114 (
            .O(N__18400),
            .I(N__18397));
    Span4Mux_s3_h I__3113 (
            .O(N__18397),
            .I(N__18393));
    InMux I__3112 (
            .O(N__18396),
            .I(N__18390));
    Odrv4 I__3111 (
            .O(N__18393),
            .I(data_5));
    LocalMux I__3110 (
            .O(N__18390),
            .I(data_5));
    InMux I__3109 (
            .O(N__18385),
            .I(\c0.n4389 ));
    InMux I__3108 (
            .O(N__18382),
            .I(N__18379));
    LocalMux I__3107 (
            .O(N__18379),
            .I(N__18375));
    InMux I__3106 (
            .O(N__18378),
            .I(N__18372));
    Odrv4 I__3105 (
            .O(N__18375),
            .I(data_6));
    LocalMux I__3104 (
            .O(N__18372),
            .I(data_6));
    InMux I__3103 (
            .O(N__18367),
            .I(\c0.n4390 ));
    CascadeMux I__3102 (
            .O(N__18364),
            .I(N__18358));
    InMux I__3101 (
            .O(N__18363),
            .I(N__18349));
    InMux I__3100 (
            .O(N__18362),
            .I(N__18349));
    InMux I__3099 (
            .O(N__18361),
            .I(N__18344));
    InMux I__3098 (
            .O(N__18358),
            .I(N__18344));
    InMux I__3097 (
            .O(N__18357),
            .I(N__18341));
    CascadeMux I__3096 (
            .O(N__18356),
            .I(N__18338));
    CascadeMux I__3095 (
            .O(N__18355),
            .I(N__18334));
    CascadeMux I__3094 (
            .O(N__18354),
            .I(N__18331));
    LocalMux I__3093 (
            .O(N__18349),
            .I(N__18325));
    LocalMux I__3092 (
            .O(N__18344),
            .I(N__18322));
    LocalMux I__3091 (
            .O(N__18341),
            .I(N__18319));
    InMux I__3090 (
            .O(N__18338),
            .I(N__18314));
    InMux I__3089 (
            .O(N__18337),
            .I(N__18314));
    InMux I__3088 (
            .O(N__18334),
            .I(N__18309));
    InMux I__3087 (
            .O(N__18331),
            .I(N__18309));
    InMux I__3086 (
            .O(N__18330),
            .I(N__18306));
    InMux I__3085 (
            .O(N__18329),
            .I(N__18301));
    InMux I__3084 (
            .O(N__18328),
            .I(N__18301));
    Span4Mux_s1_h I__3083 (
            .O(N__18325),
            .I(N__18292));
    Span4Mux_h I__3082 (
            .O(N__18322),
            .I(N__18292));
    Span4Mux_h I__3081 (
            .O(N__18319),
            .I(N__18292));
    LocalMux I__3080 (
            .O(N__18314),
            .I(N__18292));
    LocalMux I__3079 (
            .O(N__18309),
            .I(r_SM_Main_2_adj_2005));
    LocalMux I__3078 (
            .O(N__18306),
            .I(r_SM_Main_2_adj_2005));
    LocalMux I__3077 (
            .O(N__18301),
            .I(r_SM_Main_2_adj_2005));
    Odrv4 I__3076 (
            .O(N__18292),
            .I(r_SM_Main_2_adj_2005));
    InMux I__3075 (
            .O(N__18283),
            .I(N__18273));
    CascadeMux I__3074 (
            .O(N__18282),
            .I(N__18270));
    InMux I__3073 (
            .O(N__18281),
            .I(N__18261));
    InMux I__3072 (
            .O(N__18280),
            .I(N__18261));
    InMux I__3071 (
            .O(N__18279),
            .I(N__18258));
    InMux I__3070 (
            .O(N__18278),
            .I(N__18255));
    InMux I__3069 (
            .O(N__18277),
            .I(N__18252));
    InMux I__3068 (
            .O(N__18276),
            .I(N__18249));
    LocalMux I__3067 (
            .O(N__18273),
            .I(N__18243));
    InMux I__3066 (
            .O(N__18270),
            .I(N__18238));
    InMux I__3065 (
            .O(N__18269),
            .I(N__18238));
    InMux I__3064 (
            .O(N__18268),
            .I(N__18233));
    InMux I__3063 (
            .O(N__18267),
            .I(N__18233));
    InMux I__3062 (
            .O(N__18266),
            .I(N__18230));
    LocalMux I__3061 (
            .O(N__18261),
            .I(N__18227));
    LocalMux I__3060 (
            .O(N__18258),
            .I(N__18220));
    LocalMux I__3059 (
            .O(N__18255),
            .I(N__18220));
    LocalMux I__3058 (
            .O(N__18252),
            .I(N__18220));
    LocalMux I__3057 (
            .O(N__18249),
            .I(N__18217));
    InMux I__3056 (
            .O(N__18248),
            .I(N__18210));
    InMux I__3055 (
            .O(N__18247),
            .I(N__18210));
    InMux I__3054 (
            .O(N__18246),
            .I(N__18210));
    Span4Mux_v I__3053 (
            .O(N__18243),
            .I(N__18205));
    LocalMux I__3052 (
            .O(N__18238),
            .I(N__18205));
    LocalMux I__3051 (
            .O(N__18233),
            .I(\c0.rx.r_SM_Main_1 ));
    LocalMux I__3050 (
            .O(N__18230),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv4 I__3049 (
            .O(N__18227),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv12 I__3048 (
            .O(N__18220),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv4 I__3047 (
            .O(N__18217),
            .I(\c0.rx.r_SM_Main_1 ));
    LocalMux I__3046 (
            .O(N__18210),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv4 I__3045 (
            .O(N__18205),
            .I(\c0.rx.r_SM_Main_1 ));
    InMux I__3044 (
            .O(N__18190),
            .I(N__18187));
    LocalMux I__3043 (
            .O(N__18187),
            .I(\c0.rx.n5058 ));
    CascadeMux I__3042 (
            .O(N__18184),
            .I(N__18181));
    InMux I__3041 (
            .O(N__18181),
            .I(N__18171));
    InMux I__3040 (
            .O(N__18180),
            .I(N__18171));
    InMux I__3039 (
            .O(N__18179),
            .I(N__18168));
    InMux I__3038 (
            .O(N__18178),
            .I(N__18165));
    CascadeMux I__3037 (
            .O(N__18177),
            .I(N__18162));
    InMux I__3036 (
            .O(N__18176),
            .I(N__18159));
    LocalMux I__3035 (
            .O(N__18171),
            .I(N__18152));
    LocalMux I__3034 (
            .O(N__18168),
            .I(N__18152));
    LocalMux I__3033 (
            .O(N__18165),
            .I(N__18152));
    InMux I__3032 (
            .O(N__18162),
            .I(N__18149));
    LocalMux I__3031 (
            .O(N__18159),
            .I(N__18144));
    Span4Mux_h I__3030 (
            .O(N__18152),
            .I(N__18144));
    LocalMux I__3029 (
            .O(N__18149),
            .I(\c0.rx.r_Bit_Index_0 ));
    Odrv4 I__3028 (
            .O(N__18144),
            .I(\c0.rx.r_Bit_Index_0 ));
    CascadeMux I__3027 (
            .O(N__18139),
            .I(N__18133));
    InMux I__3026 (
            .O(N__18138),
            .I(N__18125));
    InMux I__3025 (
            .O(N__18137),
            .I(N__18125));
    InMux I__3024 (
            .O(N__18136),
            .I(N__18120));
    InMux I__3023 (
            .O(N__18133),
            .I(N__18120));
    InMux I__3022 (
            .O(N__18132),
            .I(N__18117));
    CascadeMux I__3021 (
            .O(N__18131),
            .I(N__18113));
    InMux I__3020 (
            .O(N__18130),
            .I(N__18106));
    LocalMux I__3019 (
            .O(N__18125),
            .I(N__18103));
    LocalMux I__3018 (
            .O(N__18120),
            .I(N__18098));
    LocalMux I__3017 (
            .O(N__18117),
            .I(N__18098));
    InMux I__3016 (
            .O(N__18116),
            .I(N__18091));
    InMux I__3015 (
            .O(N__18113),
            .I(N__18091));
    InMux I__3014 (
            .O(N__18112),
            .I(N__18091));
    InMux I__3013 (
            .O(N__18111),
            .I(N__18086));
    InMux I__3012 (
            .O(N__18110),
            .I(N__18086));
    InMux I__3011 (
            .O(N__18109),
            .I(N__18083));
    LocalMux I__3010 (
            .O(N__18106),
            .I(r_SM_Main_0_adj_2006));
    Odrv4 I__3009 (
            .O(N__18103),
            .I(r_SM_Main_0_adj_2006));
    Odrv12 I__3008 (
            .O(N__18098),
            .I(r_SM_Main_0_adj_2006));
    LocalMux I__3007 (
            .O(N__18091),
            .I(r_SM_Main_0_adj_2006));
    LocalMux I__3006 (
            .O(N__18086),
            .I(r_SM_Main_0_adj_2006));
    LocalMux I__3005 (
            .O(N__18083),
            .I(r_SM_Main_0_adj_2006));
    CascadeMux I__3004 (
            .O(N__18070),
            .I(\c0.rx.n5058_cascade_ ));
    InMux I__3003 (
            .O(N__18067),
            .I(N__18062));
    InMux I__3002 (
            .O(N__18066),
            .I(N__18057));
    InMux I__3001 (
            .O(N__18065),
            .I(N__18057));
    LocalMux I__3000 (
            .O(N__18062),
            .I(N__18050));
    LocalMux I__2999 (
            .O(N__18057),
            .I(N__18050));
    InMux I__2998 (
            .O(N__18056),
            .I(N__18041));
    InMux I__2997 (
            .O(N__18055),
            .I(N__18041));
    Span4Mux_s1_v I__2996 (
            .O(N__18050),
            .I(N__18038));
    InMux I__2995 (
            .O(N__18049),
            .I(N__18035));
    InMux I__2994 (
            .O(N__18048),
            .I(N__18030));
    InMux I__2993 (
            .O(N__18047),
            .I(N__18030));
    InMux I__2992 (
            .O(N__18046),
            .I(N__18027));
    LocalMux I__2991 (
            .O(N__18041),
            .I(\c0.rx.r_SM_Main_2_N_1824_2 ));
    Odrv4 I__2990 (
            .O(N__18038),
            .I(\c0.rx.r_SM_Main_2_N_1824_2 ));
    LocalMux I__2989 (
            .O(N__18035),
            .I(\c0.rx.r_SM_Main_2_N_1824_2 ));
    LocalMux I__2988 (
            .O(N__18030),
            .I(\c0.rx.r_SM_Main_2_N_1824_2 ));
    LocalMux I__2987 (
            .O(N__18027),
            .I(\c0.rx.r_SM_Main_2_N_1824_2 ));
    InMux I__2986 (
            .O(N__18016),
            .I(N__18012));
    InMux I__2985 (
            .O(N__18015),
            .I(N__18009));
    LocalMux I__2984 (
            .O(N__18012),
            .I(N__18004));
    LocalMux I__2983 (
            .O(N__18009),
            .I(N__18004));
    Odrv12 I__2982 (
            .O(N__18004),
            .I(n4));
    CascadeMux I__2981 (
            .O(N__18001),
            .I(n1714_cascade_));
    InMux I__2980 (
            .O(N__17998),
            .I(N__17995));
    LocalMux I__2979 (
            .O(N__17995),
            .I(N__17991));
    InMux I__2978 (
            .O(N__17994),
            .I(N__17988));
    Odrv4 I__2977 (
            .O(N__17991),
            .I(rx_data_1));
    LocalMux I__2976 (
            .O(N__17988),
            .I(rx_data_1));
    InMux I__2975 (
            .O(N__17983),
            .I(N__17978));
    InMux I__2974 (
            .O(N__17982),
            .I(N__17973));
    InMux I__2973 (
            .O(N__17981),
            .I(N__17973));
    LocalMux I__2972 (
            .O(N__17978),
            .I(data_in_0_7));
    LocalMux I__2971 (
            .O(N__17973),
            .I(data_in_0_7));
    InMux I__2970 (
            .O(N__17968),
            .I(N__17965));
    LocalMux I__2969 (
            .O(N__17965),
            .I(N__17961));
    InMux I__2968 (
            .O(N__17964),
            .I(N__17958));
    Odrv4 I__2967 (
            .O(N__17961),
            .I(n4_adj_1986));
    LocalMux I__2966 (
            .O(N__17958),
            .I(n4_adj_1986));
    CascadeMux I__2965 (
            .O(N__17953),
            .I(N__17949));
    InMux I__2964 (
            .O(N__17952),
            .I(N__17945));
    InMux I__2963 (
            .O(N__17949),
            .I(N__17940));
    InMux I__2962 (
            .O(N__17948),
            .I(N__17940));
    LocalMux I__2961 (
            .O(N__17945),
            .I(n1709));
    LocalMux I__2960 (
            .O(N__17940),
            .I(n1709));
    InMux I__2959 (
            .O(N__17935),
            .I(N__17931));
    InMux I__2958 (
            .O(N__17934),
            .I(N__17928));
    LocalMux I__2957 (
            .O(N__17931),
            .I(N__17925));
    LocalMux I__2956 (
            .O(N__17928),
            .I(N__17922));
    Span4Mux_v I__2955 (
            .O(N__17925),
            .I(N__17918));
    Span4Mux_s3_h I__2954 (
            .O(N__17922),
            .I(N__17915));
    InMux I__2953 (
            .O(N__17921),
            .I(N__17912));
    Odrv4 I__2952 (
            .O(N__17918),
            .I(data_in_16_6));
    Odrv4 I__2951 (
            .O(N__17915),
            .I(data_in_16_6));
    LocalMux I__2950 (
            .O(N__17912),
            .I(data_in_16_6));
    CascadeMux I__2949 (
            .O(N__17905),
            .I(N__17902));
    InMux I__2948 (
            .O(N__17902),
            .I(N__17899));
    LocalMux I__2947 (
            .O(N__17899),
            .I(\c0.n5731 ));
    CascadeMux I__2946 (
            .O(N__17896),
            .I(N__17893));
    InMux I__2945 (
            .O(N__17893),
            .I(N__17890));
    LocalMux I__2944 (
            .O(N__17890),
            .I(N__17887));
    Span4Mux_h I__2943 (
            .O(N__17887),
            .I(N__17884));
    Odrv4 I__2942 (
            .O(N__17884),
            .I(\c0.n5264 ));
    CascadeMux I__2941 (
            .O(N__17881),
            .I(\c0.n5264_cascade_ ));
    InMux I__2940 (
            .O(N__17878),
            .I(N__17874));
    CascadeMux I__2939 (
            .O(N__17877),
            .I(N__17871));
    LocalMux I__2938 (
            .O(N__17874),
            .I(N__17868));
    InMux I__2937 (
            .O(N__17871),
            .I(N__17863));
    Span4Mux_h I__2936 (
            .O(N__17868),
            .I(N__17860));
    InMux I__2935 (
            .O(N__17867),
            .I(N__17855));
    InMux I__2934 (
            .O(N__17866),
            .I(N__17855));
    LocalMux I__2933 (
            .O(N__17863),
            .I(N__17852));
    Odrv4 I__2932 (
            .O(N__17860),
            .I(data_in_19_1));
    LocalMux I__2931 (
            .O(N__17855),
            .I(data_in_19_1));
    Odrv12 I__2930 (
            .O(N__17852),
            .I(data_in_19_1));
    InMux I__2929 (
            .O(N__17845),
            .I(N__17841));
    InMux I__2928 (
            .O(N__17844),
            .I(N__17838));
    LocalMux I__2927 (
            .O(N__17841),
            .I(N__17833));
    LocalMux I__2926 (
            .O(N__17838),
            .I(N__17830));
    InMux I__2925 (
            .O(N__17837),
            .I(N__17827));
    InMux I__2924 (
            .O(N__17836),
            .I(N__17824));
    Odrv12 I__2923 (
            .O(N__17833),
            .I(data_in_2_3));
    Odrv4 I__2922 (
            .O(N__17830),
            .I(data_in_2_3));
    LocalMux I__2921 (
            .O(N__17827),
            .I(data_in_2_3));
    LocalMux I__2920 (
            .O(N__17824),
            .I(data_in_2_3));
    InMux I__2919 (
            .O(N__17815),
            .I(N__17812));
    LocalMux I__2918 (
            .O(N__17812),
            .I(\c0.n39 ));
    InMux I__2917 (
            .O(N__17809),
            .I(N__17806));
    LocalMux I__2916 (
            .O(N__17806),
            .I(\c0.n45_adj_1885 ));
    CascadeMux I__2915 (
            .O(N__17803),
            .I(N__17800));
    InMux I__2914 (
            .O(N__17800),
            .I(N__17797));
    LocalMux I__2913 (
            .O(N__17797),
            .I(N__17794));
    Odrv4 I__2912 (
            .O(N__17794),
            .I(\c0.n43 ));
    InMux I__2911 (
            .O(N__17791),
            .I(N__17788));
    LocalMux I__2910 (
            .O(N__17788),
            .I(N__17785));
    Span4Mux_v I__2909 (
            .O(N__17785),
            .I(N__17782));
    Odrv4 I__2908 (
            .O(N__17782),
            .I(\c0.n30 ));
    CascadeMux I__2907 (
            .O(N__17779),
            .I(\c0.n5275_cascade_ ));
    InMux I__2906 (
            .O(N__17776),
            .I(N__17773));
    LocalMux I__2905 (
            .O(N__17773),
            .I(N__17770));
    Span4Mux_h I__2904 (
            .O(N__17770),
            .I(N__17767));
    Odrv4 I__2903 (
            .O(N__17767),
            .I(\c0.n24_adj_1929 ));
    InMux I__2902 (
            .O(N__17764),
            .I(N__17761));
    LocalMux I__2901 (
            .O(N__17761),
            .I(\c0.n5182 ));
    InMux I__2900 (
            .O(N__17758),
            .I(N__17755));
    LocalMux I__2899 (
            .O(N__17755),
            .I(N__17751));
    InMux I__2898 (
            .O(N__17754),
            .I(N__17748));
    Odrv12 I__2897 (
            .O(N__17751),
            .I(\c0.n5147 ));
    LocalMux I__2896 (
            .O(N__17748),
            .I(\c0.n5147 ));
    CascadeMux I__2895 (
            .O(N__17743),
            .I(\c0.n5182_cascade_ ));
    InMux I__2894 (
            .O(N__17740),
            .I(N__17737));
    LocalMux I__2893 (
            .O(N__17737),
            .I(\c0.n40 ));
    CascadeMux I__2892 (
            .O(N__17734),
            .I(N__17729));
    CascadeMux I__2891 (
            .O(N__17733),
            .I(N__17726));
    InMux I__2890 (
            .O(N__17732),
            .I(N__17722));
    InMux I__2889 (
            .O(N__17729),
            .I(N__17717));
    InMux I__2888 (
            .O(N__17726),
            .I(N__17717));
    InMux I__2887 (
            .O(N__17725),
            .I(N__17714));
    LocalMux I__2886 (
            .O(N__17722),
            .I(N__17711));
    LocalMux I__2885 (
            .O(N__17717),
            .I(N__17708));
    LocalMux I__2884 (
            .O(N__17714),
            .I(\c0.data_in_field_119 ));
    Odrv4 I__2883 (
            .O(N__17711),
            .I(\c0.data_in_field_119 ));
    Odrv12 I__2882 (
            .O(N__17708),
            .I(\c0.data_in_field_119 ));
    InMux I__2881 (
            .O(N__17701),
            .I(N__17698));
    LocalMux I__2880 (
            .O(N__17698),
            .I(\c0.n29 ));
    InMux I__2879 (
            .O(N__17695),
            .I(N__17692));
    LocalMux I__2878 (
            .O(N__17692),
            .I(N__17689));
    Odrv4 I__2877 (
            .O(N__17689),
            .I(\c0.n20_adj_1906 ));
    InMux I__2876 (
            .O(N__17686),
            .I(N__17682));
    InMux I__2875 (
            .O(N__17685),
            .I(N__17679));
    LocalMux I__2874 (
            .O(N__17682),
            .I(N__17676));
    LocalMux I__2873 (
            .O(N__17679),
            .I(N__17673));
    Span4Mux_v I__2872 (
            .O(N__17676),
            .I(N__17670));
    Span4Mux_h I__2871 (
            .O(N__17673),
            .I(N__17666));
    Span4Mux_v I__2870 (
            .O(N__17670),
            .I(N__17663));
    InMux I__2869 (
            .O(N__17669),
            .I(N__17660));
    Odrv4 I__2868 (
            .O(N__17666),
            .I(data_in_4_3));
    Odrv4 I__2867 (
            .O(N__17663),
            .I(data_in_4_3));
    LocalMux I__2866 (
            .O(N__17660),
            .I(data_in_4_3));
    InMux I__2865 (
            .O(N__17653),
            .I(N__17650));
    LocalMux I__2864 (
            .O(N__17650),
            .I(N__17647));
    Span4Mux_h I__2863 (
            .O(N__17647),
            .I(N__17644));
    Span4Mux_s1_h I__2862 (
            .O(N__17644),
            .I(N__17641));
    Odrv4 I__2861 (
            .O(N__17641),
            .I(\c0.n15_adj_1894 ));
    CascadeMux I__2860 (
            .O(N__17638),
            .I(\c0.n16_adj_1893_cascade_ ));
    InMux I__2859 (
            .O(N__17635),
            .I(N__17632));
    LocalMux I__2858 (
            .O(N__17632),
            .I(N__17629));
    Odrv4 I__2857 (
            .O(N__17629),
            .I(\c0.n22_adj_1930 ));
    CascadeMux I__2856 (
            .O(N__17626),
            .I(N__17623));
    InMux I__2855 (
            .O(N__17623),
            .I(N__17620));
    LocalMux I__2854 (
            .O(N__17620),
            .I(N__17617));
    Odrv4 I__2853 (
            .O(N__17617),
            .I(\c0.n2058 ));
    CascadeMux I__2852 (
            .O(N__17614),
            .I(\c0.n5096_cascade_ ));
    CascadeMux I__2851 (
            .O(N__17611),
            .I(\c0.n1785_cascade_ ));
    InMux I__2850 (
            .O(N__17608),
            .I(N__17605));
    LocalMux I__2849 (
            .O(N__17605),
            .I(N__17602));
    Odrv4 I__2848 (
            .O(N__17602),
            .I(\c0.n22 ));
    CascadeMux I__2847 (
            .O(N__17599),
            .I(N__17596));
    InMux I__2846 (
            .O(N__17596),
            .I(N__17591));
    InMux I__2845 (
            .O(N__17595),
            .I(N__17588));
    InMux I__2844 (
            .O(N__17594),
            .I(N__17585));
    LocalMux I__2843 (
            .O(N__17591),
            .I(data_in_13_5));
    LocalMux I__2842 (
            .O(N__17588),
            .I(data_in_13_5));
    LocalMux I__2841 (
            .O(N__17585),
            .I(data_in_13_5));
    InMux I__2840 (
            .O(N__17578),
            .I(N__17575));
    LocalMux I__2839 (
            .O(N__17575),
            .I(N__17572));
    Sp12to4 I__2838 (
            .O(N__17572),
            .I(N__17569));
    Odrv12 I__2837 (
            .O(N__17569),
            .I(\c0.n5150 ));
    InMux I__2836 (
            .O(N__17566),
            .I(N__17563));
    LocalMux I__2835 (
            .O(N__17563),
            .I(N__17556));
    InMux I__2834 (
            .O(N__17562),
            .I(N__17547));
    InMux I__2833 (
            .O(N__17561),
            .I(N__17547));
    InMux I__2832 (
            .O(N__17560),
            .I(N__17547));
    InMux I__2831 (
            .O(N__17559),
            .I(N__17547));
    Odrv12 I__2830 (
            .O(N__17556),
            .I(\c0.data_in_field_109 ));
    LocalMux I__2829 (
            .O(N__17547),
            .I(\c0.data_in_field_109 ));
    CascadeMux I__2828 (
            .O(N__17542),
            .I(\c0.n26_adj_1915_cascade_ ));
    InMux I__2827 (
            .O(N__17539),
            .I(N__17536));
    LocalMux I__2826 (
            .O(N__17536),
            .I(N__17531));
    InMux I__2825 (
            .O(N__17535),
            .I(N__17528));
    CascadeMux I__2824 (
            .O(N__17534),
            .I(N__17525));
    Span4Mux_h I__2823 (
            .O(N__17531),
            .I(N__17522));
    LocalMux I__2822 (
            .O(N__17528),
            .I(N__17519));
    InMux I__2821 (
            .O(N__17525),
            .I(N__17516));
    Odrv4 I__2820 (
            .O(N__17522),
            .I(data_in_17_3));
    Odrv4 I__2819 (
            .O(N__17519),
            .I(data_in_17_3));
    LocalMux I__2818 (
            .O(N__17516),
            .I(data_in_17_3));
    InMux I__2817 (
            .O(N__17509),
            .I(N__17503));
    CascadeMux I__2816 (
            .O(N__17508),
            .I(N__17500));
    InMux I__2815 (
            .O(N__17507),
            .I(N__17496));
    InMux I__2814 (
            .O(N__17506),
            .I(N__17493));
    LocalMux I__2813 (
            .O(N__17503),
            .I(N__17490));
    InMux I__2812 (
            .O(N__17500),
            .I(N__17487));
    InMux I__2811 (
            .O(N__17499),
            .I(N__17484));
    LocalMux I__2810 (
            .O(N__17496),
            .I(N__17481));
    LocalMux I__2809 (
            .O(N__17493),
            .I(N__17478));
    Span4Mux_v I__2808 (
            .O(N__17490),
            .I(N__17473));
    LocalMux I__2807 (
            .O(N__17487),
            .I(N__17473));
    LocalMux I__2806 (
            .O(N__17484),
            .I(\c0.data_in_field_71 ));
    Odrv4 I__2805 (
            .O(N__17481),
            .I(\c0.data_in_field_71 ));
    Odrv12 I__2804 (
            .O(N__17478),
            .I(\c0.data_in_field_71 ));
    Odrv4 I__2803 (
            .O(N__17473),
            .I(\c0.data_in_field_71 ));
    CascadeMux I__2802 (
            .O(N__17464),
            .I(\c0.n26_cascade_ ));
    InMux I__2801 (
            .O(N__17461),
            .I(N__17458));
    LocalMux I__2800 (
            .O(N__17458),
            .I(\c0.n27_adj_1919 ));
    InMux I__2799 (
            .O(N__17455),
            .I(N__17452));
    LocalMux I__2798 (
            .O(N__17452),
            .I(\c0.n5250 ));
    CascadeMux I__2797 (
            .O(N__17449),
            .I(\c0.n28_adj_1917_cascade_ ));
    InMux I__2796 (
            .O(N__17446),
            .I(N__17443));
    LocalMux I__2795 (
            .O(N__17443),
            .I(\c0.n26_adj_1939 ));
    InMux I__2794 (
            .O(N__17440),
            .I(N__17437));
    LocalMux I__2793 (
            .O(N__17437),
            .I(N__17432));
    CascadeMux I__2792 (
            .O(N__17436),
            .I(N__17429));
    InMux I__2791 (
            .O(N__17435),
            .I(N__17426));
    Span4Mux_v I__2790 (
            .O(N__17432),
            .I(N__17423));
    InMux I__2789 (
            .O(N__17429),
            .I(N__17418));
    LocalMux I__2788 (
            .O(N__17426),
            .I(N__17413));
    Span4Mux_h I__2787 (
            .O(N__17423),
            .I(N__17413));
    InMux I__2786 (
            .O(N__17422),
            .I(N__17408));
    InMux I__2785 (
            .O(N__17421),
            .I(N__17408));
    LocalMux I__2784 (
            .O(N__17418),
            .I(\c0.data_in_field_41 ));
    Odrv4 I__2783 (
            .O(N__17413),
            .I(\c0.data_in_field_41 ));
    LocalMux I__2782 (
            .O(N__17408),
            .I(\c0.data_in_field_41 ));
    CascadeMux I__2781 (
            .O(N__17401),
            .I(\c0.n14_cascade_ ));
    InMux I__2780 (
            .O(N__17398),
            .I(N__17394));
    InMux I__2779 (
            .O(N__17397),
            .I(N__17391));
    LocalMux I__2778 (
            .O(N__17394),
            .I(\c0.data_in_frame_18_2 ));
    LocalMux I__2777 (
            .O(N__17391),
            .I(\c0.data_in_frame_18_2 ));
    CascadeMux I__2776 (
            .O(N__17386),
            .I(N__17383));
    InMux I__2775 (
            .O(N__17383),
            .I(N__17380));
    LocalMux I__2774 (
            .O(N__17380),
            .I(N__17377));
    Span4Mux_h I__2773 (
            .O(N__17377),
            .I(N__17374));
    Odrv4 I__2772 (
            .O(N__17374),
            .I(\c0.n5965 ));
    CascadeMux I__2771 (
            .O(N__17371),
            .I(N__17367));
    InMux I__2770 (
            .O(N__17370),
            .I(N__17364));
    InMux I__2769 (
            .O(N__17367),
            .I(N__17361));
    LocalMux I__2768 (
            .O(N__17364),
            .I(N__17356));
    LocalMux I__2767 (
            .O(N__17361),
            .I(N__17353));
    InMux I__2766 (
            .O(N__17360),
            .I(N__17350));
    InMux I__2765 (
            .O(N__17359),
            .I(N__17347));
    Span4Mux_v I__2764 (
            .O(N__17356),
            .I(N__17344));
    Span4Mux_v I__2763 (
            .O(N__17353),
            .I(N__17341));
    LocalMux I__2762 (
            .O(N__17350),
            .I(data_in_19_6));
    LocalMux I__2761 (
            .O(N__17347),
            .I(data_in_19_6));
    Odrv4 I__2760 (
            .O(N__17344),
            .I(data_in_19_6));
    Odrv4 I__2759 (
            .O(N__17341),
            .I(data_in_19_6));
    CascadeMux I__2758 (
            .O(N__17332),
            .I(\c0.n22_adj_1901_cascade_ ));
    InMux I__2757 (
            .O(N__17329),
            .I(N__17326));
    LocalMux I__2756 (
            .O(N__17326),
            .I(\c0.n23_adj_1932 ));
    CascadeMux I__2755 (
            .O(N__17323),
            .I(\c0.n30_adj_1940_cascade_ ));
    InMux I__2754 (
            .O(N__17320),
            .I(N__17310));
    InMux I__2753 (
            .O(N__17319),
            .I(N__17310));
    InMux I__2752 (
            .O(N__17318),
            .I(N__17310));
    InMux I__2751 (
            .O(N__17317),
            .I(N__17307));
    LocalMux I__2750 (
            .O(N__17310),
            .I(\c0.n3563 ));
    LocalMux I__2749 (
            .O(N__17307),
            .I(\c0.n3563 ));
    InMux I__2748 (
            .O(N__17302),
            .I(N__17299));
    LocalMux I__2747 (
            .O(N__17299),
            .I(\c0.n5280 ));
    InMux I__2746 (
            .O(N__17296),
            .I(N__17293));
    LocalMux I__2745 (
            .O(N__17293),
            .I(\c0.n5277 ));
    InMux I__2744 (
            .O(N__17290),
            .I(N__17287));
    LocalMux I__2743 (
            .O(N__17287),
            .I(\c0.n25_adj_1941 ));
    InMux I__2742 (
            .O(N__17284),
            .I(N__17281));
    LocalMux I__2741 (
            .O(N__17281),
            .I(N__17278));
    Span4Mux_h I__2740 (
            .O(N__17278),
            .I(N__17274));
    InMux I__2739 (
            .O(N__17277),
            .I(N__17271));
    Odrv4 I__2738 (
            .O(N__17274),
            .I(\c0.n5072 ));
    LocalMux I__2737 (
            .O(N__17271),
            .I(\c0.n5072 ));
    InMux I__2736 (
            .O(N__17266),
            .I(N__17260));
    InMux I__2735 (
            .O(N__17265),
            .I(N__17260));
    LocalMux I__2734 (
            .O(N__17260),
            .I(r_Tx_Data_3));
    InMux I__2733 (
            .O(N__17257),
            .I(N__17253));
    InMux I__2732 (
            .O(N__17256),
            .I(N__17250));
    LocalMux I__2731 (
            .O(N__17253),
            .I(N__17247));
    LocalMux I__2730 (
            .O(N__17250),
            .I(r_Tx_Data_2));
    Odrv4 I__2729 (
            .O(N__17247),
            .I(r_Tx_Data_2));
    CascadeMux I__2728 (
            .O(N__17242),
            .I(N__17239));
    InMux I__2727 (
            .O(N__17239),
            .I(N__17230));
    CascadeMux I__2726 (
            .O(N__17238),
            .I(N__17227));
    InMux I__2725 (
            .O(N__17237),
            .I(N__17224));
    InMux I__2724 (
            .O(N__17236),
            .I(N__17221));
    InMux I__2723 (
            .O(N__17235),
            .I(N__17218));
    InMux I__2722 (
            .O(N__17234),
            .I(N__17215));
    InMux I__2721 (
            .O(N__17233),
            .I(N__17212));
    LocalMux I__2720 (
            .O(N__17230),
            .I(N__17209));
    InMux I__2719 (
            .O(N__17227),
            .I(N__17206));
    LocalMux I__2718 (
            .O(N__17224),
            .I(r_Bit_Index_1));
    LocalMux I__2717 (
            .O(N__17221),
            .I(r_Bit_Index_1));
    LocalMux I__2716 (
            .O(N__17218),
            .I(r_Bit_Index_1));
    LocalMux I__2715 (
            .O(N__17215),
            .I(r_Bit_Index_1));
    LocalMux I__2714 (
            .O(N__17212),
            .I(r_Bit_Index_1));
    Odrv4 I__2713 (
            .O(N__17209),
            .I(r_Bit_Index_1));
    LocalMux I__2712 (
            .O(N__17206),
            .I(r_Bit_Index_1));
    CascadeMux I__2711 (
            .O(N__17191),
            .I(N__17187));
    InMux I__2710 (
            .O(N__17190),
            .I(N__17180));
    InMux I__2709 (
            .O(N__17187),
            .I(N__17173));
    InMux I__2708 (
            .O(N__17186),
            .I(N__17173));
    InMux I__2707 (
            .O(N__17185),
            .I(N__17173));
    InMux I__2706 (
            .O(N__17184),
            .I(N__17170));
    InMux I__2705 (
            .O(N__17183),
            .I(N__17167));
    LocalMux I__2704 (
            .O(N__17180),
            .I(r_Bit_Index_0));
    LocalMux I__2703 (
            .O(N__17173),
            .I(r_Bit_Index_0));
    LocalMux I__2702 (
            .O(N__17170),
            .I(r_Bit_Index_0));
    LocalMux I__2701 (
            .O(N__17167),
            .I(r_Bit_Index_0));
    InMux I__2700 (
            .O(N__17158),
            .I(N__17155));
    LocalMux I__2699 (
            .O(N__17155),
            .I(\c0.tx.n5719 ));
    InMux I__2698 (
            .O(N__17152),
            .I(N__17147));
    InMux I__2697 (
            .O(N__17151),
            .I(N__17144));
    InMux I__2696 (
            .O(N__17150),
            .I(N__17141));
    LocalMux I__2695 (
            .O(N__17147),
            .I(r_Bit_Index_2));
    LocalMux I__2694 (
            .O(N__17144),
            .I(r_Bit_Index_2));
    LocalMux I__2693 (
            .O(N__17141),
            .I(r_Bit_Index_2));
    InMux I__2692 (
            .O(N__17134),
            .I(N__17131));
    LocalMux I__2691 (
            .O(N__17131),
            .I(\c0.tx.n5716 ));
    InMux I__2690 (
            .O(N__17128),
            .I(N__17125));
    LocalMux I__2689 (
            .O(N__17125),
            .I(\c0.tx.n5722 ));
    InMux I__2688 (
            .O(N__17122),
            .I(N__17111));
    InMux I__2687 (
            .O(N__17121),
            .I(N__17111));
    InMux I__2686 (
            .O(N__17120),
            .I(N__17104));
    InMux I__2685 (
            .O(N__17119),
            .I(N__17104));
    InMux I__2684 (
            .O(N__17118),
            .I(N__17104));
    InMux I__2683 (
            .O(N__17117),
            .I(N__17101));
    InMux I__2682 (
            .O(N__17116),
            .I(N__17094));
    LocalMux I__2681 (
            .O(N__17111),
            .I(N__17091));
    LocalMux I__2680 (
            .O(N__17104),
            .I(N__17086));
    LocalMux I__2679 (
            .O(N__17101),
            .I(N__17086));
    InMux I__2678 (
            .O(N__17100),
            .I(N__17081));
    InMux I__2677 (
            .O(N__17099),
            .I(N__17081));
    InMux I__2676 (
            .O(N__17098),
            .I(N__17076));
    InMux I__2675 (
            .O(N__17097),
            .I(N__17076));
    LocalMux I__2674 (
            .O(N__17094),
            .I(r_SM_Main_1));
    Odrv4 I__2673 (
            .O(N__17091),
            .I(r_SM_Main_1));
    Odrv4 I__2672 (
            .O(N__17086),
            .I(r_SM_Main_1));
    LocalMux I__2671 (
            .O(N__17081),
            .I(r_SM_Main_1));
    LocalMux I__2670 (
            .O(N__17076),
            .I(r_SM_Main_1));
    CascadeMux I__2669 (
            .O(N__17065),
            .I(\c0.tx.o_Tx_Serial_N_1798_cascade_ ));
    InMux I__2668 (
            .O(N__17062),
            .I(N__17055));
    InMux I__2667 (
            .O(N__17061),
            .I(N__17052));
    CascadeMux I__2666 (
            .O(N__17060),
            .I(N__17046));
    InMux I__2665 (
            .O(N__17059),
            .I(N__17041));
    InMux I__2664 (
            .O(N__17058),
            .I(N__17038));
    LocalMux I__2663 (
            .O(N__17055),
            .I(N__17035));
    LocalMux I__2662 (
            .O(N__17052),
            .I(N__17032));
    InMux I__2661 (
            .O(N__17051),
            .I(N__17029));
    InMux I__2660 (
            .O(N__17050),
            .I(N__17026));
    InMux I__2659 (
            .O(N__17049),
            .I(N__17017));
    InMux I__2658 (
            .O(N__17046),
            .I(N__17017));
    InMux I__2657 (
            .O(N__17045),
            .I(N__17017));
    InMux I__2656 (
            .O(N__17044),
            .I(N__17017));
    LocalMux I__2655 (
            .O(N__17041),
            .I(r_SM_Main_0));
    LocalMux I__2654 (
            .O(N__17038),
            .I(r_SM_Main_0));
    Odrv4 I__2653 (
            .O(N__17035),
            .I(r_SM_Main_0));
    Odrv4 I__2652 (
            .O(N__17032),
            .I(r_SM_Main_0));
    LocalMux I__2651 (
            .O(N__17029),
            .I(r_SM_Main_0));
    LocalMux I__2650 (
            .O(N__17026),
            .I(r_SM_Main_0));
    LocalMux I__2649 (
            .O(N__17017),
            .I(r_SM_Main_0));
    CascadeMux I__2648 (
            .O(N__17002),
            .I(N__16993));
    CascadeMux I__2647 (
            .O(N__17001),
            .I(N__16989));
    CascadeMux I__2646 (
            .O(N__17000),
            .I(N__16986));
    CascadeMux I__2645 (
            .O(N__16999),
            .I(N__16980));
    CascadeMux I__2644 (
            .O(N__16998),
            .I(N__16974));
    CascadeMux I__2643 (
            .O(N__16997),
            .I(N__16969));
    InMux I__2642 (
            .O(N__16996),
            .I(N__16962));
    InMux I__2641 (
            .O(N__16993),
            .I(N__16962));
    InMux I__2640 (
            .O(N__16992),
            .I(N__16959));
    InMux I__2639 (
            .O(N__16989),
            .I(N__16950));
    InMux I__2638 (
            .O(N__16986),
            .I(N__16950));
    InMux I__2637 (
            .O(N__16985),
            .I(N__16950));
    InMux I__2636 (
            .O(N__16984),
            .I(N__16950));
    CascadeMux I__2635 (
            .O(N__16983),
            .I(N__16946));
    InMux I__2634 (
            .O(N__16980),
            .I(N__16937));
    InMux I__2633 (
            .O(N__16979),
            .I(N__16937));
    InMux I__2632 (
            .O(N__16978),
            .I(N__16937));
    InMux I__2631 (
            .O(N__16977),
            .I(N__16937));
    InMux I__2630 (
            .O(N__16974),
            .I(N__16932));
    InMux I__2629 (
            .O(N__16973),
            .I(N__16932));
    InMux I__2628 (
            .O(N__16972),
            .I(N__16923));
    InMux I__2627 (
            .O(N__16969),
            .I(N__16923));
    InMux I__2626 (
            .O(N__16968),
            .I(N__16923));
    InMux I__2625 (
            .O(N__16967),
            .I(N__16923));
    LocalMux I__2624 (
            .O(N__16962),
            .I(N__16920));
    LocalMux I__2623 (
            .O(N__16959),
            .I(N__16915));
    LocalMux I__2622 (
            .O(N__16950),
            .I(N__16915));
    InMux I__2621 (
            .O(N__16949),
            .I(N__16912));
    InMux I__2620 (
            .O(N__16946),
            .I(N__16909));
    LocalMux I__2619 (
            .O(N__16937),
            .I(r_SM_Main_2));
    LocalMux I__2618 (
            .O(N__16932),
            .I(r_SM_Main_2));
    LocalMux I__2617 (
            .O(N__16923),
            .I(r_SM_Main_2));
    Odrv4 I__2616 (
            .O(N__16920),
            .I(r_SM_Main_2));
    Odrv12 I__2615 (
            .O(N__16915),
            .I(r_SM_Main_2));
    LocalMux I__2614 (
            .O(N__16912),
            .I(r_SM_Main_2));
    LocalMux I__2613 (
            .O(N__16909),
            .I(r_SM_Main_2));
    CascadeMux I__2612 (
            .O(N__16894),
            .I(\c0.tx.n3_cascade_ ));
    InMux I__2611 (
            .O(N__16891),
            .I(N__16887));
    IoInMux I__2610 (
            .O(N__16890),
            .I(N__16884));
    LocalMux I__2609 (
            .O(N__16887),
            .I(N__16879));
    LocalMux I__2608 (
            .O(N__16884),
            .I(N__16879));
    Span4Mux_s3_v I__2607 (
            .O(N__16879),
            .I(N__16876));
    Span4Mux_h I__2606 (
            .O(N__16876),
            .I(N__16873));
    Span4Mux_v I__2605 (
            .O(N__16873),
            .I(N__16870));
    Span4Mux_v I__2604 (
            .O(N__16870),
            .I(N__16866));
    InMux I__2603 (
            .O(N__16869),
            .I(N__16863));
    Odrv4 I__2602 (
            .O(N__16866),
            .I(tx_o));
    LocalMux I__2601 (
            .O(N__16863),
            .I(tx_o));
    CascadeMux I__2600 (
            .O(N__16858),
            .I(N__16855));
    InMux I__2599 (
            .O(N__16855),
            .I(N__16852));
    LocalMux I__2598 (
            .O(N__16852),
            .I(\c0.n2018 ));
    InMux I__2597 (
            .O(N__16849),
            .I(N__16846));
    LocalMux I__2596 (
            .O(N__16846),
            .I(\c0.n5519 ));
    InMux I__2595 (
            .O(N__16843),
            .I(N__16840));
    LocalMux I__2594 (
            .O(N__16840),
            .I(N__16837));
    Span4Mux_h I__2593 (
            .O(N__16837),
            .I(N__16834));
    Odrv4 I__2592 (
            .O(N__16834),
            .I(\c0.n5980 ));
    InMux I__2591 (
            .O(N__16831),
            .I(N__16828));
    LocalMux I__2590 (
            .O(N__16828),
            .I(N__16824));
    InMux I__2589 (
            .O(N__16827),
            .I(N__16821));
    Span4Mux_h I__2588 (
            .O(N__16824),
            .I(N__16818));
    LocalMux I__2587 (
            .O(N__16821),
            .I(r_Tx_Data_4));
    Odrv4 I__2586 (
            .O(N__16818),
            .I(r_Tx_Data_4));
    CascadeMux I__2585 (
            .O(N__16813),
            .I(\c0.tx.n5713_cascade_ ));
    InMux I__2584 (
            .O(N__16810),
            .I(N__16804));
    InMux I__2583 (
            .O(N__16809),
            .I(N__16801));
    InMux I__2582 (
            .O(N__16808),
            .I(N__16798));
    InMux I__2581 (
            .O(N__16807),
            .I(N__16793));
    LocalMux I__2580 (
            .O(N__16804),
            .I(N__16790));
    LocalMux I__2579 (
            .O(N__16801),
            .I(N__16787));
    LocalMux I__2578 (
            .O(N__16798),
            .I(N__16784));
    InMux I__2577 (
            .O(N__16797),
            .I(N__16779));
    InMux I__2576 (
            .O(N__16796),
            .I(N__16779));
    LocalMux I__2575 (
            .O(N__16793),
            .I(N__16770));
    Span4Mux_v I__2574 (
            .O(N__16790),
            .I(N__16770));
    Span4Mux_v I__2573 (
            .O(N__16787),
            .I(N__16770));
    Span4Mux_v I__2572 (
            .O(N__16784),
            .I(N__16770));
    LocalMux I__2571 (
            .O(N__16779),
            .I(data_out_11_1));
    Odrv4 I__2570 (
            .O(N__16770),
            .I(data_out_11_1));
    CascadeMux I__2569 (
            .O(N__16765),
            .I(N__16762));
    InMux I__2568 (
            .O(N__16762),
            .I(N__16759));
    LocalMux I__2567 (
            .O(N__16759),
            .I(\c0.n9_adj_1880 ));
    CascadeMux I__2566 (
            .O(N__16756),
            .I(N__16753));
    InMux I__2565 (
            .O(N__16753),
            .I(N__16750));
    LocalMux I__2564 (
            .O(N__16750),
            .I(N__16747));
    Odrv4 I__2563 (
            .O(N__16747),
            .I(\c0.n9_adj_1890 ));
    InMux I__2562 (
            .O(N__16744),
            .I(N__16741));
    LocalMux I__2561 (
            .O(N__16741),
            .I(N__16738));
    Odrv12 I__2560 (
            .O(N__16738),
            .I(\c0.n5489 ));
    CascadeMux I__2559 (
            .O(N__16735),
            .I(\c0.n991_cascade_ ));
    CascadeMux I__2558 (
            .O(N__16732),
            .I(tx_data_5_N_keep_cascade_));
    InMux I__2557 (
            .O(N__16729),
            .I(N__16723));
    InMux I__2556 (
            .O(N__16728),
            .I(N__16723));
    LocalMux I__2555 (
            .O(N__16723),
            .I(r_Tx_Data_5));
    InMux I__2554 (
            .O(N__16720),
            .I(N__16717));
    LocalMux I__2553 (
            .O(N__16717),
            .I(N__16714));
    Odrv4 I__2552 (
            .O(N__16714),
            .I(tx_data_3_N_keep));
    InMux I__2551 (
            .O(N__16711),
            .I(N__16707));
    CascadeMux I__2550 (
            .O(N__16710),
            .I(N__16704));
    LocalMux I__2549 (
            .O(N__16707),
            .I(N__16700));
    InMux I__2548 (
            .O(N__16704),
            .I(N__16695));
    InMux I__2547 (
            .O(N__16703),
            .I(N__16695));
    Odrv4 I__2546 (
            .O(N__16700),
            .I(n5135));
    LocalMux I__2545 (
            .O(N__16695),
            .I(n5135));
    InMux I__2544 (
            .O(N__16690),
            .I(N__16687));
    LocalMux I__2543 (
            .O(N__16687),
            .I(n5117));
    CascadeMux I__2542 (
            .O(N__16684),
            .I(n5117_cascade_));
    InMux I__2541 (
            .O(N__16681),
            .I(N__16674));
    InMux I__2540 (
            .O(N__16680),
            .I(N__16658));
    InMux I__2539 (
            .O(N__16679),
            .I(N__16658));
    InMux I__2538 (
            .O(N__16678),
            .I(N__16655));
    InMux I__2537 (
            .O(N__16677),
            .I(N__16652));
    LocalMux I__2536 (
            .O(N__16674),
            .I(N__16649));
    InMux I__2535 (
            .O(N__16673),
            .I(N__16646));
    InMux I__2534 (
            .O(N__16672),
            .I(N__16643));
    InMux I__2533 (
            .O(N__16671),
            .I(N__16640));
    InMux I__2532 (
            .O(N__16670),
            .I(N__16631));
    InMux I__2531 (
            .O(N__16669),
            .I(N__16631));
    InMux I__2530 (
            .O(N__16668),
            .I(N__16631));
    InMux I__2529 (
            .O(N__16667),
            .I(N__16631));
    InMux I__2528 (
            .O(N__16666),
            .I(N__16626));
    InMux I__2527 (
            .O(N__16665),
            .I(N__16626));
    InMux I__2526 (
            .O(N__16664),
            .I(N__16621));
    InMux I__2525 (
            .O(N__16663),
            .I(N__16621));
    LocalMux I__2524 (
            .O(N__16658),
            .I(n4316));
    LocalMux I__2523 (
            .O(N__16655),
            .I(n4316));
    LocalMux I__2522 (
            .O(N__16652),
            .I(n4316));
    Odrv4 I__2521 (
            .O(N__16649),
            .I(n4316));
    LocalMux I__2520 (
            .O(N__16646),
            .I(n4316));
    LocalMux I__2519 (
            .O(N__16643),
            .I(n4316));
    LocalMux I__2518 (
            .O(N__16640),
            .I(n4316));
    LocalMux I__2517 (
            .O(N__16631),
            .I(n4316));
    LocalMux I__2516 (
            .O(N__16626),
            .I(n4316));
    LocalMux I__2515 (
            .O(N__16621),
            .I(n4316));
    CascadeMux I__2514 (
            .O(N__16600),
            .I(N__16596));
    InMux I__2513 (
            .O(N__16599),
            .I(N__16591));
    InMux I__2512 (
            .O(N__16596),
            .I(N__16591));
    LocalMux I__2511 (
            .O(N__16591),
            .I(data_out_19_5));
    InMux I__2510 (
            .O(N__16588),
            .I(N__16585));
    LocalMux I__2509 (
            .O(N__16585),
            .I(tx_data_2_N_keep));
    InMux I__2508 (
            .O(N__16582),
            .I(N__16576));
    InMux I__2507 (
            .O(N__16581),
            .I(N__16571));
    InMux I__2506 (
            .O(N__16580),
            .I(N__16571));
    InMux I__2505 (
            .O(N__16579),
            .I(N__16567));
    LocalMux I__2504 (
            .O(N__16576),
            .I(N__16562));
    LocalMux I__2503 (
            .O(N__16571),
            .I(N__16559));
    InMux I__2502 (
            .O(N__16570),
            .I(N__16555));
    LocalMux I__2501 (
            .O(N__16567),
            .I(N__16552));
    CascadeMux I__2500 (
            .O(N__16566),
            .I(N__16549));
    InMux I__2499 (
            .O(N__16565),
            .I(N__16546));
    Span4Mux_v I__2498 (
            .O(N__16562),
            .I(N__16541));
    Span4Mux_v I__2497 (
            .O(N__16559),
            .I(N__16541));
    InMux I__2496 (
            .O(N__16558),
            .I(N__16538));
    LocalMux I__2495 (
            .O(N__16555),
            .I(N__16533));
    Span4Mux_h I__2494 (
            .O(N__16552),
            .I(N__16533));
    InMux I__2493 (
            .O(N__16549),
            .I(N__16530));
    LocalMux I__2492 (
            .O(N__16546),
            .I(data_out_11_3));
    Odrv4 I__2491 (
            .O(N__16541),
            .I(data_out_11_3));
    LocalMux I__2490 (
            .O(N__16538),
            .I(data_out_11_3));
    Odrv4 I__2489 (
            .O(N__16533),
            .I(data_out_11_3));
    LocalMux I__2488 (
            .O(N__16530),
            .I(data_out_11_3));
    InMux I__2487 (
            .O(N__16519),
            .I(N__16516));
    LocalMux I__2486 (
            .O(N__16516),
            .I(N__16509));
    CascadeMux I__2485 (
            .O(N__16515),
            .I(N__16506));
    CascadeMux I__2484 (
            .O(N__16514),
            .I(N__16503));
    CascadeMux I__2483 (
            .O(N__16513),
            .I(N__16500));
    InMux I__2482 (
            .O(N__16512),
            .I(N__16497));
    Span4Mux_v I__2481 (
            .O(N__16509),
            .I(N__16494));
    InMux I__2480 (
            .O(N__16506),
            .I(N__16489));
    InMux I__2479 (
            .O(N__16503),
            .I(N__16489));
    InMux I__2478 (
            .O(N__16500),
            .I(N__16486));
    LocalMux I__2477 (
            .O(N__16497),
            .I(data_out_11_2));
    Odrv4 I__2476 (
            .O(N__16494),
            .I(data_out_11_2));
    LocalMux I__2475 (
            .O(N__16489),
            .I(data_out_11_2));
    LocalMux I__2474 (
            .O(N__16486),
            .I(data_out_11_2));
    CascadeMux I__2473 (
            .O(N__16477),
            .I(\c0.n1805_cascade_ ));
    InMux I__2472 (
            .O(N__16474),
            .I(N__16471));
    LocalMux I__2471 (
            .O(N__16471),
            .I(N__16466));
    InMux I__2470 (
            .O(N__16470),
            .I(N__16463));
    InMux I__2469 (
            .O(N__16469),
            .I(N__16460));
    Span4Mux_h I__2468 (
            .O(N__16466),
            .I(N__16457));
    LocalMux I__2467 (
            .O(N__16463),
            .I(n135));
    LocalMux I__2466 (
            .O(N__16460),
            .I(n135));
    Odrv4 I__2465 (
            .O(N__16457),
            .I(n135));
    InMux I__2464 (
            .O(N__16450),
            .I(N__16447));
    LocalMux I__2463 (
            .O(N__16447),
            .I(\c0.n1805 ));
    InMux I__2462 (
            .O(N__16444),
            .I(N__16441));
    LocalMux I__2461 (
            .O(N__16441),
            .I(N__16438));
    Odrv12 I__2460 (
            .O(N__16438),
            .I(n5173));
    InMux I__2459 (
            .O(N__16435),
            .I(N__16427));
    InMux I__2458 (
            .O(N__16434),
            .I(N__16420));
    InMux I__2457 (
            .O(N__16433),
            .I(N__16420));
    InMux I__2456 (
            .O(N__16432),
            .I(N__16420));
    InMux I__2455 (
            .O(N__16431),
            .I(N__16417));
    InMux I__2454 (
            .O(N__16430),
            .I(N__16412));
    LocalMux I__2453 (
            .O(N__16427),
            .I(N__16407));
    LocalMux I__2452 (
            .O(N__16420),
            .I(N__16407));
    LocalMux I__2451 (
            .O(N__16417),
            .I(N__16404));
    InMux I__2450 (
            .O(N__16416),
            .I(N__16401));
    InMux I__2449 (
            .O(N__16415),
            .I(N__16398));
    LocalMux I__2448 (
            .O(N__16412),
            .I(N__16395));
    Span4Mux_v I__2447 (
            .O(N__16407),
            .I(N__16392));
    Span4Mux_s2_h I__2446 (
            .O(N__16404),
            .I(N__16389));
    LocalMux I__2445 (
            .O(N__16401),
            .I(data_out_11_7));
    LocalMux I__2444 (
            .O(N__16398),
            .I(data_out_11_7));
    Odrv12 I__2443 (
            .O(N__16395),
            .I(data_out_11_7));
    Odrv4 I__2442 (
            .O(N__16392),
            .I(data_out_11_7));
    Odrv4 I__2441 (
            .O(N__16389),
            .I(data_out_11_7));
    CascadeMux I__2440 (
            .O(N__16378),
            .I(N__16375));
    InMux I__2439 (
            .O(N__16375),
            .I(N__16372));
    LocalMux I__2438 (
            .O(N__16372),
            .I(N__16367));
    InMux I__2437 (
            .O(N__16371),
            .I(N__16364));
    CascadeMux I__2436 (
            .O(N__16370),
            .I(N__16360));
    Span4Mux_h I__2435 (
            .O(N__16367),
            .I(N__16355));
    LocalMux I__2434 (
            .O(N__16364),
            .I(N__16355));
    InMux I__2433 (
            .O(N__16363),
            .I(N__16351));
    InMux I__2432 (
            .O(N__16360),
            .I(N__16348));
    Span4Mux_v I__2431 (
            .O(N__16355),
            .I(N__16345));
    InMux I__2430 (
            .O(N__16354),
            .I(N__16341));
    LocalMux I__2429 (
            .O(N__16351),
            .I(N__16338));
    LocalMux I__2428 (
            .O(N__16348),
            .I(N__16335));
    Span4Mux_s1_h I__2427 (
            .O(N__16345),
            .I(N__16332));
    InMux I__2426 (
            .O(N__16344),
            .I(N__16329));
    LocalMux I__2425 (
            .O(N__16341),
            .I(data_out_10_7));
    Odrv4 I__2424 (
            .O(N__16338),
            .I(data_out_10_7));
    Odrv12 I__2423 (
            .O(N__16335),
            .I(data_out_10_7));
    Odrv4 I__2422 (
            .O(N__16332),
            .I(data_out_10_7));
    LocalMux I__2421 (
            .O(N__16329),
            .I(data_out_10_7));
    InMux I__2420 (
            .O(N__16318),
            .I(N__16315));
    LocalMux I__2419 (
            .O(N__16315),
            .I(N__16312));
    Odrv4 I__2418 (
            .O(N__16312),
            .I(n5079));
    CascadeMux I__2417 (
            .O(N__16309),
            .I(N__16305));
    CascadeMux I__2416 (
            .O(N__16308),
            .I(N__16302));
    InMux I__2415 (
            .O(N__16305),
            .I(N__16299));
    InMux I__2414 (
            .O(N__16302),
            .I(N__16296));
    LocalMux I__2413 (
            .O(N__16299),
            .I(data_out_19_1));
    LocalMux I__2412 (
            .O(N__16296),
            .I(data_out_19_1));
    CascadeMux I__2411 (
            .O(N__16291),
            .I(N__16288));
    InMux I__2410 (
            .O(N__16288),
            .I(N__16285));
    LocalMux I__2409 (
            .O(N__16285),
            .I(N__16280));
    InMux I__2408 (
            .O(N__16284),
            .I(N__16277));
    InMux I__2407 (
            .O(N__16283),
            .I(N__16274));
    Span4Mux_v I__2406 (
            .O(N__16280),
            .I(N__16264));
    LocalMux I__2405 (
            .O(N__16277),
            .I(N__16264));
    LocalMux I__2404 (
            .O(N__16274),
            .I(N__16264));
    InMux I__2403 (
            .O(N__16273),
            .I(N__16261));
    InMux I__2402 (
            .O(N__16272),
            .I(N__16256));
    InMux I__2401 (
            .O(N__16271),
            .I(N__16256));
    Span4Mux_h I__2400 (
            .O(N__16264),
            .I(N__16253));
    LocalMux I__2399 (
            .O(N__16261),
            .I(data_out_11_0));
    LocalMux I__2398 (
            .O(N__16256),
            .I(data_out_11_0));
    Odrv4 I__2397 (
            .O(N__16253),
            .I(data_out_11_0));
    InMux I__2396 (
            .O(N__16246),
            .I(N__16242));
    InMux I__2395 (
            .O(N__16245),
            .I(N__16239));
    LocalMux I__2394 (
            .O(N__16242),
            .I(data_out_18_2));
    LocalMux I__2393 (
            .O(N__16239),
            .I(data_out_18_2));
    CascadeMux I__2392 (
            .O(N__16234),
            .I(N__16231));
    InMux I__2391 (
            .O(N__16231),
            .I(N__16228));
    LocalMux I__2390 (
            .O(N__16228),
            .I(N__16224));
    InMux I__2389 (
            .O(N__16227),
            .I(N__16221));
    Span4Mux_h I__2388 (
            .O(N__16224),
            .I(N__16218));
    LocalMux I__2387 (
            .O(N__16221),
            .I(data_out_19_2));
    Odrv4 I__2386 (
            .O(N__16218),
            .I(data_out_19_2));
    InMux I__2385 (
            .O(N__16213),
            .I(N__16210));
    LocalMux I__2384 (
            .O(N__16210),
            .I(\c0.n2249 ));
    CascadeMux I__2383 (
            .O(N__16207),
            .I(\c0.n5522_cascade_ ));
    InMux I__2382 (
            .O(N__16204),
            .I(N__16201));
    LocalMux I__2381 (
            .O(N__16201),
            .I(n4_adj_1991));
    InMux I__2380 (
            .O(N__16198),
            .I(N__16194));
    InMux I__2379 (
            .O(N__16197),
            .I(N__16191));
    LocalMux I__2378 (
            .O(N__16194),
            .I(data_out_18_5));
    LocalMux I__2377 (
            .O(N__16191),
            .I(data_out_18_5));
    InMux I__2376 (
            .O(N__16186),
            .I(N__16183));
    LocalMux I__2375 (
            .O(N__16183),
            .I(N__16180));
    Odrv12 I__2374 (
            .O(N__16180),
            .I(n4_adj_1994));
    CascadeMux I__2373 (
            .O(N__16177),
            .I(\c0.rx.n2151_cascade_ ));
    CascadeMux I__2372 (
            .O(N__16174),
            .I(n1709_cascade_));
    InMux I__2371 (
            .O(N__16171),
            .I(N__16167));
    InMux I__2370 (
            .O(N__16170),
            .I(N__16164));
    LocalMux I__2369 (
            .O(N__16167),
            .I(N__16161));
    LocalMux I__2368 (
            .O(N__16164),
            .I(n4_adj_1990));
    Odrv4 I__2367 (
            .O(N__16161),
            .I(n4_adj_1990));
    InMux I__2366 (
            .O(N__16156),
            .I(N__16152));
    InMux I__2365 (
            .O(N__16155),
            .I(N__16149));
    LocalMux I__2364 (
            .O(N__16152),
            .I(rx_data_4));
    LocalMux I__2363 (
            .O(N__16149),
            .I(rx_data_4));
    CascadeMux I__2362 (
            .O(N__16144),
            .I(N__16141));
    InMux I__2361 (
            .O(N__16141),
            .I(N__16138));
    LocalMux I__2360 (
            .O(N__16138),
            .I(N__16135));
    Span4Mux_h I__2359 (
            .O(N__16135),
            .I(N__16132));
    Odrv4 I__2358 (
            .O(N__16132),
            .I(n4_adj_1992));
    InMux I__2357 (
            .O(N__16129),
            .I(N__16126));
    LocalMux I__2356 (
            .O(N__16126),
            .I(N__16122));
    InMux I__2355 (
            .O(N__16125),
            .I(N__16119));
    Span4Mux_v I__2354 (
            .O(N__16122),
            .I(N__16116));
    LocalMux I__2353 (
            .O(N__16119),
            .I(\c0.data_in_frame_18_6 ));
    Odrv4 I__2352 (
            .O(N__16116),
            .I(\c0.data_in_frame_18_6 ));
    InMux I__2351 (
            .O(N__16111),
            .I(N__16108));
    LocalMux I__2350 (
            .O(N__16108),
            .I(N__16104));
    InMux I__2349 (
            .O(N__16107),
            .I(N__16099));
    Span4Mux_v I__2348 (
            .O(N__16104),
            .I(N__16096));
    InMux I__2347 (
            .O(N__16103),
            .I(N__16091));
    InMux I__2346 (
            .O(N__16102),
            .I(N__16091));
    LocalMux I__2345 (
            .O(N__16099),
            .I(data_in_2_5));
    Odrv4 I__2344 (
            .O(N__16096),
            .I(data_in_2_5));
    LocalMux I__2343 (
            .O(N__16091),
            .I(data_in_2_5));
    InMux I__2342 (
            .O(N__16084),
            .I(N__16081));
    LocalMux I__2341 (
            .O(N__16081),
            .I(N__16077));
    InMux I__2340 (
            .O(N__16080),
            .I(N__16074));
    Odrv4 I__2339 (
            .O(N__16077),
            .I(rx_data_6));
    LocalMux I__2338 (
            .O(N__16074),
            .I(rx_data_6));
    CascadeMux I__2337 (
            .O(N__16069),
            .I(\c0.n5222_cascade_ ));
    InMux I__2336 (
            .O(N__16066),
            .I(N__16063));
    LocalMux I__2335 (
            .O(N__16063),
            .I(\c0.n42 ));
    CascadeMux I__2334 (
            .O(N__16060),
            .I(\c0.n33_cascade_ ));
    CascadeMux I__2333 (
            .O(N__16057),
            .I(\c0.n2008_cascade_ ));
    CascadeMux I__2332 (
            .O(N__16054),
            .I(\c0.n38_cascade_ ));
    InMux I__2331 (
            .O(N__16051),
            .I(N__16048));
    LocalMux I__2330 (
            .O(N__16048),
            .I(N__16045));
    Span4Mux_s3_h I__2329 (
            .O(N__16045),
            .I(N__16042));
    Odrv4 I__2328 (
            .O(N__16042),
            .I(\c0.n5462 ));
    CascadeMux I__2327 (
            .O(N__16039),
            .I(N__16036));
    InMux I__2326 (
            .O(N__16036),
            .I(N__16030));
    InMux I__2325 (
            .O(N__16035),
            .I(N__16030));
    LocalMux I__2324 (
            .O(N__16030),
            .I(N__16026));
    InMux I__2323 (
            .O(N__16029),
            .I(N__16023));
    Span4Mux_s3_h I__2322 (
            .O(N__16026),
            .I(N__16020));
    LocalMux I__2321 (
            .O(N__16023),
            .I(data_in_12_5));
    Odrv4 I__2320 (
            .O(N__16020),
            .I(data_in_12_5));
    InMux I__2319 (
            .O(N__16015),
            .I(N__16012));
    LocalMux I__2318 (
            .O(N__16012),
            .I(N__16008));
    InMux I__2317 (
            .O(N__16011),
            .I(N__16005));
    Span4Mux_v I__2316 (
            .O(N__16008),
            .I(N__16002));
    LocalMux I__2315 (
            .O(N__16005),
            .I(\c0.data_in_frame_18_0 ));
    Odrv4 I__2314 (
            .O(N__16002),
            .I(\c0.data_in_frame_18_0 ));
    InMux I__2313 (
            .O(N__15997),
            .I(N__15994));
    LocalMux I__2312 (
            .O(N__15994),
            .I(N__15990));
    InMux I__2311 (
            .O(N__15993),
            .I(N__15987));
    Span4Mux_s3_h I__2310 (
            .O(N__15990),
            .I(N__15984));
    LocalMux I__2309 (
            .O(N__15987),
            .I(\c0.data_in_frame_18_4 ));
    Odrv4 I__2308 (
            .O(N__15984),
            .I(\c0.data_in_frame_18_4 ));
    InMux I__2307 (
            .O(N__15979),
            .I(N__15976));
    LocalMux I__2306 (
            .O(N__15976),
            .I(\c0.n22_adj_1881 ));
    InMux I__2305 (
            .O(N__15973),
            .I(N__15970));
    LocalMux I__2304 (
            .O(N__15970),
            .I(\c0.n5266 ));
    CascadeMux I__2303 (
            .O(N__15967),
            .I(N__15964));
    InMux I__2302 (
            .O(N__15964),
            .I(N__15960));
    InMux I__2301 (
            .O(N__15963),
            .I(N__15955));
    LocalMux I__2300 (
            .O(N__15960),
            .I(N__15952));
    InMux I__2299 (
            .O(N__15959),
            .I(N__15949));
    InMux I__2298 (
            .O(N__15958),
            .I(N__15946));
    LocalMux I__2297 (
            .O(N__15955),
            .I(N__15941));
    Span4Mux_v I__2296 (
            .O(N__15952),
            .I(N__15941));
    LocalMux I__2295 (
            .O(N__15949),
            .I(N__15938));
    LocalMux I__2294 (
            .O(N__15946),
            .I(N__15935));
    Odrv4 I__2293 (
            .O(N__15941),
            .I(\c0.data_in_field_101 ));
    Odrv4 I__2292 (
            .O(N__15938),
            .I(\c0.data_in_field_101 ));
    Odrv4 I__2291 (
            .O(N__15935),
            .I(\c0.data_in_field_101 ));
    CascadeMux I__2290 (
            .O(N__15928),
            .I(\c0.n18_adj_1882_cascade_ ));
    InMux I__2289 (
            .O(N__15925),
            .I(N__15922));
    LocalMux I__2288 (
            .O(N__15922),
            .I(\c0.n26_adj_1883 ));
    CascadeMux I__2287 (
            .O(N__15919),
            .I(\c0.n30_adj_1897_cascade_ ));
    CascadeMux I__2286 (
            .O(N__15916),
            .I(\c0.n36_cascade_ ));
    CascadeMux I__2285 (
            .O(N__15913),
            .I(\c0.n5080_cascade_ ));
    InMux I__2284 (
            .O(N__15910),
            .I(N__15907));
    LocalMux I__2283 (
            .O(N__15907),
            .I(\c0.n1990 ));
    InMux I__2282 (
            .O(N__15904),
            .I(N__15901));
    LocalMux I__2281 (
            .O(N__15901),
            .I(N__15898));
    Odrv4 I__2280 (
            .O(N__15898),
            .I(\c0.n5192 ));
    InMux I__2279 (
            .O(N__15895),
            .I(N__15892));
    LocalMux I__2278 (
            .O(N__15892),
            .I(\c0.n5080 ));
    InMux I__2277 (
            .O(N__15889),
            .I(N__15886));
    LocalMux I__2276 (
            .O(N__15886),
            .I(\c0.n23_adj_1931 ));
    InMux I__2275 (
            .O(N__15883),
            .I(N__15880));
    LocalMux I__2274 (
            .O(N__15880),
            .I(\c0.n21_adj_1928 ));
    CascadeMux I__2273 (
            .O(N__15877),
            .I(\c0.n22_adj_1927_cascade_ ));
    InMux I__2272 (
            .O(N__15874),
            .I(N__15871));
    LocalMux I__2271 (
            .O(N__15871),
            .I(N__15868));
    Odrv4 I__2270 (
            .O(N__15868),
            .I(\c0.n24_adj_1907 ));
    CascadeMux I__2269 (
            .O(N__15865),
            .I(N__15862));
    InMux I__2268 (
            .O(N__15862),
            .I(N__15858));
    InMux I__2267 (
            .O(N__15861),
            .I(N__15854));
    LocalMux I__2266 (
            .O(N__15858),
            .I(N__15850));
    InMux I__2265 (
            .O(N__15857),
            .I(N__15847));
    LocalMux I__2264 (
            .O(N__15854),
            .I(N__15844));
    InMux I__2263 (
            .O(N__15853),
            .I(N__15841));
    Span4Mux_h I__2262 (
            .O(N__15850),
            .I(N__15838));
    LocalMux I__2261 (
            .O(N__15847),
            .I(data_in_19_3));
    Odrv4 I__2260 (
            .O(N__15844),
            .I(data_in_19_3));
    LocalMux I__2259 (
            .O(N__15841),
            .I(data_in_19_3));
    Odrv4 I__2258 (
            .O(N__15838),
            .I(data_in_19_3));
    InMux I__2257 (
            .O(N__15829),
            .I(N__15826));
    LocalMux I__2256 (
            .O(N__15826),
            .I(\c0.n3414 ));
    CascadeMux I__2255 (
            .O(N__15823),
            .I(N__15818));
    InMux I__2254 (
            .O(N__15822),
            .I(N__15813));
    InMux I__2253 (
            .O(N__15821),
            .I(N__15813));
    InMux I__2252 (
            .O(N__15818),
            .I(N__15810));
    LocalMux I__2251 (
            .O(N__15813),
            .I(N__15807));
    LocalMux I__2250 (
            .O(N__15810),
            .I(N__15804));
    Span4Mux_v I__2249 (
            .O(N__15807),
            .I(N__15801));
    Span4Mux_v I__2248 (
            .O(N__15804),
            .I(N__15798));
    Odrv4 I__2247 (
            .O(N__15801),
            .I(\c0.FRAME_MATCHER_wait_for_transmission_N_909 ));
    Odrv4 I__2246 (
            .O(N__15798),
            .I(\c0.FRAME_MATCHER_wait_for_transmission_N_909 ));
    CascadeMux I__2245 (
            .O(N__15793),
            .I(N__15790));
    InMux I__2244 (
            .O(N__15790),
            .I(N__15787));
    LocalMux I__2243 (
            .O(N__15787),
            .I(N__15784));
    Span4Mux_v I__2242 (
            .O(N__15784),
            .I(N__15777));
    InMux I__2241 (
            .O(N__15783),
            .I(N__15772));
    InMux I__2240 (
            .O(N__15782),
            .I(N__15772));
    InMux I__2239 (
            .O(N__15781),
            .I(N__15767));
    InMux I__2238 (
            .O(N__15780),
            .I(N__15767));
    Sp12to4 I__2237 (
            .O(N__15777),
            .I(N__15762));
    LocalMux I__2236 (
            .O(N__15772),
            .I(N__15762));
    LocalMux I__2235 (
            .O(N__15767),
            .I(\c0.r_SM_Main_2_N_1770_0 ));
    Odrv12 I__2234 (
            .O(N__15762),
            .I(\c0.r_SM_Main_2_N_1770_0 ));
    InMux I__2233 (
            .O(N__15757),
            .I(N__15753));
    InMux I__2232 (
            .O(N__15756),
            .I(N__15750));
    LocalMux I__2231 (
            .O(N__15753),
            .I(N__15744));
    LocalMux I__2230 (
            .O(N__15750),
            .I(N__15744));
    InMux I__2229 (
            .O(N__15749),
            .I(N__15741));
    Span4Mux_h I__2228 (
            .O(N__15744),
            .I(N__15738));
    LocalMux I__2227 (
            .O(N__15741),
            .I(tx2_active));
    Odrv4 I__2226 (
            .O(N__15738),
            .I(tx2_active));
    CEMux I__2225 (
            .O(N__15733),
            .I(N__15730));
    LocalMux I__2224 (
            .O(N__15730),
            .I(N__15727));
    Odrv4 I__2223 (
            .O(N__15727),
            .I(\c0.n195 ));
    CascadeMux I__2222 (
            .O(N__15724),
            .I(\c0.n5845_cascade_ ));
    SRMux I__2221 (
            .O(N__15721),
            .I(N__15718));
    LocalMux I__2220 (
            .O(N__15718),
            .I(N__15715));
    Span4Mux_v I__2219 (
            .O(N__15715),
            .I(N__15712));
    Odrv4 I__2218 (
            .O(N__15712),
            .I(\c0.n2275 ));
    InMux I__2217 (
            .O(N__15709),
            .I(N__15706));
    LocalMux I__2216 (
            .O(N__15706),
            .I(N__15703));
    Span4Mux_h I__2215 (
            .O(N__15703),
            .I(N__15697));
    InMux I__2214 (
            .O(N__15702),
            .I(N__15690));
    InMux I__2213 (
            .O(N__15701),
            .I(N__15690));
    InMux I__2212 (
            .O(N__15700),
            .I(N__15690));
    Odrv4 I__2211 (
            .O(N__15697),
            .I(\c0.data_in_field_81 ));
    LocalMux I__2210 (
            .O(N__15690),
            .I(\c0.data_in_field_81 ));
    CascadeMux I__2209 (
            .O(N__15685),
            .I(\c0.n1918_cascade_ ));
    CascadeMux I__2208 (
            .O(N__15682),
            .I(\c0.n5192_cascade_ ));
    CascadeMux I__2207 (
            .O(N__15679),
            .I(\c0.tx.n3507_cascade_ ));
    InMux I__2206 (
            .O(N__15676),
            .I(N__15670));
    InMux I__2205 (
            .O(N__15675),
            .I(N__15670));
    LocalMux I__2204 (
            .O(N__15670),
            .I(n2307));
    InMux I__2203 (
            .O(N__15667),
            .I(N__15655));
    InMux I__2202 (
            .O(N__15666),
            .I(N__15655));
    InMux I__2201 (
            .O(N__15665),
            .I(N__15655));
    InMux I__2200 (
            .O(N__15664),
            .I(N__15655));
    LocalMux I__2199 (
            .O(N__15655),
            .I(n2200));
    CascadeMux I__2198 (
            .O(N__15652),
            .I(n2307_cascade_));
    InMux I__2197 (
            .O(N__15649),
            .I(N__15646));
    LocalMux I__2196 (
            .O(N__15646),
            .I(N__15643));
    Odrv4 I__2195 (
            .O(N__15643),
            .I(n805));
    InMux I__2194 (
            .O(N__15640),
            .I(N__15634));
    InMux I__2193 (
            .O(N__15639),
            .I(N__15634));
    LocalMux I__2192 (
            .O(N__15634),
            .I(N__15628));
    InMux I__2191 (
            .O(N__15633),
            .I(N__15625));
    InMux I__2190 (
            .O(N__15632),
            .I(N__15619));
    InMux I__2189 (
            .O(N__15631),
            .I(N__15619));
    Span4Mux_h I__2188 (
            .O(N__15628),
            .I(N__15614));
    LocalMux I__2187 (
            .O(N__15625),
            .I(N__15614));
    InMux I__2186 (
            .O(N__15624),
            .I(N__15611));
    LocalMux I__2185 (
            .O(N__15619),
            .I(\c0.tx2.r_Bit_Index_0 ));
    Odrv4 I__2184 (
            .O(N__15614),
            .I(\c0.tx2.r_Bit_Index_0 ));
    LocalMux I__2183 (
            .O(N__15611),
            .I(\c0.tx2.r_Bit_Index_0 ));
    CascadeMux I__2182 (
            .O(N__15604),
            .I(N__15599));
    InMux I__2181 (
            .O(N__15603),
            .I(N__15595));
    CascadeMux I__2180 (
            .O(N__15602),
            .I(N__15591));
    InMux I__2179 (
            .O(N__15599),
            .I(N__15587));
    InMux I__2178 (
            .O(N__15598),
            .I(N__15584));
    LocalMux I__2177 (
            .O(N__15595),
            .I(N__15581));
    InMux I__2176 (
            .O(N__15594),
            .I(N__15576));
    InMux I__2175 (
            .O(N__15591),
            .I(N__15576));
    CascadeMux I__2174 (
            .O(N__15590),
            .I(N__15573));
    LocalMux I__2173 (
            .O(N__15587),
            .I(N__15569));
    LocalMux I__2172 (
            .O(N__15584),
            .I(N__15566));
    Span4Mux_s2_h I__2171 (
            .O(N__15581),
            .I(N__15561));
    LocalMux I__2170 (
            .O(N__15576),
            .I(N__15561));
    InMux I__2169 (
            .O(N__15573),
            .I(N__15556));
    InMux I__2168 (
            .O(N__15572),
            .I(N__15556));
    Span4Mux_s3_h I__2167 (
            .O(N__15569),
            .I(N__15553));
    Span4Mux_s3_h I__2166 (
            .O(N__15566),
            .I(N__15550));
    Span4Mux_v I__2165 (
            .O(N__15561),
            .I(N__15547));
    LocalMux I__2164 (
            .O(N__15556),
            .I(\c0.tx2.r_Bit_Index_1 ));
    Odrv4 I__2163 (
            .O(N__15553),
            .I(\c0.tx2.r_Bit_Index_1 ));
    Odrv4 I__2162 (
            .O(N__15550),
            .I(\c0.tx2.r_Bit_Index_1 ));
    Odrv4 I__2161 (
            .O(N__15547),
            .I(\c0.tx2.r_Bit_Index_1 ));
    InMux I__2160 (
            .O(N__15538),
            .I(N__15534));
    InMux I__2159 (
            .O(N__15537),
            .I(N__15531));
    LocalMux I__2158 (
            .O(N__15534),
            .I(N__15527));
    LocalMux I__2157 (
            .O(N__15531),
            .I(N__15524));
    InMux I__2156 (
            .O(N__15530),
            .I(N__15521));
    Span4Mux_s3_h I__2155 (
            .O(N__15527),
            .I(N__15518));
    Span4Mux_v I__2154 (
            .O(N__15524),
            .I(N__15515));
    LocalMux I__2153 (
            .O(N__15521),
            .I(\c0.tx2.r_Bit_Index_2 ));
    Odrv4 I__2152 (
            .O(N__15518),
            .I(\c0.tx2.r_Bit_Index_2 ));
    Odrv4 I__2151 (
            .O(N__15515),
            .I(\c0.tx2.r_Bit_Index_2 ));
    CEMux I__2150 (
            .O(N__15508),
            .I(N__15505));
    LocalMux I__2149 (
            .O(N__15505),
            .I(N__15502));
    Odrv12 I__2148 (
            .O(N__15502),
            .I(\c0.tx2.n2218 ));
    SRMux I__2147 (
            .O(N__15499),
            .I(N__15496));
    LocalMux I__2146 (
            .O(N__15496),
            .I(\c0.tx2.n2319 ));
    CascadeMux I__2145 (
            .O(N__15493),
            .I(N__15490));
    InMux I__2144 (
            .O(N__15490),
            .I(N__15487));
    LocalMux I__2143 (
            .O(N__15487),
            .I(N__15483));
    InMux I__2142 (
            .O(N__15486),
            .I(N__15480));
    Span4Mux_v I__2141 (
            .O(N__15483),
            .I(N__15477));
    LocalMux I__2140 (
            .O(N__15480),
            .I(N__15474));
    Odrv4 I__2139 (
            .O(N__15477),
            .I(n5153));
    Odrv12 I__2138 (
            .O(N__15474),
            .I(n5153));
    CascadeMux I__2137 (
            .O(N__15469),
            .I(\c0.n3414_cascade_ ));
    CascadeMux I__2136 (
            .O(N__15466),
            .I(N__15463));
    InMux I__2135 (
            .O(N__15463),
            .I(N__15460));
    LocalMux I__2134 (
            .O(N__15460),
            .I(N__15457));
    Span4Mux_h I__2133 (
            .O(N__15457),
            .I(N__15454));
    Odrv4 I__2132 (
            .O(N__15454),
            .I(\c0.n9 ));
    InMux I__2131 (
            .O(N__15451),
            .I(N__15448));
    LocalMux I__2130 (
            .O(N__15448),
            .I(N__15445));
    Odrv4 I__2129 (
            .O(N__15445),
            .I(\c0.n5501 ));
    CascadeMux I__2128 (
            .O(N__15442),
            .I(\c0.n1173_cascade_ ));
    CascadeMux I__2127 (
            .O(N__15439),
            .I(tx_data_0_N_keep_cascade_));
    CascadeMux I__2126 (
            .O(N__15436),
            .I(N__15432));
    InMux I__2125 (
            .O(N__15435),
            .I(N__15427));
    InMux I__2124 (
            .O(N__15432),
            .I(N__15427));
    LocalMux I__2123 (
            .O(N__15427),
            .I(r_Tx_Data_0));
    InMux I__2122 (
            .O(N__15424),
            .I(N__15421));
    LocalMux I__2121 (
            .O(N__15421),
            .I(\c0.n5531 ));
    CascadeMux I__2120 (
            .O(N__15418),
            .I(\c0.n15_cascade_ ));
    InMux I__2119 (
            .O(N__15415),
            .I(N__15412));
    LocalMux I__2118 (
            .O(N__15412),
            .I(N__15409));
    Odrv12 I__2117 (
            .O(N__15409),
            .I(tx_data_1_N_keep));
    InMux I__2116 (
            .O(N__15406),
            .I(N__15393));
    InMux I__2115 (
            .O(N__15405),
            .I(N__15393));
    InMux I__2114 (
            .O(N__15404),
            .I(N__15393));
    InMux I__2113 (
            .O(N__15403),
            .I(N__15393));
    InMux I__2112 (
            .O(N__15402),
            .I(N__15390));
    LocalMux I__2111 (
            .O(N__15393),
            .I(\c0.tx.r_SM_Main_2_N_1767_1 ));
    LocalMux I__2110 (
            .O(N__15390),
            .I(\c0.tx.r_SM_Main_2_N_1767_1 ));
    CascadeMux I__2109 (
            .O(N__15385),
            .I(N__15382));
    InMux I__2108 (
            .O(N__15382),
            .I(N__15379));
    LocalMux I__2107 (
            .O(N__15379),
            .I(\c0.tx.n3507 ));
    InMux I__2106 (
            .O(N__15376),
            .I(N__15373));
    LocalMux I__2105 (
            .O(N__15373),
            .I(n5156));
    CascadeMux I__2104 (
            .O(N__15370),
            .I(N__15367));
    InMux I__2103 (
            .O(N__15367),
            .I(N__15364));
    LocalMux I__2102 (
            .O(N__15364),
            .I(N__15361));
    Odrv4 I__2101 (
            .O(N__15361),
            .I(n5063));
    CascadeMux I__2100 (
            .O(N__15358),
            .I(N__15354));
    InMux I__2099 (
            .O(N__15357),
            .I(N__15351));
    InMux I__2098 (
            .O(N__15354),
            .I(N__15348));
    LocalMux I__2097 (
            .O(N__15351),
            .I(data_out_18_3));
    LocalMux I__2096 (
            .O(N__15348),
            .I(data_out_18_3));
    InMux I__2095 (
            .O(N__15343),
            .I(N__15339));
    InMux I__2094 (
            .O(N__15342),
            .I(N__15336));
    LocalMux I__2093 (
            .O(N__15339),
            .I(N__15333));
    LocalMux I__2092 (
            .O(N__15336),
            .I(data_out_19_7));
    Odrv4 I__2091 (
            .O(N__15333),
            .I(data_out_19_7));
    InMux I__2090 (
            .O(N__15328),
            .I(N__15325));
    LocalMux I__2089 (
            .O(N__15325),
            .I(N__15322));
    Odrv12 I__2088 (
            .O(N__15322),
            .I(n7_adj_1998));
    CascadeMux I__2087 (
            .O(N__15319),
            .I(N__15316));
    InMux I__2086 (
            .O(N__15316),
            .I(N__15313));
    LocalMux I__2085 (
            .O(N__15313),
            .I(n8_adj_1997));
    InMux I__2084 (
            .O(N__15310),
            .I(N__15304));
    InMux I__2083 (
            .O(N__15309),
            .I(N__15304));
    LocalMux I__2082 (
            .O(N__15304),
            .I(data_out_18_7));
    CascadeMux I__2081 (
            .O(N__15301),
            .I(N__15298));
    InMux I__2080 (
            .O(N__15298),
            .I(N__15292));
    InMux I__2079 (
            .O(N__15297),
            .I(N__15292));
    LocalMux I__2078 (
            .O(N__15292),
            .I(data_out_19_3));
    InMux I__2077 (
            .O(N__15289),
            .I(N__15285));
    InMux I__2076 (
            .O(N__15288),
            .I(N__15282));
    LocalMux I__2075 (
            .O(N__15285),
            .I(N__15279));
    LocalMux I__2074 (
            .O(N__15282),
            .I(data_out_18_1));
    Odrv4 I__2073 (
            .O(N__15279),
            .I(data_out_18_1));
    CascadeMux I__2072 (
            .O(N__15274),
            .I(N__15271));
    InMux I__2071 (
            .O(N__15271),
            .I(N__15268));
    LocalMux I__2070 (
            .O(N__15268),
            .I(n4_adj_2007));
    InMux I__2069 (
            .O(N__15265),
            .I(N__15261));
    InMux I__2068 (
            .O(N__15264),
            .I(N__15258));
    LocalMux I__2067 (
            .O(N__15261),
            .I(N__15255));
    LocalMux I__2066 (
            .O(N__15258),
            .I(r_Tx_Data_1));
    Odrv4 I__2065 (
            .O(N__15255),
            .I(r_Tx_Data_1));
    CascadeMux I__2064 (
            .O(N__15250),
            .I(N__15246));
    InMux I__2063 (
            .O(N__15249),
            .I(N__15243));
    InMux I__2062 (
            .O(N__15246),
            .I(N__15240));
    LocalMux I__2061 (
            .O(N__15243),
            .I(data_out_19_0));
    LocalMux I__2060 (
            .O(N__15240),
            .I(data_out_19_0));
    CascadeMux I__2059 (
            .O(N__15235),
            .I(N__15232));
    InMux I__2058 (
            .O(N__15232),
            .I(N__15226));
    InMux I__2057 (
            .O(N__15231),
            .I(N__15226));
    LocalMux I__2056 (
            .O(N__15226),
            .I(\c0.delay_counter_9 ));
    InMux I__2055 (
            .O(N__15223),
            .I(N__15219));
    InMux I__2054 (
            .O(N__15222),
            .I(N__15216));
    LocalMux I__2053 (
            .O(N__15219),
            .I(\c0.delay_counter_2 ));
    LocalMux I__2052 (
            .O(N__15216),
            .I(\c0.delay_counter_2 ));
    CascadeMux I__2051 (
            .O(N__15211),
            .I(N__15207));
    CascadeMux I__2050 (
            .O(N__15210),
            .I(N__15204));
    InMux I__2049 (
            .O(N__15207),
            .I(N__15201));
    InMux I__2048 (
            .O(N__15204),
            .I(N__15198));
    LocalMux I__2047 (
            .O(N__15201),
            .I(\c0.delay_counter_0 ));
    LocalMux I__2046 (
            .O(N__15198),
            .I(\c0.delay_counter_0 ));
    InMux I__2045 (
            .O(N__15193),
            .I(N__15189));
    InMux I__2044 (
            .O(N__15192),
            .I(N__15186));
    LocalMux I__2043 (
            .O(N__15189),
            .I(\c0.delay_counter_7 ));
    LocalMux I__2042 (
            .O(N__15186),
            .I(\c0.delay_counter_7 ));
    InMux I__2041 (
            .O(N__15181),
            .I(N__15178));
    LocalMux I__2040 (
            .O(N__15178),
            .I(\c0.n18_adj_1908 ));
    InMux I__2039 (
            .O(N__15175),
            .I(N__15172));
    LocalMux I__2038 (
            .O(N__15172),
            .I(N__15169));
    Odrv4 I__2037 (
            .O(N__15169),
            .I(n4_adj_2000));
    CascadeMux I__2036 (
            .O(N__15166),
            .I(n5086_cascade_));
    InMux I__2035 (
            .O(N__15163),
            .I(N__15159));
    InMux I__2034 (
            .O(N__15162),
            .I(N__15156));
    LocalMux I__2033 (
            .O(N__15159),
            .I(N__15152));
    LocalMux I__2032 (
            .O(N__15156),
            .I(N__15149));
    InMux I__2031 (
            .O(N__15155),
            .I(N__15146));
    Span4Mux_v I__2030 (
            .O(N__15152),
            .I(N__15143));
    Span4Mux_v I__2029 (
            .O(N__15149),
            .I(N__15140));
    LocalMux I__2028 (
            .O(N__15146),
            .I(N__15137));
    Odrv4 I__2027 (
            .O(N__15143),
            .I(n1525));
    Odrv4 I__2026 (
            .O(N__15140),
            .I(n1525));
    Odrv12 I__2025 (
            .O(N__15137),
            .I(n1525));
    CascadeMux I__2024 (
            .O(N__15130),
            .I(n5156_cascade_));
    InMux I__2023 (
            .O(N__15127),
            .I(N__15123));
    InMux I__2022 (
            .O(N__15126),
            .I(N__15120));
    LocalMux I__2021 (
            .O(N__15123),
            .I(data_out_18_0));
    LocalMux I__2020 (
            .O(N__15120),
            .I(data_out_18_0));
    InMux I__2019 (
            .O(N__15115),
            .I(\c0.n4406 ));
    InMux I__2018 (
            .O(N__15112),
            .I(N__15108));
    InMux I__2017 (
            .O(N__15111),
            .I(N__15105));
    LocalMux I__2016 (
            .O(N__15108),
            .I(\c0.delay_counter_4 ));
    LocalMux I__2015 (
            .O(N__15105),
            .I(\c0.delay_counter_4 ));
    InMux I__2014 (
            .O(N__15100),
            .I(\c0.n4407 ));
    InMux I__2013 (
            .O(N__15097),
            .I(N__15093));
    InMux I__2012 (
            .O(N__15096),
            .I(N__15090));
    LocalMux I__2011 (
            .O(N__15093),
            .I(\c0.delay_counter_5 ));
    LocalMux I__2010 (
            .O(N__15090),
            .I(\c0.delay_counter_5 ));
    InMux I__2009 (
            .O(N__15085),
            .I(\c0.n4408 ));
    CascadeMux I__2008 (
            .O(N__15082),
            .I(N__15078));
    InMux I__2007 (
            .O(N__15081),
            .I(N__15075));
    InMux I__2006 (
            .O(N__15078),
            .I(N__15072));
    LocalMux I__2005 (
            .O(N__15075),
            .I(\c0.delay_counter_6 ));
    LocalMux I__2004 (
            .O(N__15072),
            .I(\c0.delay_counter_6 ));
    InMux I__2003 (
            .O(N__15067),
            .I(\c0.n4409 ));
    InMux I__2002 (
            .O(N__15064),
            .I(\c0.n4410 ));
    CascadeMux I__2001 (
            .O(N__15061),
            .I(N__15058));
    InMux I__2000 (
            .O(N__15058),
            .I(N__15054));
    InMux I__1999 (
            .O(N__15057),
            .I(N__15051));
    LocalMux I__1998 (
            .O(N__15054),
            .I(\c0.delay_counter_8 ));
    LocalMux I__1997 (
            .O(N__15051),
            .I(\c0.delay_counter_8 ));
    InMux I__1996 (
            .O(N__15046),
            .I(bfn_4_17_0_));
    InMux I__1995 (
            .O(N__15043),
            .I(\c0.n4412 ));
    InMux I__1994 (
            .O(N__15040),
            .I(\c0.n4413 ));
    InMux I__1993 (
            .O(N__15037),
            .I(N__15033));
    InMux I__1992 (
            .O(N__15036),
            .I(N__15030));
    LocalMux I__1991 (
            .O(N__15033),
            .I(\c0.delay_counter_10 ));
    LocalMux I__1990 (
            .O(N__15030),
            .I(\c0.delay_counter_10 ));
    InMux I__1989 (
            .O(N__15025),
            .I(N__15022));
    LocalMux I__1988 (
            .O(N__15022),
            .I(N__15018));
    InMux I__1987 (
            .O(N__15021),
            .I(N__15015));
    Span4Mux_h I__1986 (
            .O(N__15018),
            .I(N__15012));
    LocalMux I__1985 (
            .O(N__15015),
            .I(N__15009));
    Odrv4 I__1984 (
            .O(N__15012),
            .I(n5077));
    Odrv4 I__1983 (
            .O(N__15009),
            .I(n5077));
    CascadeMux I__1982 (
            .O(N__15004),
            .I(N__15001));
    InMux I__1981 (
            .O(N__15001),
            .I(N__14998));
    LocalMux I__1980 (
            .O(N__14998),
            .I(N__14995));
    Odrv4 I__1979 (
            .O(N__14995),
            .I(n4_adj_1988));
    CEMux I__1978 (
            .O(N__14992),
            .I(N__14989));
    LocalMux I__1977 (
            .O(N__14989),
            .I(N__14985));
    InMux I__1976 (
            .O(N__14988),
            .I(N__14982));
    Odrv12 I__1975 (
            .O(N__14985),
            .I(\c0.rx.n2213 ));
    LocalMux I__1974 (
            .O(N__14982),
            .I(\c0.rx.n2213 ));
    SRMux I__1973 (
            .O(N__14977),
            .I(N__14974));
    LocalMux I__1972 (
            .O(N__14974),
            .I(N__14971));
    Odrv4 I__1971 (
            .O(N__14971),
            .I(\c0.rx.n2317 ));
    InMux I__1970 (
            .O(N__14968),
            .I(N__14951));
    InMux I__1969 (
            .O(N__14967),
            .I(N__14951));
    InMux I__1968 (
            .O(N__14966),
            .I(N__14951));
    InMux I__1967 (
            .O(N__14965),
            .I(N__14951));
    InMux I__1966 (
            .O(N__14964),
            .I(N__14951));
    InMux I__1965 (
            .O(N__14963),
            .I(N__14946));
    InMux I__1964 (
            .O(N__14962),
            .I(N__14946));
    LocalMux I__1963 (
            .O(N__14951),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__1962 (
            .O(N__14946),
            .I(\c0.rx.r_Bit_Index_1 ));
    CascadeMux I__1961 (
            .O(N__14941),
            .I(N__14935));
    InMux I__1960 (
            .O(N__14940),
            .I(N__14924));
    InMux I__1959 (
            .O(N__14939),
            .I(N__14924));
    InMux I__1958 (
            .O(N__14938),
            .I(N__14924));
    InMux I__1957 (
            .O(N__14935),
            .I(N__14924));
    InMux I__1956 (
            .O(N__14934),
            .I(N__14919));
    InMux I__1955 (
            .O(N__14933),
            .I(N__14919));
    LocalMux I__1954 (
            .O(N__14924),
            .I(\c0.rx.r_Bit_Index_2 ));
    LocalMux I__1953 (
            .O(N__14919),
            .I(\c0.rx.r_Bit_Index_2 ));
    InMux I__1952 (
            .O(N__14914),
            .I(N__14908));
    CascadeMux I__1951 (
            .O(N__14913),
            .I(N__14905));
    InMux I__1950 (
            .O(N__14912),
            .I(N__14902));
    InMux I__1949 (
            .O(N__14911),
            .I(N__14899));
    LocalMux I__1948 (
            .O(N__14908),
            .I(N__14896));
    InMux I__1947 (
            .O(N__14905),
            .I(N__14893));
    LocalMux I__1946 (
            .O(N__14902),
            .I(r_Clock_Count_0));
    LocalMux I__1945 (
            .O(N__14899),
            .I(r_Clock_Count_0));
    Odrv4 I__1944 (
            .O(N__14896),
            .I(r_Clock_Count_0));
    LocalMux I__1943 (
            .O(N__14893),
            .I(r_Clock_Count_0));
    CascadeMux I__1942 (
            .O(N__14884),
            .I(N__14878));
    InMux I__1941 (
            .O(N__14883),
            .I(N__14875));
    InMux I__1940 (
            .O(N__14882),
            .I(N__14871));
    InMux I__1939 (
            .O(N__14881),
            .I(N__14868));
    InMux I__1938 (
            .O(N__14878),
            .I(N__14865));
    LocalMux I__1937 (
            .O(N__14875),
            .I(N__14862));
    InMux I__1936 (
            .O(N__14874),
            .I(N__14859));
    LocalMux I__1935 (
            .O(N__14871),
            .I(r_Clock_Count_6));
    LocalMux I__1934 (
            .O(N__14868),
            .I(r_Clock_Count_6));
    LocalMux I__1933 (
            .O(N__14865),
            .I(r_Clock_Count_6));
    Odrv4 I__1932 (
            .O(N__14862),
            .I(r_Clock_Count_6));
    LocalMux I__1931 (
            .O(N__14859),
            .I(r_Clock_Count_6));
    InMux I__1930 (
            .O(N__14848),
            .I(N__14845));
    LocalMux I__1929 (
            .O(N__14845),
            .I(n8_adj_1996));
    IoInMux I__1928 (
            .O(N__14842),
            .I(N__14839));
    LocalMux I__1927 (
            .O(N__14839),
            .I(tx_enable));
    InMux I__1926 (
            .O(N__14836),
            .I(N__14832));
    InMux I__1925 (
            .O(N__14835),
            .I(N__14829));
    LocalMux I__1924 (
            .O(N__14832),
            .I(\c0.delay_counter_1 ));
    LocalMux I__1923 (
            .O(N__14829),
            .I(\c0.delay_counter_1 ));
    InMux I__1922 (
            .O(N__14824),
            .I(\c0.n4404 ));
    InMux I__1921 (
            .O(N__14821),
            .I(\c0.n4405 ));
    InMux I__1920 (
            .O(N__14818),
            .I(N__14814));
    InMux I__1919 (
            .O(N__14817),
            .I(N__14811));
    LocalMux I__1918 (
            .O(N__14814),
            .I(N__14808));
    LocalMux I__1917 (
            .O(N__14811),
            .I(\c0.delay_counter_3 ));
    Odrv4 I__1916 (
            .O(N__14808),
            .I(\c0.delay_counter_3 ));
    InMux I__1915 (
            .O(N__14803),
            .I(N__14800));
    LocalMux I__1914 (
            .O(N__14800),
            .I(\c0.n5671 ));
    InMux I__1913 (
            .O(N__14797),
            .I(N__14794));
    LocalMux I__1912 (
            .O(N__14794),
            .I(N__14790));
    InMux I__1911 (
            .O(N__14793),
            .I(N__14787));
    Odrv4 I__1910 (
            .O(N__14790),
            .I(rx_data_3));
    LocalMux I__1909 (
            .O(N__14787),
            .I(rx_data_3));
    InMux I__1908 (
            .O(N__14782),
            .I(N__14779));
    LocalMux I__1907 (
            .O(N__14779),
            .I(N__14775));
    InMux I__1906 (
            .O(N__14778),
            .I(N__14772));
    Odrv12 I__1905 (
            .O(N__14775),
            .I(rx_data_5));
    LocalMux I__1904 (
            .O(N__14772),
            .I(rx_data_5));
    CascadeMux I__1903 (
            .O(N__14767),
            .I(N__14762));
    InMux I__1902 (
            .O(N__14766),
            .I(N__14757));
    InMux I__1901 (
            .O(N__14765),
            .I(N__14754));
    InMux I__1900 (
            .O(N__14762),
            .I(N__14751));
    InMux I__1899 (
            .O(N__14761),
            .I(N__14746));
    InMux I__1898 (
            .O(N__14760),
            .I(N__14746));
    LocalMux I__1897 (
            .O(N__14757),
            .I(N__14743));
    LocalMux I__1896 (
            .O(N__14754),
            .I(N__14740));
    LocalMux I__1895 (
            .O(N__14751),
            .I(r_Clock_Count_7_adj_2004));
    LocalMux I__1894 (
            .O(N__14746),
            .I(r_Clock_Count_7_adj_2004));
    Odrv4 I__1893 (
            .O(N__14743),
            .I(r_Clock_Count_7_adj_2004));
    Odrv4 I__1892 (
            .O(N__14740),
            .I(r_Clock_Count_7_adj_2004));
    InMux I__1891 (
            .O(N__14731),
            .I(N__14726));
    InMux I__1890 (
            .O(N__14730),
            .I(N__14721));
    InMux I__1889 (
            .O(N__14729),
            .I(N__14718));
    LocalMux I__1888 (
            .O(N__14726),
            .I(N__14715));
    InMux I__1887 (
            .O(N__14725),
            .I(N__14710));
    InMux I__1886 (
            .O(N__14724),
            .I(N__14710));
    LocalMux I__1885 (
            .O(N__14721),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__1884 (
            .O(N__14718),
            .I(\c0.rx.r_Clock_Count_2 ));
    Odrv4 I__1883 (
            .O(N__14715),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__1882 (
            .O(N__14710),
            .I(\c0.rx.r_Clock_Count_2 ));
    InMux I__1881 (
            .O(N__14701),
            .I(N__14698));
    LocalMux I__1880 (
            .O(N__14698),
            .I(N__14695));
    Odrv4 I__1879 (
            .O(N__14695),
            .I(\c0.rx.n6 ));
    InMux I__1878 (
            .O(N__14692),
            .I(N__14686));
    InMux I__1877 (
            .O(N__14691),
            .I(N__14683));
    InMux I__1876 (
            .O(N__14690),
            .I(N__14678));
    InMux I__1875 (
            .O(N__14689),
            .I(N__14678));
    LocalMux I__1874 (
            .O(N__14686),
            .I(\c0.data_in_field_131 ));
    LocalMux I__1873 (
            .O(N__14683),
            .I(\c0.data_in_field_131 ));
    LocalMux I__1872 (
            .O(N__14678),
            .I(\c0.data_in_field_131 ));
    CascadeMux I__1871 (
            .O(N__14671),
            .I(\c0.n2036_cascade_ ));
    CascadeMux I__1870 (
            .O(N__14668),
            .I(\c0.n5273_cascade_ ));
    InMux I__1869 (
            .O(N__14665),
            .I(N__14662));
    LocalMux I__1868 (
            .O(N__14662),
            .I(N__14658));
    InMux I__1867 (
            .O(N__14661),
            .I(N__14655));
    Span4Mux_s3_h I__1866 (
            .O(N__14658),
            .I(N__14652));
    LocalMux I__1865 (
            .O(N__14655),
            .I(\c0.data_in_frame_18_7 ));
    Odrv4 I__1864 (
            .O(N__14652),
            .I(\c0.data_in_frame_18_7 ));
    InMux I__1863 (
            .O(N__14647),
            .I(N__14643));
    CascadeMux I__1862 (
            .O(N__14646),
            .I(N__14640));
    LocalMux I__1861 (
            .O(N__14643),
            .I(N__14636));
    InMux I__1860 (
            .O(N__14640),
            .I(N__14630));
    InMux I__1859 (
            .O(N__14639),
            .I(N__14630));
    Span4Mux_v I__1858 (
            .O(N__14636),
            .I(N__14627));
    InMux I__1857 (
            .O(N__14635),
            .I(N__14624));
    LocalMux I__1856 (
            .O(N__14630),
            .I(data_in_18_3));
    Odrv4 I__1855 (
            .O(N__14627),
            .I(data_in_18_3));
    LocalMux I__1854 (
            .O(N__14624),
            .I(data_in_18_3));
    CascadeMux I__1853 (
            .O(N__14617),
            .I(\c0.n1893_cascade_ ));
    InMux I__1852 (
            .O(N__14614),
            .I(N__14611));
    LocalMux I__1851 (
            .O(N__14611),
            .I(\c0.n20_adj_1921 ));
    InMux I__1850 (
            .O(N__14608),
            .I(N__14605));
    LocalMux I__1849 (
            .O(N__14605),
            .I(\c0.n5459 ));
    InMux I__1848 (
            .O(N__14602),
            .I(N__14599));
    LocalMux I__1847 (
            .O(N__14599),
            .I(N__14596));
    Odrv4 I__1846 (
            .O(N__14596),
            .I(\c0.n5737 ));
    CascadeMux I__1845 (
            .O(N__14593),
            .I(N__14590));
    InMux I__1844 (
            .O(N__14590),
            .I(N__14587));
    LocalMux I__1843 (
            .O(N__14587),
            .I(N__14583));
    InMux I__1842 (
            .O(N__14586),
            .I(N__14580));
    Span12Mux_s2_h I__1841 (
            .O(N__14583),
            .I(N__14577));
    LocalMux I__1840 (
            .O(N__14580),
            .I(\c0.data_in_frame_19_1 ));
    Odrv12 I__1839 (
            .O(N__14577),
            .I(\c0.data_in_frame_19_1 ));
    CascadeMux I__1838 (
            .O(N__14572),
            .I(N__14569));
    InMux I__1837 (
            .O(N__14569),
            .I(N__14566));
    LocalMux I__1836 (
            .O(N__14566),
            .I(N__14563));
    Odrv4 I__1835 (
            .O(N__14563),
            .I(\c0.n5944 ));
    CascadeMux I__1834 (
            .O(N__14560),
            .I(N__14556));
    CascadeMux I__1833 (
            .O(N__14559),
            .I(N__14553));
    InMux I__1832 (
            .O(N__14556),
            .I(N__14550));
    InMux I__1831 (
            .O(N__14553),
            .I(N__14547));
    LocalMux I__1830 (
            .O(N__14550),
            .I(\c0.data_in_frame_19_6 ));
    LocalMux I__1829 (
            .O(N__14547),
            .I(\c0.data_in_frame_19_6 ));
    InMux I__1828 (
            .O(N__14542),
            .I(N__14539));
    LocalMux I__1827 (
            .O(N__14539),
            .I(\c0.n5456 ));
    InMux I__1826 (
            .O(N__14536),
            .I(\c0.n4403 ));
    CascadeMux I__1825 (
            .O(N__14533),
            .I(N__14527));
    InMux I__1824 (
            .O(N__14532),
            .I(N__14518));
    InMux I__1823 (
            .O(N__14531),
            .I(N__14518));
    InMux I__1822 (
            .O(N__14530),
            .I(N__14518));
    InMux I__1821 (
            .O(N__14527),
            .I(N__14515));
    InMux I__1820 (
            .O(N__14526),
            .I(N__14512));
    InMux I__1819 (
            .O(N__14525),
            .I(N__14506));
    LocalMux I__1818 (
            .O(N__14518),
            .I(N__14500));
    LocalMux I__1817 (
            .O(N__14515),
            .I(N__14500));
    LocalMux I__1816 (
            .O(N__14512),
            .I(N__14497));
    InMux I__1815 (
            .O(N__14511),
            .I(N__14490));
    InMux I__1814 (
            .O(N__14510),
            .I(N__14490));
    InMux I__1813 (
            .O(N__14509),
            .I(N__14490));
    LocalMux I__1812 (
            .O(N__14506),
            .I(N__14487));
    InMux I__1811 (
            .O(N__14505),
            .I(N__14484));
    Span4Mux_s3_h I__1810 (
            .O(N__14500),
            .I(N__14481));
    Odrv4 I__1809 (
            .O(N__14497),
            .I(\c0.byte_transmit_counter2_4 ));
    LocalMux I__1808 (
            .O(N__14490),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__1807 (
            .O(N__14487),
            .I(\c0.byte_transmit_counter2_4 ));
    LocalMux I__1806 (
            .O(N__14484),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__1805 (
            .O(N__14481),
            .I(\c0.byte_transmit_counter2_4 ));
    CascadeMux I__1804 (
            .O(N__14470),
            .I(\c0.n5785_cascade_ ));
    InMux I__1803 (
            .O(N__14467),
            .I(N__14464));
    LocalMux I__1802 (
            .O(N__14464),
            .I(N__14461));
    Odrv4 I__1801 (
            .O(N__14461),
            .I(\c0.n5426 ));
    InMux I__1800 (
            .O(N__14458),
            .I(N__14455));
    LocalMux I__1799 (
            .O(N__14455),
            .I(\c0.n5788 ));
    CascadeMux I__1798 (
            .O(N__14452),
            .I(N__14449));
    InMux I__1797 (
            .O(N__14449),
            .I(N__14446));
    LocalMux I__1796 (
            .O(N__14446),
            .I(\c0.n5968 ));
    CascadeMux I__1795 (
            .O(N__14443),
            .I(N__14440));
    InMux I__1794 (
            .O(N__14440),
            .I(N__14437));
    LocalMux I__1793 (
            .O(N__14437),
            .I(N__14434));
    Odrv12 I__1792 (
            .O(N__14434),
            .I(\c0.n5363 ));
    CascadeMux I__1791 (
            .O(N__14431),
            .I(N__14428));
    InMux I__1790 (
            .O(N__14428),
            .I(N__14424));
    InMux I__1789 (
            .O(N__14427),
            .I(N__14421));
    LocalMux I__1788 (
            .O(N__14424),
            .I(N__14418));
    LocalMux I__1787 (
            .O(N__14421),
            .I(N__14415));
    Span4Mux_s2_h I__1786 (
            .O(N__14418),
            .I(N__14412));
    Odrv4 I__1785 (
            .O(N__14415),
            .I(\c0.data_in_frame_19_7 ));
    Odrv4 I__1784 (
            .O(N__14412),
            .I(\c0.data_in_frame_19_7 ));
    CascadeMux I__1783 (
            .O(N__14407),
            .I(N__14404));
    InMux I__1782 (
            .O(N__14404),
            .I(N__14401));
    LocalMux I__1781 (
            .O(N__14401),
            .I(\c0.n5935 ));
    InMux I__1780 (
            .O(N__14398),
            .I(N__14394));
    CascadeMux I__1779 (
            .O(N__14397),
            .I(N__14382));
    LocalMux I__1778 (
            .O(N__14394),
            .I(N__14379));
    InMux I__1777 (
            .O(N__14393),
            .I(N__14372));
    InMux I__1776 (
            .O(N__14392),
            .I(N__14372));
    InMux I__1775 (
            .O(N__14391),
            .I(N__14372));
    CascadeMux I__1774 (
            .O(N__14390),
            .I(N__14369));
    CascadeMux I__1773 (
            .O(N__14389),
            .I(N__14365));
    InMux I__1772 (
            .O(N__14388),
            .I(N__14362));
    InMux I__1771 (
            .O(N__14387),
            .I(N__14353));
    InMux I__1770 (
            .O(N__14386),
            .I(N__14353));
    InMux I__1769 (
            .O(N__14385),
            .I(N__14353));
    InMux I__1768 (
            .O(N__14382),
            .I(N__14353));
    Span4Mux_v I__1767 (
            .O(N__14379),
            .I(N__14350));
    LocalMux I__1766 (
            .O(N__14372),
            .I(N__14347));
    InMux I__1765 (
            .O(N__14369),
            .I(N__14344));
    InMux I__1764 (
            .O(N__14368),
            .I(N__14339));
    InMux I__1763 (
            .O(N__14365),
            .I(N__14339));
    LocalMux I__1762 (
            .O(N__14362),
            .I(r_SM_Main_1_adj_2010));
    LocalMux I__1761 (
            .O(N__14353),
            .I(r_SM_Main_1_adj_2010));
    Odrv4 I__1760 (
            .O(N__14350),
            .I(r_SM_Main_1_adj_2010));
    Odrv12 I__1759 (
            .O(N__14347),
            .I(r_SM_Main_1_adj_2010));
    LocalMux I__1758 (
            .O(N__14344),
            .I(r_SM_Main_1_adj_2010));
    LocalMux I__1757 (
            .O(N__14339),
            .I(r_SM_Main_1_adj_2010));
    CascadeMux I__1756 (
            .O(N__14326),
            .I(\c0.tx2.n2218_cascade_ ));
    InMux I__1755 (
            .O(N__14323),
            .I(N__14319));
    CascadeMux I__1754 (
            .O(N__14322),
            .I(N__14315));
    LocalMux I__1753 (
            .O(N__14319),
            .I(N__14312));
    InMux I__1752 (
            .O(N__14318),
            .I(N__14309));
    InMux I__1751 (
            .O(N__14315),
            .I(N__14306));
    Span4Mux_v I__1750 (
            .O(N__14312),
            .I(N__14303));
    LocalMux I__1749 (
            .O(N__14309),
            .I(\c0.tx2.n3577 ));
    LocalMux I__1748 (
            .O(N__14306),
            .I(\c0.tx2.n3577 ));
    Odrv4 I__1747 (
            .O(N__14303),
            .I(\c0.tx2.n3577 ));
    CascadeMux I__1746 (
            .O(N__14296),
            .I(N__14293));
    InMux I__1745 (
            .O(N__14293),
            .I(N__14290));
    LocalMux I__1744 (
            .O(N__14290),
            .I(N__14287));
    Odrv4 I__1743 (
            .O(N__14287),
            .I(\c0.n5953 ));
    CascadeMux I__1742 (
            .O(N__14284),
            .I(N__14281));
    InMux I__1741 (
            .O(N__14281),
            .I(N__14278));
    LocalMux I__1740 (
            .O(N__14278),
            .I(N__14275));
    Span4Mux_s2_h I__1739 (
            .O(N__14275),
            .I(N__14272));
    Odrv4 I__1738 (
            .O(N__14272),
            .I(\c0.n5956 ));
    InMux I__1737 (
            .O(N__14269),
            .I(N__14266));
    LocalMux I__1736 (
            .O(N__14266),
            .I(n2392));
    CascadeMux I__1735 (
            .O(N__14263),
            .I(N__14245));
    CascadeMux I__1734 (
            .O(N__14262),
            .I(N__14242));
    CascadeMux I__1733 (
            .O(N__14261),
            .I(N__14229));
    CascadeMux I__1732 (
            .O(N__14260),
            .I(N__14226));
    CascadeMux I__1731 (
            .O(N__14259),
            .I(N__14223));
    CascadeMux I__1730 (
            .O(N__14258),
            .I(N__14220));
    CascadeMux I__1729 (
            .O(N__14257),
            .I(N__14217));
    CascadeMux I__1728 (
            .O(N__14256),
            .I(N__14214));
    CascadeMux I__1727 (
            .O(N__14255),
            .I(N__14211));
    CascadeMux I__1726 (
            .O(N__14254),
            .I(N__14208));
    InMux I__1725 (
            .O(N__14253),
            .I(N__14204));
    CascadeMux I__1724 (
            .O(N__14252),
            .I(N__14201));
    CascadeMux I__1723 (
            .O(N__14251),
            .I(N__14198));
    CascadeMux I__1722 (
            .O(N__14250),
            .I(N__14195));
    CascadeMux I__1721 (
            .O(N__14249),
            .I(N__14192));
    InMux I__1720 (
            .O(N__14248),
            .I(N__14181));
    InMux I__1719 (
            .O(N__14245),
            .I(N__14181));
    InMux I__1718 (
            .O(N__14242),
            .I(N__14181));
    InMux I__1717 (
            .O(N__14241),
            .I(N__14181));
    InMux I__1716 (
            .O(N__14240),
            .I(N__14181));
    InMux I__1715 (
            .O(N__14239),
            .I(N__14174));
    InMux I__1714 (
            .O(N__14238),
            .I(N__14174));
    InMux I__1713 (
            .O(N__14237),
            .I(N__14174));
    InMux I__1712 (
            .O(N__14236),
            .I(N__14169));
    InMux I__1711 (
            .O(N__14235),
            .I(N__14169));
    InMux I__1710 (
            .O(N__14234),
            .I(N__14162));
    InMux I__1709 (
            .O(N__14233),
            .I(N__14162));
    InMux I__1708 (
            .O(N__14232),
            .I(N__14162));
    InMux I__1707 (
            .O(N__14229),
            .I(N__14153));
    InMux I__1706 (
            .O(N__14226),
            .I(N__14153));
    InMux I__1705 (
            .O(N__14223),
            .I(N__14153));
    InMux I__1704 (
            .O(N__14220),
            .I(N__14153));
    InMux I__1703 (
            .O(N__14217),
            .I(N__14144));
    InMux I__1702 (
            .O(N__14214),
            .I(N__14144));
    InMux I__1701 (
            .O(N__14211),
            .I(N__14144));
    InMux I__1700 (
            .O(N__14208),
            .I(N__14144));
    InMux I__1699 (
            .O(N__14207),
            .I(N__14141));
    LocalMux I__1698 (
            .O(N__14204),
            .I(N__14138));
    InMux I__1697 (
            .O(N__14201),
            .I(N__14135));
    InMux I__1696 (
            .O(N__14198),
            .I(N__14128));
    InMux I__1695 (
            .O(N__14195),
            .I(N__14128));
    InMux I__1694 (
            .O(N__14192),
            .I(N__14128));
    LocalMux I__1693 (
            .O(N__14181),
            .I(N__14121));
    LocalMux I__1692 (
            .O(N__14174),
            .I(N__14121));
    LocalMux I__1691 (
            .O(N__14169),
            .I(N__14121));
    LocalMux I__1690 (
            .O(N__14162),
            .I(N__14114));
    LocalMux I__1689 (
            .O(N__14153),
            .I(N__14114));
    LocalMux I__1688 (
            .O(N__14144),
            .I(N__14114));
    LocalMux I__1687 (
            .O(N__14141),
            .I(r_SM_Main_2_adj_2009));
    Odrv4 I__1686 (
            .O(N__14138),
            .I(r_SM_Main_2_adj_2009));
    LocalMux I__1685 (
            .O(N__14135),
            .I(r_SM_Main_2_adj_2009));
    LocalMux I__1684 (
            .O(N__14128),
            .I(r_SM_Main_2_adj_2009));
    Odrv4 I__1683 (
            .O(N__14121),
            .I(r_SM_Main_2_adj_2009));
    Odrv4 I__1682 (
            .O(N__14114),
            .I(r_SM_Main_2_adj_2009));
    InMux I__1681 (
            .O(N__14101),
            .I(N__14098));
    LocalMux I__1680 (
            .O(N__14098),
            .I(N__14093));
    InMux I__1679 (
            .O(N__14097),
            .I(N__14088));
    InMux I__1678 (
            .O(N__14096),
            .I(N__14088));
    Span4Mux_v I__1677 (
            .O(N__14093),
            .I(N__14080));
    LocalMux I__1676 (
            .O(N__14088),
            .I(N__14077));
    InMux I__1675 (
            .O(N__14087),
            .I(N__14068));
    InMux I__1674 (
            .O(N__14086),
            .I(N__14068));
    InMux I__1673 (
            .O(N__14085),
            .I(N__14068));
    InMux I__1672 (
            .O(N__14084),
            .I(N__14068));
    InMux I__1671 (
            .O(N__14083),
            .I(N__14065));
    Odrv4 I__1670 (
            .O(N__14080),
            .I(n5037));
    Odrv4 I__1669 (
            .O(N__14077),
            .I(n5037));
    LocalMux I__1668 (
            .O(N__14068),
            .I(n5037));
    LocalMux I__1667 (
            .O(N__14065),
            .I(n5037));
    InMux I__1666 (
            .O(N__14056),
            .I(N__14051));
    InMux I__1665 (
            .O(N__14055),
            .I(N__14048));
    InMux I__1664 (
            .O(N__14054),
            .I(N__14045));
    LocalMux I__1663 (
            .O(N__14051),
            .I(\c0.tx2.r_Clock_Count_3 ));
    LocalMux I__1662 (
            .O(N__14048),
            .I(\c0.tx2.r_Clock_Count_3 ));
    LocalMux I__1661 (
            .O(N__14045),
            .I(\c0.tx2.r_Clock_Count_3 ));
    InMux I__1660 (
            .O(N__14038),
            .I(\c0.n4400 ));
    InMux I__1659 (
            .O(N__14035),
            .I(\c0.n4401 ));
    InMux I__1658 (
            .O(N__14032),
            .I(\c0.n4402 ));
    CascadeMux I__1657 (
            .O(N__14029),
            .I(\c0.tx.n12_cascade_ ));
    InMux I__1656 (
            .O(N__14026),
            .I(N__14019));
    InMux I__1655 (
            .O(N__14025),
            .I(N__14014));
    InMux I__1654 (
            .O(N__14024),
            .I(N__14014));
    InMux I__1653 (
            .O(N__14023),
            .I(N__14011));
    InMux I__1652 (
            .O(N__14022),
            .I(N__14008));
    LocalMux I__1651 (
            .O(N__14019),
            .I(r_Clock_Count_8));
    LocalMux I__1650 (
            .O(N__14014),
            .I(r_Clock_Count_8));
    LocalMux I__1649 (
            .O(N__14011),
            .I(r_Clock_Count_8));
    LocalMux I__1648 (
            .O(N__14008),
            .I(r_Clock_Count_8));
    CascadeMux I__1647 (
            .O(N__13999),
            .I(n1307_cascade_));
    InMux I__1646 (
            .O(N__13996),
            .I(N__13992));
    InMux I__1645 (
            .O(N__13995),
            .I(N__13989));
    LocalMux I__1644 (
            .O(N__13992),
            .I(n3595));
    LocalMux I__1643 (
            .O(N__13989),
            .I(n3595));
    InMux I__1642 (
            .O(N__13984),
            .I(N__13973));
    InMux I__1641 (
            .O(N__13983),
            .I(N__13968));
    InMux I__1640 (
            .O(N__13982),
            .I(N__13968));
    InMux I__1639 (
            .O(N__13981),
            .I(N__13963));
    InMux I__1638 (
            .O(N__13980),
            .I(N__13963));
    InMux I__1637 (
            .O(N__13979),
            .I(N__13954));
    InMux I__1636 (
            .O(N__13978),
            .I(N__13954));
    InMux I__1635 (
            .O(N__13977),
            .I(N__13954));
    InMux I__1634 (
            .O(N__13976),
            .I(N__13954));
    LocalMux I__1633 (
            .O(N__13973),
            .I(N__13951));
    LocalMux I__1632 (
            .O(N__13968),
            .I(n4221));
    LocalMux I__1631 (
            .O(N__13963),
            .I(n4221));
    LocalMux I__1630 (
            .O(N__13954),
            .I(n4221));
    Odrv4 I__1629 (
            .O(N__13951),
            .I(n4221));
    InMux I__1628 (
            .O(N__13942),
            .I(N__13939));
    LocalMux I__1627 (
            .O(N__13939),
            .I(n2));
    InMux I__1626 (
            .O(N__13936),
            .I(N__13933));
    LocalMux I__1625 (
            .O(N__13933),
            .I(n1307));
    CascadeMux I__1624 (
            .O(N__13930),
            .I(n4_adj_2003_cascade_));
    CascadeMux I__1623 (
            .O(N__13927),
            .I(N__13923));
    InMux I__1622 (
            .O(N__13926),
            .I(N__13920));
    InMux I__1621 (
            .O(N__13923),
            .I(N__13917));
    LocalMux I__1620 (
            .O(N__13920),
            .I(n4155));
    LocalMux I__1619 (
            .O(N__13917),
            .I(n4155));
    CascadeMux I__1618 (
            .O(N__13912),
            .I(N__13909));
    InMux I__1617 (
            .O(N__13909),
            .I(N__13906));
    LocalMux I__1616 (
            .O(N__13906),
            .I(n2372));
    InMux I__1615 (
            .O(N__13903),
            .I(N__13898));
    InMux I__1614 (
            .O(N__13902),
            .I(N__13895));
    InMux I__1613 (
            .O(N__13901),
            .I(N__13892));
    LocalMux I__1612 (
            .O(N__13898),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__1611 (
            .O(N__13895),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__1610 (
            .O(N__13892),
            .I(\c0.tx2.r_Clock_Count_7 ));
    InMux I__1609 (
            .O(N__13885),
            .I(N__13882));
    LocalMux I__1608 (
            .O(N__13882),
            .I(n2395));
    InMux I__1607 (
            .O(N__13879),
            .I(N__13874));
    InMux I__1606 (
            .O(N__13878),
            .I(N__13871));
    InMux I__1605 (
            .O(N__13877),
            .I(N__13868));
    LocalMux I__1604 (
            .O(N__13874),
            .I(\c0.tx2.r_Clock_Count_2 ));
    LocalMux I__1603 (
            .O(N__13871),
            .I(\c0.tx2.r_Clock_Count_2 ));
    LocalMux I__1602 (
            .O(N__13868),
            .I(\c0.tx2.r_Clock_Count_2 ));
    InMux I__1601 (
            .O(N__13861),
            .I(N__13857));
    InMux I__1600 (
            .O(N__13860),
            .I(N__13847));
    LocalMux I__1599 (
            .O(N__13857),
            .I(N__13844));
    InMux I__1598 (
            .O(N__13856),
            .I(N__13841));
    InMux I__1597 (
            .O(N__13855),
            .I(N__13838));
    InMux I__1596 (
            .O(N__13854),
            .I(N__13831));
    InMux I__1595 (
            .O(N__13853),
            .I(N__13831));
    InMux I__1594 (
            .O(N__13852),
            .I(N__13831));
    InMux I__1593 (
            .O(N__13851),
            .I(N__13826));
    InMux I__1592 (
            .O(N__13850),
            .I(N__13826));
    LocalMux I__1591 (
            .O(N__13847),
            .I(N__13819));
    Span4Mux_v I__1590 (
            .O(N__13844),
            .I(N__13819));
    LocalMux I__1589 (
            .O(N__13841),
            .I(N__13819));
    LocalMux I__1588 (
            .O(N__13838),
            .I(N__13816));
    LocalMux I__1587 (
            .O(N__13831),
            .I(r_SM_Main_0_adj_2011));
    LocalMux I__1586 (
            .O(N__13826),
            .I(r_SM_Main_0_adj_2011));
    Odrv4 I__1585 (
            .O(N__13819),
            .I(r_SM_Main_0_adj_2011));
    Odrv4 I__1584 (
            .O(N__13816),
            .I(r_SM_Main_0_adj_2011));
    InMux I__1583 (
            .O(N__13807),
            .I(N__13796));
    InMux I__1582 (
            .O(N__13806),
            .I(N__13796));
    InMux I__1581 (
            .O(N__13805),
            .I(N__13796));
    InMux I__1580 (
            .O(N__13804),
            .I(N__13790));
    InMux I__1579 (
            .O(N__13803),
            .I(N__13790));
    LocalMux I__1578 (
            .O(N__13796),
            .I(N__13787));
    InMux I__1577 (
            .O(N__13795),
            .I(N__13784));
    LocalMux I__1576 (
            .O(N__13790),
            .I(r_SM_Main_2_N_1767_1));
    Odrv4 I__1575 (
            .O(N__13787),
            .I(r_SM_Main_2_N_1767_1));
    LocalMux I__1574 (
            .O(N__13784),
            .I(r_SM_Main_2_N_1767_1));
    InMux I__1573 (
            .O(N__13777),
            .I(N__13773));
    InMux I__1572 (
            .O(N__13776),
            .I(N__13770));
    LocalMux I__1571 (
            .O(N__13773),
            .I(N__13765));
    LocalMux I__1570 (
            .O(N__13770),
            .I(N__13765));
    Odrv4 I__1569 (
            .O(N__13765),
            .I(data_out_19_4));
    InMux I__1568 (
            .O(N__13762),
            .I(N__13756));
    InMux I__1567 (
            .O(N__13761),
            .I(N__13756));
    LocalMux I__1566 (
            .O(N__13756),
            .I(data_out_18_4));
    CascadeMux I__1565 (
            .O(N__13753),
            .I(\c0.n17_cascade_ ));
    CascadeMux I__1564 (
            .O(N__13750),
            .I(tx_data_4_N_keep_cascade_));
    InMux I__1563 (
            .O(N__13747),
            .I(N__13744));
    LocalMux I__1562 (
            .O(N__13744),
            .I(N__13741));
    Odrv4 I__1561 (
            .O(N__13741),
            .I(n8_adj_2001));
    CascadeMux I__1560 (
            .O(N__13738),
            .I(\c0.tx.r_SM_Main_2_N_1767_1_cascade_ ));
    InMux I__1559 (
            .O(N__13735),
            .I(N__13732));
    LocalMux I__1558 (
            .O(N__13732),
            .I(n5041));
    InMux I__1557 (
            .O(N__13729),
            .I(N__13726));
    LocalMux I__1556 (
            .O(N__13726),
            .I(N__13720));
    InMux I__1555 (
            .O(N__13725),
            .I(N__13717));
    InMux I__1554 (
            .O(N__13724),
            .I(N__13714));
    CascadeMux I__1553 (
            .O(N__13723),
            .I(N__13711));
    Span4Mux_v I__1552 (
            .O(N__13720),
            .I(N__13703));
    LocalMux I__1551 (
            .O(N__13717),
            .I(N__13703));
    LocalMux I__1550 (
            .O(N__13714),
            .I(N__13703));
    InMux I__1549 (
            .O(N__13711),
            .I(N__13697));
    InMux I__1548 (
            .O(N__13710),
            .I(N__13697));
    Span4Mux_v I__1547 (
            .O(N__13703),
            .I(N__13694));
    InMux I__1546 (
            .O(N__13702),
            .I(N__13691));
    LocalMux I__1545 (
            .O(N__13697),
            .I(\c0.tx_transmit ));
    Odrv4 I__1544 (
            .O(N__13694),
            .I(\c0.tx_transmit ));
    LocalMux I__1543 (
            .O(N__13691),
            .I(\c0.tx_transmit ));
    CascadeMux I__1542 (
            .O(N__13684),
            .I(n4316_cascade_));
    CascadeMux I__1541 (
            .O(N__13681),
            .I(N__13678));
    InMux I__1540 (
            .O(N__13678),
            .I(N__13675));
    LocalMux I__1539 (
            .O(N__13675),
            .I(n7_adj_2002));
    InMux I__1538 (
            .O(N__13672),
            .I(N__13668));
    InMux I__1537 (
            .O(N__13671),
            .I(N__13665));
    LocalMux I__1536 (
            .O(N__13668),
            .I(N__13662));
    LocalMux I__1535 (
            .O(N__13665),
            .I(n5066));
    Odrv4 I__1534 (
            .O(N__13662),
            .I(n5066));
    CascadeMux I__1533 (
            .O(N__13657),
            .I(N__13651));
    InMux I__1532 (
            .O(N__13656),
            .I(N__13646));
    InMux I__1531 (
            .O(N__13655),
            .I(N__13646));
    InMux I__1530 (
            .O(N__13654),
            .I(N__13643));
    InMux I__1529 (
            .O(N__13651),
            .I(N__13638));
    LocalMux I__1528 (
            .O(N__13646),
            .I(N__13635));
    LocalMux I__1527 (
            .O(N__13643),
            .I(N__13632));
    InMux I__1526 (
            .O(N__13642),
            .I(N__13627));
    InMux I__1525 (
            .O(N__13641),
            .I(N__13627));
    LocalMux I__1524 (
            .O(N__13638),
            .I(tx_active));
    Odrv4 I__1523 (
            .O(N__13635),
            .I(tx_active));
    Odrv4 I__1522 (
            .O(N__13632),
            .I(tx_active));
    LocalMux I__1521 (
            .O(N__13627),
            .I(tx_active));
    InMux I__1520 (
            .O(N__13618),
            .I(N__13614));
    InMux I__1519 (
            .O(N__13617),
            .I(N__13611));
    LocalMux I__1518 (
            .O(N__13614),
            .I(\c0.tx_transmit_N_568_5 ));
    LocalMux I__1517 (
            .O(N__13611),
            .I(\c0.tx_transmit_N_568_5 ));
    InMux I__1516 (
            .O(N__13606),
            .I(N__13602));
    InMux I__1515 (
            .O(N__13605),
            .I(N__13599));
    LocalMux I__1514 (
            .O(N__13602),
            .I(\c0.tx_transmit_N_568_6 ));
    LocalMux I__1513 (
            .O(N__13599),
            .I(\c0.tx_transmit_N_568_6 ));
    InMux I__1512 (
            .O(N__13594),
            .I(N__13590));
    InMux I__1511 (
            .O(N__13593),
            .I(N__13587));
    LocalMux I__1510 (
            .O(N__13590),
            .I(\c0.tx_transmit_N_568_7 ));
    LocalMux I__1509 (
            .O(N__13587),
            .I(\c0.tx_transmit_N_568_7 ));
    InMux I__1508 (
            .O(N__13582),
            .I(N__13576));
    InMux I__1507 (
            .O(N__13581),
            .I(N__13571));
    InMux I__1506 (
            .O(N__13580),
            .I(N__13571));
    InMux I__1505 (
            .O(N__13579),
            .I(N__13568));
    LocalMux I__1504 (
            .O(N__13576),
            .I(\c0.tx_transmit_N_568_4 ));
    LocalMux I__1503 (
            .O(N__13571),
            .I(\c0.tx_transmit_N_568_4 ));
    LocalMux I__1502 (
            .O(N__13568),
            .I(\c0.tx_transmit_N_568_4 ));
    InMux I__1501 (
            .O(N__13561),
            .I(N__13557));
    InMux I__1500 (
            .O(N__13560),
            .I(N__13554));
    LocalMux I__1499 (
            .O(N__13557),
            .I(\c0.n103 ));
    LocalMux I__1498 (
            .O(N__13554),
            .I(\c0.n103 ));
    InMux I__1497 (
            .O(N__13549),
            .I(N__13546));
    LocalMux I__1496 (
            .O(N__13546),
            .I(\c0.n109 ));
    InMux I__1495 (
            .O(N__13543),
            .I(N__13534));
    InMux I__1494 (
            .O(N__13542),
            .I(N__13534));
    InMux I__1493 (
            .O(N__13541),
            .I(N__13529));
    InMux I__1492 (
            .O(N__13540),
            .I(N__13529));
    InMux I__1491 (
            .O(N__13539),
            .I(N__13526));
    LocalMux I__1490 (
            .O(N__13534),
            .I(\c0.n45 ));
    LocalMux I__1489 (
            .O(N__13529),
            .I(\c0.n45 ));
    LocalMux I__1488 (
            .O(N__13526),
            .I(\c0.n45 ));
    CascadeMux I__1487 (
            .O(N__13519),
            .I(\c0.n109_cascade_ ));
    CascadeMux I__1486 (
            .O(N__13516),
            .I(n4315_cascade_));
    InMux I__1485 (
            .O(N__13513),
            .I(N__13510));
    LocalMux I__1484 (
            .O(N__13510),
            .I(N__13506));
    CascadeMux I__1483 (
            .O(N__13509),
            .I(N__13503));
    Span4Mux_v I__1482 (
            .O(N__13506),
            .I(N__13500));
    InMux I__1481 (
            .O(N__13503),
            .I(N__13497));
    Odrv4 I__1480 (
            .O(N__13500),
            .I(\c0.rx.n3573 ));
    LocalMux I__1479 (
            .O(N__13497),
            .I(\c0.rx.n3573 ));
    CascadeMux I__1478 (
            .O(N__13492),
            .I(\c0.rx.n3573_cascade_ ));
    CascadeMux I__1477 (
            .O(N__13489),
            .I(\c0.n20_adj_1918_cascade_ ));
    CascadeMux I__1476 (
            .O(N__13486),
            .I(N__13482));
    CascadeMux I__1475 (
            .O(N__13485),
            .I(N__13479));
    InMux I__1474 (
            .O(N__13482),
            .I(N__13465));
    InMux I__1473 (
            .O(N__13479),
            .I(N__13465));
    InMux I__1472 (
            .O(N__13478),
            .I(N__13465));
    InMux I__1471 (
            .O(N__13477),
            .I(N__13465));
    InMux I__1470 (
            .O(N__13476),
            .I(N__13465));
    LocalMux I__1469 (
            .O(N__13465),
            .I(\c0.n87 ));
    CascadeMux I__1468 (
            .O(N__13462),
            .I(\c0.n87_cascade_ ));
    InMux I__1467 (
            .O(N__13459),
            .I(N__13456));
    LocalMux I__1466 (
            .O(N__13456),
            .I(\c0.n16_adj_1909 ));
    CascadeMux I__1465 (
            .O(N__13453),
            .I(\c0.rx.n4_adj_1866_cascade_ ));
    InMux I__1464 (
            .O(N__13450),
            .I(N__13441));
    InMux I__1463 (
            .O(N__13449),
            .I(N__13441));
    InMux I__1462 (
            .O(N__13448),
            .I(N__13441));
    LocalMux I__1461 (
            .O(N__13441),
            .I(N__13436));
    InMux I__1460 (
            .O(N__13440),
            .I(N__13431));
    InMux I__1459 (
            .O(N__13439),
            .I(N__13431));
    Span4Mux_s1_h I__1458 (
            .O(N__13436),
            .I(N__13428));
    LocalMux I__1457 (
            .O(N__13431),
            .I(\c0.rx.n4011 ));
    Odrv4 I__1456 (
            .O(N__13428),
            .I(\c0.rx.n4011 ));
    InMux I__1455 (
            .O(N__13423),
            .I(N__13419));
    InMux I__1454 (
            .O(N__13422),
            .I(N__13416));
    LocalMux I__1453 (
            .O(N__13419),
            .I(N__13411));
    LocalMux I__1452 (
            .O(N__13416),
            .I(N__13411));
    Span4Mux_v I__1451 (
            .O(N__13411),
            .I(N__13407));
    InMux I__1450 (
            .O(N__13410),
            .I(N__13404));
    Odrv4 I__1449 (
            .O(N__13407),
            .I(data_in_5_1));
    LocalMux I__1448 (
            .O(N__13404),
            .I(data_in_5_1));
    InMux I__1447 (
            .O(N__13399),
            .I(N__13393));
    InMux I__1446 (
            .O(N__13398),
            .I(N__13390));
    InMux I__1445 (
            .O(N__13397),
            .I(N__13387));
    InMux I__1444 (
            .O(N__13396),
            .I(N__13384));
    LocalMux I__1443 (
            .O(N__13393),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__1442 (
            .O(N__13390),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__1441 (
            .O(N__13387),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__1440 (
            .O(N__13384),
            .I(\c0.rx.r_Clock_Count_5 ));
    InMux I__1439 (
            .O(N__13375),
            .I(N__13369));
    InMux I__1438 (
            .O(N__13374),
            .I(N__13366));
    InMux I__1437 (
            .O(N__13373),
            .I(N__13363));
    InMux I__1436 (
            .O(N__13372),
            .I(N__13360));
    LocalMux I__1435 (
            .O(N__13369),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__1434 (
            .O(N__13366),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__1433 (
            .O(N__13363),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__1432 (
            .O(N__13360),
            .I(\c0.rx.r_Clock_Count_4 ));
    InMux I__1431 (
            .O(N__13351),
            .I(N__13348));
    LocalMux I__1430 (
            .O(N__13348),
            .I(\c0.rx.n37 ));
    InMux I__1429 (
            .O(N__13345),
            .I(N__13341));
    InMux I__1428 (
            .O(N__13344),
            .I(N__13335));
    LocalMux I__1427 (
            .O(N__13341),
            .I(N__13332));
    InMux I__1426 (
            .O(N__13340),
            .I(N__13329));
    InMux I__1425 (
            .O(N__13339),
            .I(N__13326));
    InMux I__1424 (
            .O(N__13338),
            .I(N__13323));
    LocalMux I__1423 (
            .O(N__13335),
            .I(\c0.rx.r_Clock_Count_1 ));
    Odrv4 I__1422 (
            .O(N__13332),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__1421 (
            .O(N__13329),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__1420 (
            .O(N__13326),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__1419 (
            .O(N__13323),
            .I(\c0.rx.r_Clock_Count_1 ));
    CascadeMux I__1418 (
            .O(N__13312),
            .I(\c0.rx.n37_cascade_ ));
    InMux I__1417 (
            .O(N__13309),
            .I(N__13302));
    InMux I__1416 (
            .O(N__13308),
            .I(N__13299));
    InMux I__1415 (
            .O(N__13307),
            .I(N__13296));
    InMux I__1414 (
            .O(N__13306),
            .I(N__13291));
    InMux I__1413 (
            .O(N__13305),
            .I(N__13291));
    LocalMux I__1412 (
            .O(N__13302),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__1411 (
            .O(N__13299),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__1410 (
            .O(N__13296),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__1409 (
            .O(N__13291),
            .I(\c0.rx.r_Clock_Count_3 ));
    InMux I__1408 (
            .O(N__13282),
            .I(N__13275));
    InMux I__1407 (
            .O(N__13281),
            .I(N__13272));
    InMux I__1406 (
            .O(N__13280),
            .I(N__13265));
    InMux I__1405 (
            .O(N__13279),
            .I(N__13265));
    InMux I__1404 (
            .O(N__13278),
            .I(N__13265));
    LocalMux I__1403 (
            .O(N__13275),
            .I(r_SM_Main_2_N_1830_0));
    LocalMux I__1402 (
            .O(N__13272),
            .I(r_SM_Main_2_N_1830_0));
    LocalMux I__1401 (
            .O(N__13265),
            .I(r_SM_Main_2_N_1830_0));
    InMux I__1400 (
            .O(N__13258),
            .I(N__13255));
    LocalMux I__1399 (
            .O(N__13255),
            .I(\c0.rx.r_Rx_Data_R ));
    CascadeMux I__1398 (
            .O(N__13252),
            .I(n12_adj_1995_cascade_));
    InMux I__1397 (
            .O(N__13249),
            .I(N__13246));
    LocalMux I__1396 (
            .O(N__13246),
            .I(n5316));
    InMux I__1395 (
            .O(N__13243),
            .I(N__13233));
    InMux I__1394 (
            .O(N__13242),
            .I(N__13233));
    InMux I__1393 (
            .O(N__13241),
            .I(N__13226));
    InMux I__1392 (
            .O(N__13240),
            .I(N__13226));
    InMux I__1391 (
            .O(N__13239),
            .I(N__13226));
    InMux I__1390 (
            .O(N__13238),
            .I(N__13219));
    LocalMux I__1389 (
            .O(N__13233),
            .I(N__13216));
    LocalMux I__1388 (
            .O(N__13226),
            .I(N__13213));
    InMux I__1387 (
            .O(N__13225),
            .I(N__13206));
    InMux I__1386 (
            .O(N__13224),
            .I(N__13206));
    InMux I__1385 (
            .O(N__13223),
            .I(N__13206));
    InMux I__1384 (
            .O(N__13222),
            .I(N__13203));
    LocalMux I__1383 (
            .O(N__13219),
            .I(n16_adj_1993));
    Odrv12 I__1382 (
            .O(N__13216),
            .I(n16_adj_1993));
    Odrv4 I__1381 (
            .O(N__13213),
            .I(n16_adj_1993));
    LocalMux I__1380 (
            .O(N__13206),
            .I(n16_adj_1993));
    LocalMux I__1379 (
            .O(N__13203),
            .I(n16_adj_1993));
    InMux I__1378 (
            .O(N__13192),
            .I(N__13189));
    LocalMux I__1377 (
            .O(N__13189),
            .I(n5491));
    InMux I__1376 (
            .O(N__13186),
            .I(N__13183));
    LocalMux I__1375 (
            .O(N__13183),
            .I(\c0.rx.n5535 ));
    InMux I__1374 (
            .O(N__13180),
            .I(N__13177));
    LocalMux I__1373 (
            .O(N__13177),
            .I(\c0.rx.n2157 ));
    InMux I__1372 (
            .O(N__13174),
            .I(N__13171));
    LocalMux I__1371 (
            .O(N__13171),
            .I(\c0.rx.n5538 ));
    InMux I__1370 (
            .O(N__13168),
            .I(N__13165));
    LocalMux I__1369 (
            .O(N__13165),
            .I(\c0.rx.n5539 ));
    InMux I__1368 (
            .O(N__13162),
            .I(N__13159));
    LocalMux I__1367 (
            .O(N__13159),
            .I(\c0.rx.n40 ));
    CascadeMux I__1366 (
            .O(N__13156),
            .I(\c0.rx.r_SM_Main_2_N_1824_2_cascade_ ));
    InMux I__1365 (
            .O(N__13153),
            .I(N__13150));
    LocalMux I__1364 (
            .O(N__13150),
            .I(n4474));
    InMux I__1363 (
            .O(N__13147),
            .I(N__13144));
    LocalMux I__1362 (
            .O(N__13144),
            .I(n2156));
    CascadeMux I__1361 (
            .O(N__13141),
            .I(n4474_cascade_));
    InMux I__1360 (
            .O(N__13138),
            .I(N__13134));
    InMux I__1359 (
            .O(N__13137),
            .I(N__13131));
    LocalMux I__1358 (
            .O(N__13134),
            .I(N__13128));
    LocalMux I__1357 (
            .O(N__13131),
            .I(\c0.data_in_frame_18_1 ));
    Odrv4 I__1356 (
            .O(N__13128),
            .I(\c0.data_in_frame_18_1 ));
    InMux I__1355 (
            .O(N__13123),
            .I(N__13120));
    LocalMux I__1354 (
            .O(N__13120),
            .I(N__13117));
    Odrv4 I__1353 (
            .O(N__13117),
            .I(\c0.n5369 ));
    InMux I__1352 (
            .O(N__13114),
            .I(N__13111));
    LocalMux I__1351 (
            .O(N__13111),
            .I(N__13108));
    Odrv4 I__1350 (
            .O(N__13108),
            .I(\c0.n5869 ));
    CascadeMux I__1349 (
            .O(N__13105),
            .I(N__13102));
    InMux I__1348 (
            .O(N__13102),
            .I(N__13099));
    LocalMux I__1347 (
            .O(N__13099),
            .I(\c0.n5959 ));
    CascadeMux I__1346 (
            .O(N__13096),
            .I(N__13093));
    InMux I__1345 (
            .O(N__13093),
            .I(N__13090));
    LocalMux I__1344 (
            .O(N__13090),
            .I(N__13087));
    Odrv12 I__1343 (
            .O(N__13087),
            .I(\c0.n5962 ));
    InMux I__1342 (
            .O(N__13084),
            .I(N__13080));
    InMux I__1341 (
            .O(N__13083),
            .I(N__13077));
    LocalMux I__1340 (
            .O(N__13080),
            .I(N__13074));
    LocalMux I__1339 (
            .O(N__13077),
            .I(\c0.data_in_frame_18_3 ));
    Odrv4 I__1338 (
            .O(N__13074),
            .I(\c0.data_in_frame_18_3 ));
    InMux I__1337 (
            .O(N__13069),
            .I(N__13066));
    LocalMux I__1336 (
            .O(N__13066),
            .I(n5051));
    CascadeMux I__1335 (
            .O(N__13063),
            .I(\c0.n5725_cascade_ ));
    InMux I__1334 (
            .O(N__13060),
            .I(N__13049));
    InMux I__1333 (
            .O(N__13059),
            .I(N__13049));
    InMux I__1332 (
            .O(N__13058),
            .I(N__13049));
    InMux I__1331 (
            .O(N__13057),
            .I(N__13042));
    InMux I__1330 (
            .O(N__13056),
            .I(N__13039));
    LocalMux I__1329 (
            .O(N__13049),
            .I(N__13036));
    InMux I__1328 (
            .O(N__13048),
            .I(N__13029));
    InMux I__1327 (
            .O(N__13047),
            .I(N__13029));
    InMux I__1326 (
            .O(N__13046),
            .I(N__13029));
    InMux I__1325 (
            .O(N__13045),
            .I(N__13026));
    LocalMux I__1324 (
            .O(N__13042),
            .I(N__13021));
    LocalMux I__1323 (
            .O(N__13039),
            .I(N__13021));
    Odrv4 I__1322 (
            .O(N__13036),
            .I(\c0.n1058 ));
    LocalMux I__1321 (
            .O(N__13029),
            .I(\c0.n1058 ));
    LocalMux I__1320 (
            .O(N__13026),
            .I(\c0.n1058 ));
    Odrv4 I__1319 (
            .O(N__13021),
            .I(\c0.n1058 ));
    CascadeMux I__1318 (
            .O(N__13012),
            .I(\c0.n5728_cascade_ ));
    InMux I__1317 (
            .O(N__13009),
            .I(N__13006));
    LocalMux I__1316 (
            .O(N__13006),
            .I(\c0.n5974 ));
    InMux I__1315 (
            .O(N__13003),
            .I(N__13000));
    LocalMux I__1314 (
            .O(N__13000),
            .I(N__12997));
    Odrv4 I__1313 (
            .O(N__12997),
            .I(\c0.tx2.r_Tx_Data_1 ));
    CEMux I__1312 (
            .O(N__12994),
            .I(N__12989));
    CEMux I__1311 (
            .O(N__12993),
            .I(N__12986));
    CEMux I__1310 (
            .O(N__12992),
            .I(N__12983));
    LocalMux I__1309 (
            .O(N__12989),
            .I(N__12977));
    LocalMux I__1308 (
            .O(N__12986),
            .I(N__12977));
    LocalMux I__1307 (
            .O(N__12983),
            .I(N__12974));
    CEMux I__1306 (
            .O(N__12982),
            .I(N__12971));
    Span4Mux_v I__1305 (
            .O(N__12977),
            .I(N__12968));
    Span4Mux_s1_h I__1304 (
            .O(N__12974),
            .I(N__12963));
    LocalMux I__1303 (
            .O(N__12971),
            .I(N__12963));
    Odrv4 I__1302 (
            .O(N__12968),
            .I(\c0.tx2.n1592 ));
    Odrv4 I__1301 (
            .O(N__12963),
            .I(\c0.tx2.n1592 ));
    CascadeMux I__1300 (
            .O(N__12958),
            .I(\c0.n5803_cascade_ ));
    InMux I__1299 (
            .O(N__12955),
            .I(N__12952));
    LocalMux I__1298 (
            .O(N__12952),
            .I(\c0.tx2.r_Tx_Data_3 ));
    CascadeMux I__1297 (
            .O(N__12949),
            .I(\c0.n5665_cascade_ ));
    CascadeMux I__1296 (
            .O(N__12946),
            .I(\c0.n5372_cascade_ ));
    InMux I__1295 (
            .O(N__12943),
            .I(N__12940));
    LocalMux I__1294 (
            .O(N__12940),
            .I(\c0.n5659 ));
    CascadeMux I__1293 (
            .O(N__12937),
            .I(N__12934));
    InMux I__1292 (
            .O(N__12934),
            .I(N__12931));
    LocalMux I__1291 (
            .O(N__12931),
            .I(\c0.n5938 ));
    CascadeMux I__1290 (
            .O(N__12928),
            .I(\c0.n5971_cascade_ ));
    CascadeMux I__1289 (
            .O(N__12925),
            .I(N__12922));
    InMux I__1288 (
            .O(N__12922),
            .I(N__12919));
    LocalMux I__1287 (
            .O(N__12919),
            .I(\c0.tx2.r_Tx_Data_0 ));
    InMux I__1286 (
            .O(N__12916),
            .I(N__12913));
    LocalMux I__1285 (
            .O(N__12913),
            .I(\c0.tx2.n5947 ));
    InMux I__1284 (
            .O(N__12910),
            .I(N__12907));
    LocalMux I__1283 (
            .O(N__12907),
            .I(\c0.tx2.n5950 ));
    InMux I__1282 (
            .O(N__12904),
            .I(N__12901));
    LocalMux I__1281 (
            .O(N__12901),
            .I(n1345));
    InMux I__1280 (
            .O(N__12898),
            .I(N__12895));
    LocalMux I__1279 (
            .O(N__12895),
            .I(\c0.tx2.r_Tx_Data_4 ));
    InMux I__1278 (
            .O(N__12892),
            .I(N__12889));
    LocalMux I__1277 (
            .O(N__12889),
            .I(\c0.tx2.r_Tx_Data_2 ));
    CascadeMux I__1276 (
            .O(N__12886),
            .I(N__12881));
    InMux I__1275 (
            .O(N__12885),
            .I(N__12878));
    InMux I__1274 (
            .O(N__12884),
            .I(N__12875));
    InMux I__1273 (
            .O(N__12881),
            .I(N__12872));
    LocalMux I__1272 (
            .O(N__12878),
            .I(\c0.tx2.r_Clock_Count_1 ));
    LocalMux I__1271 (
            .O(N__12875),
            .I(\c0.tx2.r_Clock_Count_1 ));
    LocalMux I__1270 (
            .O(N__12872),
            .I(\c0.tx2.r_Clock_Count_1 ));
    InMux I__1269 (
            .O(N__12865),
            .I(N__12862));
    LocalMux I__1268 (
            .O(N__12862),
            .I(n2399));
    InMux I__1267 (
            .O(N__12859),
            .I(\c0.tx2.n4429 ));
    InMux I__1266 (
            .O(N__12856),
            .I(\c0.tx2.n4430 ));
    InMux I__1265 (
            .O(N__12853),
            .I(\c0.tx2.n4431 ));
    InMux I__1264 (
            .O(N__12850),
            .I(N__12845));
    InMux I__1263 (
            .O(N__12849),
            .I(N__12842));
    InMux I__1262 (
            .O(N__12848),
            .I(N__12839));
    LocalMux I__1261 (
            .O(N__12845),
            .I(\c0.tx2.r_Clock_Count_4 ));
    LocalMux I__1260 (
            .O(N__12842),
            .I(\c0.tx2.r_Clock_Count_4 ));
    LocalMux I__1259 (
            .O(N__12839),
            .I(\c0.tx2.r_Clock_Count_4 ));
    InMux I__1258 (
            .O(N__12832),
            .I(N__12829));
    LocalMux I__1257 (
            .O(N__12829),
            .I(N__12826));
    Odrv4 I__1256 (
            .O(N__12826),
            .I(n2382));
    InMux I__1255 (
            .O(N__12823),
            .I(\c0.tx2.n4432 ));
    InMux I__1254 (
            .O(N__12820),
            .I(N__12815));
    InMux I__1253 (
            .O(N__12819),
            .I(N__12812));
    InMux I__1252 (
            .O(N__12818),
            .I(N__12809));
    LocalMux I__1251 (
            .O(N__12815),
            .I(\c0.tx2.r_Clock_Count_5 ));
    LocalMux I__1250 (
            .O(N__12812),
            .I(\c0.tx2.r_Clock_Count_5 ));
    LocalMux I__1249 (
            .O(N__12809),
            .I(\c0.tx2.r_Clock_Count_5 ));
    InMux I__1248 (
            .O(N__12802),
            .I(N__12799));
    LocalMux I__1247 (
            .O(N__12799),
            .I(N__12796));
    Odrv4 I__1246 (
            .O(N__12796),
            .I(n2379));
    InMux I__1245 (
            .O(N__12793),
            .I(\c0.tx2.n4433 ));
    InMux I__1244 (
            .O(N__12790),
            .I(N__12785));
    InMux I__1243 (
            .O(N__12789),
            .I(N__12782));
    InMux I__1242 (
            .O(N__12788),
            .I(N__12779));
    LocalMux I__1241 (
            .O(N__12785),
            .I(\c0.tx2.r_Clock_Count_6 ));
    LocalMux I__1240 (
            .O(N__12782),
            .I(\c0.tx2.r_Clock_Count_6 ));
    LocalMux I__1239 (
            .O(N__12779),
            .I(\c0.tx2.r_Clock_Count_6 ));
    InMux I__1238 (
            .O(N__12772),
            .I(N__12769));
    LocalMux I__1237 (
            .O(N__12769),
            .I(N__12766));
    Odrv4 I__1236 (
            .O(N__12766),
            .I(n2376));
    InMux I__1235 (
            .O(N__12763),
            .I(\c0.tx2.n4434 ));
    InMux I__1234 (
            .O(N__12760),
            .I(\c0.tx2.n4435 ));
    InMux I__1233 (
            .O(N__12757),
            .I(N__12752));
    InMux I__1232 (
            .O(N__12756),
            .I(N__12749));
    InMux I__1231 (
            .O(N__12755),
            .I(N__12745));
    LocalMux I__1230 (
            .O(N__12752),
            .I(N__12740));
    LocalMux I__1229 (
            .O(N__12749),
            .I(N__12740));
    InMux I__1228 (
            .O(N__12748),
            .I(N__12737));
    LocalMux I__1227 (
            .O(N__12745),
            .I(r_Clock_Count_8_adj_2012));
    Odrv4 I__1226 (
            .O(N__12740),
            .I(r_Clock_Count_8_adj_2012));
    LocalMux I__1225 (
            .O(N__12737),
            .I(r_Clock_Count_8_adj_2012));
    InMux I__1224 (
            .O(N__12730),
            .I(bfn_2_24_0_));
    InMux I__1223 (
            .O(N__12727),
            .I(N__12724));
    LocalMux I__1222 (
            .O(N__12724),
            .I(N__12721));
    Odrv4 I__1221 (
            .O(N__12721),
            .I(n2369));
    CascadeMux I__1220 (
            .O(N__12718),
            .I(\c0.tx2.n5_cascade_ ));
    InMux I__1219 (
            .O(N__12715),
            .I(N__12712));
    LocalMux I__1218 (
            .O(N__12712),
            .I(\c0.tx2.n3591 ));
    CascadeMux I__1217 (
            .O(N__12709),
            .I(\c0.tx2.n3591_cascade_ ));
    CascadeMux I__1216 (
            .O(N__12706),
            .I(r_SM_Main_2_N_1767_1_cascade_));
    InMux I__1215 (
            .O(N__12703),
            .I(N__12699));
    InMux I__1214 (
            .O(N__12702),
            .I(N__12696));
    LocalMux I__1213 (
            .O(N__12699),
            .I(N__12691));
    LocalMux I__1212 (
            .O(N__12696),
            .I(N__12691));
    Odrv4 I__1211 (
            .O(N__12691),
            .I(\c0.tx2.r_Clock_Count_0 ));
    CascadeMux I__1210 (
            .O(N__12688),
            .I(N__12685));
    InMux I__1209 (
            .O(N__12685),
            .I(N__12682));
    LocalMux I__1208 (
            .O(N__12682),
            .I(n2460));
    InMux I__1207 (
            .O(N__12679),
            .I(bfn_2_23_0_));
    CascadeMux I__1206 (
            .O(N__12676),
            .I(N__12673));
    InMux I__1205 (
            .O(N__12673),
            .I(N__12669));
    InMux I__1204 (
            .O(N__12672),
            .I(N__12666));
    LocalMux I__1203 (
            .O(N__12669),
            .I(\c0.tx.r_Clock_Count_0 ));
    LocalMux I__1202 (
            .O(N__12666),
            .I(\c0.tx.r_Clock_Count_0 ));
    InMux I__1201 (
            .O(N__12661),
            .I(N__12658));
    LocalMux I__1200 (
            .O(N__12658),
            .I(\c0.tx.n313 ));
    InMux I__1199 (
            .O(N__12655),
            .I(N__12652));
    LocalMux I__1198 (
            .O(N__12652),
            .I(n316));
    InMux I__1197 (
            .O(N__12649),
            .I(N__12646));
    LocalMux I__1196 (
            .O(N__12646),
            .I(n314));
    CascadeMux I__1195 (
            .O(N__12643),
            .I(N__12640));
    InMux I__1194 (
            .O(N__12640),
            .I(N__12637));
    LocalMux I__1193 (
            .O(N__12637),
            .I(n317));
    CascadeMux I__1192 (
            .O(N__12634),
            .I(N__12631));
    InMux I__1191 (
            .O(N__12631),
            .I(N__12626));
    InMux I__1190 (
            .O(N__12630),
            .I(N__12623));
    InMux I__1189 (
            .O(N__12629),
            .I(N__12620));
    LocalMux I__1188 (
            .O(N__12626),
            .I(r_Clock_Count_2));
    LocalMux I__1187 (
            .O(N__12623),
            .I(r_Clock_Count_2));
    LocalMux I__1186 (
            .O(N__12620),
            .I(r_Clock_Count_2));
    InMux I__1185 (
            .O(N__12613),
            .I(N__12608));
    InMux I__1184 (
            .O(N__12612),
            .I(N__12605));
    InMux I__1183 (
            .O(N__12611),
            .I(N__12602));
    LocalMux I__1182 (
            .O(N__12608),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__1181 (
            .O(N__12605),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__1180 (
            .O(N__12602),
            .I(\c0.tx.r_Clock_Count_6 ));
    CascadeMux I__1179 (
            .O(N__12595),
            .I(N__12591));
    CascadeMux I__1178 (
            .O(N__12594),
            .I(N__12587));
    InMux I__1177 (
            .O(N__12591),
            .I(N__12584));
    InMux I__1176 (
            .O(N__12590),
            .I(N__12581));
    InMux I__1175 (
            .O(N__12587),
            .I(N__12578));
    LocalMux I__1174 (
            .O(N__12584),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__1173 (
            .O(N__12581),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__1172 (
            .O(N__12578),
            .I(\c0.tx.r_Clock_Count_1 ));
    InMux I__1171 (
            .O(N__12571),
            .I(N__12566));
    InMux I__1170 (
            .O(N__12570),
            .I(N__12561));
    InMux I__1169 (
            .O(N__12569),
            .I(N__12561));
    LocalMux I__1168 (
            .O(N__12566),
            .I(r_Clock_Count_5));
    LocalMux I__1167 (
            .O(N__12561),
            .I(r_Clock_Count_5));
    InMux I__1166 (
            .O(N__12556),
            .I(N__12551));
    InMux I__1165 (
            .O(N__12555),
            .I(N__12546));
    InMux I__1164 (
            .O(N__12554),
            .I(N__12546));
    LocalMux I__1163 (
            .O(N__12551),
            .I(r_Clock_Count_4));
    LocalMux I__1162 (
            .O(N__12546),
            .I(r_Clock_Count_4));
    CascadeMux I__1161 (
            .O(N__12541),
            .I(\c0.tx.n5_cascade_ ));
    InMux I__1160 (
            .O(N__12538),
            .I(N__12533));
    InMux I__1159 (
            .O(N__12537),
            .I(N__12528));
    InMux I__1158 (
            .O(N__12536),
            .I(N__12528));
    LocalMux I__1157 (
            .O(N__12533),
            .I(r_Clock_Count_7));
    LocalMux I__1156 (
            .O(N__12528),
            .I(r_Clock_Count_7));
    CascadeMux I__1155 (
            .O(N__12523),
            .I(n3595_cascade_));
    CascadeMux I__1154 (
            .O(N__12520),
            .I(N__12517));
    InMux I__1153 (
            .O(N__12517),
            .I(N__12514));
    LocalMux I__1152 (
            .O(N__12514),
            .I(\c0.tx.n5520 ));
    InMux I__1151 (
            .O(N__12511),
            .I(N__12506));
    InMux I__1150 (
            .O(N__12510),
            .I(N__12501));
    InMux I__1149 (
            .O(N__12509),
            .I(N__12501));
    LocalMux I__1148 (
            .O(N__12506),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__1147 (
            .O(N__12501),
            .I(\c0.tx.r_Clock_Count_3 ));
    InMux I__1146 (
            .O(N__12496),
            .I(N__12493));
    LocalMux I__1145 (
            .O(N__12493),
            .I(n1760));
    CascadeMux I__1144 (
            .O(N__12490),
            .I(\c0.n1529_cascade_ ));
    InMux I__1143 (
            .O(N__12487),
            .I(N__12484));
    LocalMux I__1142 (
            .O(N__12484),
            .I(\c0.n1801 ));
    InMux I__1141 (
            .O(N__12481),
            .I(N__12478));
    LocalMux I__1140 (
            .O(N__12478),
            .I(\c0.tx.n315 ));
    InMux I__1139 (
            .O(N__12475),
            .I(N__12472));
    LocalMux I__1138 (
            .O(N__12472),
            .I(n319));
    InMux I__1137 (
            .O(N__12469),
            .I(N__12466));
    LocalMux I__1136 (
            .O(N__12466),
            .I(\c0.tx.n320 ));
    InMux I__1135 (
            .O(N__12463),
            .I(N__12460));
    LocalMux I__1134 (
            .O(N__12460),
            .I(\c0.tx.n321 ));
    InMux I__1133 (
            .O(N__12457),
            .I(N__12454));
    LocalMux I__1132 (
            .O(N__12454),
            .I(\c0.n50 ));
    InMux I__1131 (
            .O(N__12451),
            .I(N__12448));
    LocalMux I__1130 (
            .O(N__12448),
            .I(\c0.tx_active_prev ));
    CascadeMux I__1129 (
            .O(N__12445),
            .I(\c0.n5540_cascade_ ));
    CascadeMux I__1128 (
            .O(N__12442),
            .I(\c0.n5977_cascade_ ));
    CascadeMux I__1127 (
            .O(N__12439),
            .I(n1760_cascade_));
    InMux I__1126 (
            .O(N__12436),
            .I(\c0.n4378 ));
    InMux I__1125 (
            .O(N__12433),
            .I(N__12427));
    InMux I__1124 (
            .O(N__12432),
            .I(N__12427));
    LocalMux I__1123 (
            .O(N__12427),
            .I(\c0.tx_transmit_N_568_2 ));
    InMux I__1122 (
            .O(N__12424),
            .I(\c0.n4379 ));
    InMux I__1121 (
            .O(N__12421),
            .I(N__12415));
    InMux I__1120 (
            .O(N__12420),
            .I(N__12415));
    LocalMux I__1119 (
            .O(N__12415),
            .I(\c0.tx_transmit_N_568_3 ));
    InMux I__1118 (
            .O(N__12412),
            .I(\c0.n4380 ));
    InMux I__1117 (
            .O(N__12409),
            .I(\c0.n4381 ));
    InMux I__1116 (
            .O(N__12406),
            .I(N__12403));
    LocalMux I__1115 (
            .O(N__12403),
            .I(\c0.byte_transmit_counter_5 ));
    InMux I__1114 (
            .O(N__12400),
            .I(\c0.n4382 ));
    InMux I__1113 (
            .O(N__12397),
            .I(N__12394));
    LocalMux I__1112 (
            .O(N__12394),
            .I(\c0.byte_transmit_counter_6 ));
    InMux I__1111 (
            .O(N__12391),
            .I(\c0.n4383 ));
    InMux I__1110 (
            .O(N__12388),
            .I(N__12385));
    LocalMux I__1109 (
            .O(N__12385),
            .I(\c0.byte_transmit_counter_7 ));
    InMux I__1108 (
            .O(N__12382),
            .I(\c0.n4384 ));
    InMux I__1107 (
            .O(N__12379),
            .I(N__12376));
    LocalMux I__1106 (
            .O(N__12376),
            .I(n5490));
    CascadeMux I__1105 (
            .O(N__12373),
            .I(\c0.rx.n3980_cascade_ ));
    InMux I__1104 (
            .O(N__12370),
            .I(N__12367));
    LocalMux I__1103 (
            .O(N__12367),
            .I(\c0.rx.n5532 ));
    CascadeMux I__1102 (
            .O(N__12364),
            .I(\c0.rx.n5298_cascade_ ));
    InMux I__1101 (
            .O(N__12361),
            .I(N__12358));
    LocalMux I__1100 (
            .O(N__12358),
            .I(\c0.rx.n5536 ));
    InMux I__1099 (
            .O(N__12355),
            .I(N__12349));
    InMux I__1098 (
            .O(N__12354),
            .I(N__12349));
    LocalMux I__1097 (
            .O(N__12349),
            .I(\c0.rx.n5049 ));
    InMux I__1096 (
            .O(N__12346),
            .I(N__12343));
    LocalMux I__1095 (
            .O(N__12343),
            .I(n5050));
    CascadeMux I__1094 (
            .O(N__12340),
            .I(\c0.rx.n5923_cascade_ ));
    CascadeMux I__1093 (
            .O(N__12337),
            .I(\c0.rx.n5926_cascade_ ));
    InMux I__1092 (
            .O(N__12334),
            .I(N__12331));
    LocalMux I__1091 (
            .O(N__12331),
            .I(N__12328));
    Odrv4 I__1090 (
            .O(N__12328),
            .I(\c0.rx.n5537 ));
    InMux I__1089 (
            .O(N__12325),
            .I(\c0.rx.n4422 ));
    InMux I__1088 (
            .O(N__12322),
            .I(\c0.rx.n4423 ));
    InMux I__1087 (
            .O(N__12319),
            .I(\c0.rx.n4424 ));
    InMux I__1086 (
            .O(N__12316),
            .I(\c0.rx.n4425 ));
    InMux I__1085 (
            .O(N__12313),
            .I(\c0.rx.n4426 ));
    InMux I__1084 (
            .O(N__12310),
            .I(\c0.rx.n4427 ));
    InMux I__1083 (
            .O(N__12307),
            .I(\c0.rx.n4428 ));
    CascadeMux I__1082 (
            .O(N__12304),
            .I(n2156_cascade_));
    InMux I__1081 (
            .O(N__12301),
            .I(N__12298));
    LocalMux I__1080 (
            .O(N__12298),
            .I(n8));
    CascadeMux I__1079 (
            .O(N__12295),
            .I(N__12292));
    InMux I__1078 (
            .O(N__12292),
            .I(N__12288));
    InMux I__1077 (
            .O(N__12291),
            .I(N__12285));
    LocalMux I__1076 (
            .O(N__12288),
            .I(N__12282));
    LocalMux I__1075 (
            .O(N__12285),
            .I(\c0.data_in_frame_19_0 ));
    Odrv12 I__1074 (
            .O(N__12282),
            .I(\c0.data_in_frame_19_0 ));
    InMux I__1073 (
            .O(N__12277),
            .I(N__12272));
    IoInMux I__1072 (
            .O(N__12276),
            .I(N__12269));
    InMux I__1071 (
            .O(N__12275),
            .I(N__12266));
    LocalMux I__1070 (
            .O(N__12272),
            .I(N__12263));
    LocalMux I__1069 (
            .O(N__12269),
            .I(tx2_o));
    LocalMux I__1068 (
            .O(N__12266),
            .I(tx2_o));
    Odrv4 I__1067 (
            .O(N__12263),
            .I(tx2_o));
    IoInMux I__1066 (
            .O(N__12256),
            .I(N__12253));
    LocalMux I__1065 (
            .O(N__12253),
            .I(tx2_enable));
    InMux I__1064 (
            .O(N__12250),
            .I(N__12247));
    LocalMux I__1063 (
            .O(N__12247),
            .I(\c0.n5402 ));
    CascadeMux I__1062 (
            .O(N__12244),
            .I(N__12240));
    InMux I__1061 (
            .O(N__12243),
            .I(N__12237));
    InMux I__1060 (
            .O(N__12240),
            .I(N__12234));
    LocalMux I__1059 (
            .O(N__12237),
            .I(\c0.data_in_frame_19_3 ));
    LocalMux I__1058 (
            .O(N__12234),
            .I(\c0.data_in_frame_19_3 ));
    InMux I__1057 (
            .O(N__12229),
            .I(N__12226));
    LocalMux I__1056 (
            .O(N__12226),
            .I(\c0.n5863 ));
    InMux I__1055 (
            .O(N__12223),
            .I(bfn_1_30_0_));
    CascadeMux I__1054 (
            .O(N__12220),
            .I(\c0.n5920_cascade_ ));
    InMux I__1053 (
            .O(N__12217),
            .I(N__12214));
    LocalMux I__1052 (
            .O(N__12214),
            .I(\c0.n5662 ));
    CascadeMux I__1051 (
            .O(N__12211),
            .I(N__12208));
    InMux I__1050 (
            .O(N__12208),
            .I(N__12205));
    LocalMux I__1049 (
            .O(N__12205),
            .I(\c0.tx2.r_Tx_Data_7 ));
    InMux I__1048 (
            .O(N__12202),
            .I(N__12199));
    LocalMux I__1047 (
            .O(N__12199),
            .I(\c0.tx2.n5929 ));
    InMux I__1046 (
            .O(N__12196),
            .I(N__12193));
    LocalMux I__1045 (
            .O(N__12193),
            .I(\c0.tx2.r_Tx_Data_6 ));
    InMux I__1044 (
            .O(N__12190),
            .I(N__12187));
    LocalMux I__1043 (
            .O(N__12187),
            .I(N__12184));
    Odrv4 I__1042 (
            .O(N__12184),
            .I(\c0.tx2.r_Tx_Data_5 ));
    CascadeMux I__1041 (
            .O(N__12181),
            .I(\c0.n5399_cascade_ ));
    CascadeMux I__1040 (
            .O(N__12178),
            .I(\c0.n5857_cascade_ ));
    InMux I__1039 (
            .O(N__12175),
            .I(N__12172));
    LocalMux I__1038 (
            .O(N__12172),
            .I(\c0.n5860 ));
    InMux I__1037 (
            .O(N__12169),
            .I(N__12166));
    LocalMux I__1036 (
            .O(N__12166),
            .I(N__12163));
    Odrv4 I__1035 (
            .O(N__12163),
            .I(\c0.tx2.o_Tx_Serial_N_1798 ));
    CascadeMux I__1034 (
            .O(N__12160),
            .I(n3_cascade_));
    CascadeMux I__1033 (
            .O(N__12157),
            .I(\c0.tx2.n5312_cascade_ ));
    CascadeMux I__1032 (
            .O(N__12154),
            .I(\c0.n5815_cascade_ ));
    CascadeMux I__1031 (
            .O(N__12151),
            .I(N__12148));
    InMux I__1030 (
            .O(N__12148),
            .I(N__12145));
    LocalMux I__1029 (
            .O(N__12145),
            .I(\c0.n5818 ));
    CascadeMux I__1028 (
            .O(N__12142),
            .I(\c0.tx2.n5932_cascade_ ));
    CascadeMux I__1027 (
            .O(N__12139),
            .I(\c0.n5917_cascade_ ));
    InMux I__1026 (
            .O(N__12136),
            .I(\c0.tx.n4420 ));
    InMux I__1025 (
            .O(N__12133),
            .I(bfn_1_22_0_));
    CascadeMux I__1024 (
            .O(N__12130),
            .I(n5037_cascade_));
    InMux I__1023 (
            .O(N__12127),
            .I(N__12124));
    LocalMux I__1022 (
            .O(N__12124),
            .I(n3611));
    CascadeMux I__1021 (
            .O(N__12121),
            .I(n4_adj_2008_cascade_));
    InMux I__1020 (
            .O(N__12118),
            .I(bfn_1_21_0_));
    InMux I__1019 (
            .O(N__12115),
            .I(\c0.tx.n4414 ));
    InMux I__1018 (
            .O(N__12112),
            .I(\c0.tx.n4415 ));
    InMux I__1017 (
            .O(N__12109),
            .I(\c0.tx.n4416 ));
    InMux I__1016 (
            .O(N__12106),
            .I(\c0.tx.n4417 ));
    InMux I__1015 (
            .O(N__12103),
            .I(\c0.tx.n4418 ));
    InMux I__1014 (
            .O(N__12100),
            .I(\c0.tx.n4419 ));
    IoInMux I__1013 (
            .O(N__12097),
            .I(N__12094));
    LocalMux I__1012 (
            .O(N__12094),
            .I(N__12091));
    IoSpan4Mux I__1011 (
            .O(N__12091),
            .I(N__12088));
    IoSpan4Mux I__1010 (
            .O(N__12088),
            .I(N__12085));
    IoSpan4Mux I__1009 (
            .O(N__12085),
            .I(N__12082));
    Odrv4 I__1008 (
            .O(N__12082),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_2_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_23_0_));
    defparam IN_MUX_bfv_2_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_24_0_ (
            .carryinitin(\c0.tx2.n4436 ),
            .carryinitout(bfn_2_24_0_));
    defparam IN_MUX_bfv_1_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_21_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(\c0.tx.n4421 ),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_1_30_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_30_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_4_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_17_0_ (
            .carryinitin(\c0.n4411 ),
            .carryinitout(bfn_4_17_0_));
    defparam IN_MUX_bfv_6_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_17_0_));
    defparam IN_MUX_bfv_6_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_18_0_ (
            .carryinitin(\c0.n4392 ),
            .carryinitout(bfn_6_18_0_));
    defparam IN_MUX_bfv_3_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_24_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(n4444),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_15_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_27_0_ (
            .carryinitin(n4452),
            .carryinitout(bfn_15_27_0_));
    defparam IN_MUX_bfv_15_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_28_0_ (
            .carryinitin(n4460),
            .carryinitout(bfn_15_28_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__12097),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_937_LC_1_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_937_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_937_LC_1_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_937_LC_1_19_2  (
            .in0(N__18977),
            .in1(N__20475),
            .in2(_gnd_net_),
            .in3(N__18754),
            .lcout(n5066),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_1_19_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_LC_1_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_LC_1_19_5  (
            .in0(N__16810),
            .in1(N__18978),
            .in2(N__20476),
            .in3(N__21076),
            .lcout(n7_adj_1998),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_2_lut_LC_1_21_0 .C_ON=1'b1;
    defparam \c0.tx.add_59_2_lut_LC_1_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_2_lut_LC_1_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_2_lut_LC_1_21_0  (
            .in0(_gnd_net_),
            .in1(N__12672),
            .in2(_gnd_net_),
            .in3(N__12118),
            .lcout(\c0.tx.n321 ),
            .ltout(),
            .carryin(bfn_1_21_0_),
            .carryout(\c0.tx.n4414 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_3_lut_LC_1_21_1 .C_ON=1'b1;
    defparam \c0.tx.add_59_3_lut_LC_1_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_3_lut_LC_1_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_3_lut_LC_1_21_1  (
            .in0(_gnd_net_),
            .in1(N__12590),
            .in2(_gnd_net_),
            .in3(N__12115),
            .lcout(\c0.tx.n320 ),
            .ltout(),
            .carryin(\c0.tx.n4414 ),
            .carryout(\c0.tx.n4415 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_4_lut_LC_1_21_2 .C_ON=1'b1;
    defparam \c0.tx.add_59_4_lut_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_4_lut_LC_1_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_4_lut_LC_1_21_2  (
            .in0(_gnd_net_),
            .in1(N__12630),
            .in2(_gnd_net_),
            .in3(N__12112),
            .lcout(n319),
            .ltout(),
            .carryin(\c0.tx.n4415 ),
            .carryout(\c0.tx.n4416 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_5_lut_LC_1_21_3 .C_ON=1'b1;
    defparam \c0.tx.add_59_5_lut_LC_1_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_5_lut_LC_1_21_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_5_lut_LC_1_21_3  (
            .in0(N__13984),
            .in1(N__12511),
            .in2(_gnd_net_),
            .in3(N__12109),
            .lcout(\c0.tx.n5520 ),
            .ltout(),
            .carryin(\c0.tx.n4416 ),
            .carryout(\c0.tx.n4417 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_6_lut_LC_1_21_4 .C_ON=1'b1;
    defparam \c0.tx.add_59_6_lut_LC_1_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_6_lut_LC_1_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_6_lut_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(N__12556),
            .in2(_gnd_net_),
            .in3(N__12106),
            .lcout(n317),
            .ltout(),
            .carryin(\c0.tx.n4417 ),
            .carryout(\c0.tx.n4418 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_7_lut_LC_1_21_5 .C_ON=1'b1;
    defparam \c0.tx.add_59_7_lut_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_7_lut_LC_1_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_7_lut_LC_1_21_5  (
            .in0(_gnd_net_),
            .in1(N__12571),
            .in2(_gnd_net_),
            .in3(N__12103),
            .lcout(n316),
            .ltout(),
            .carryin(\c0.tx.n4418 ),
            .carryout(\c0.tx.n4419 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_8_lut_LC_1_21_6 .C_ON=1'b1;
    defparam \c0.tx.add_59_8_lut_LC_1_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_8_lut_LC_1_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_8_lut_LC_1_21_6  (
            .in0(_gnd_net_),
            .in1(N__12612),
            .in2(_gnd_net_),
            .in3(N__12100),
            .lcout(\c0.tx.n315 ),
            .ltout(),
            .carryin(\c0.tx.n4419 ),
            .carryout(\c0.tx.n4420 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_9_lut_LC_1_21_7 .C_ON=1'b1;
    defparam \c0.tx.add_59_9_lut_LC_1_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_9_lut_LC_1_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_9_lut_LC_1_21_7  (
            .in0(_gnd_net_),
            .in1(N__12538),
            .in2(_gnd_net_),
            .in3(N__12136),
            .lcout(n314),
            .ltout(),
            .carryin(\c0.tx.n4420 ),
            .carryout(\c0.tx.n4421 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_10_lut_LC_1_22_0 .C_ON=1'b0;
    defparam \c0.tx.add_59_10_lut_LC_1_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_10_lut_LC_1_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_10_lut_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(N__14026),
            .in2(_gnd_net_),
            .in3(N__12133),
            .lcout(\c0.tx.n313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_1010_LC_1_22_4.C_ON=1'b0;
    defparam i1_4_lut_adj_1010_LC_1_22_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_1010_LC_1_22_4.LUT_INIT=16'b0000000000110010;
    LogicCell40 i1_4_lut_adj_1010_LC_1_22_4 (
            .in0(N__13856),
            .in1(N__12755),
            .in2(N__14390),
            .in3(N__12127),
            .lcout(n5037),
            .ltout(n5037_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_22_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_22_5 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i8_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(N__12727),
            .in2(N__12130),
            .in3(N__14236),
            .lcout(r_Clock_Count_8_adj_2012),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35283),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i3366_2_lut_LC_1_22_7 .C_ON=1'b0;
    defparam \c0.tx2.i3366_2_lut_LC_1_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i3366_2_lut_LC_1_22_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx2.i3366_2_lut_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(N__14235),
            .in2(_gnd_net_),
            .in3(N__12715),
            .lcout(n3611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_2_lut_3_lut_LC_1_23_0 .C_ON=1'b0;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_1_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_1_23_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx2.i2_2_lut_3_lut_LC_1_23_0  (
            .in0(N__15537),
            .in1(N__15598),
            .in2(_gnd_net_),
            .in3(N__15631),
            .lcout(\c0.tx2.n3577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5286_3_lut_4_lut_4_lut_LC_1_23_1 .C_ON=1'b0;
    defparam \c0.tx2.i5286_3_lut_4_lut_4_lut_LC_1_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5286_3_lut_4_lut_4_lut_LC_1_23_1 .LUT_INIT=16'b1001100000010000;
    LogicCell40 \c0.tx2.i5286_3_lut_4_lut_4_lut_LC_1_23_1  (
            .in0(N__13851),
            .in1(N__14385),
            .in2(N__15793),
            .in3(N__13803),
            .lcout(),
            .ltout(n4_adj_2008_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_47_LC_1_23_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_47_LC_1_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_47_LC_1_23_2 .LUT_INIT=16'b1100110001011100;
    LogicCell40 \c0.tx2.r_Tx_Active_47_LC_1_23_2  (
            .in0(N__14387),
            .in1(N__15749),
            .in2(N__12121),
            .in3(N__14239),
            .lcout(tx2_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35289),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i0_LC_1_23_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i0_LC_1_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i0_LC_1_23_5 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \c0.tx2.r_Clock_Count__i0_LC_1_23_5  (
            .in0(N__14238),
            .in1(_gnd_net_),
            .in2(N__12688),
            .in3(N__14083),
            .lcout(\c0.tx2.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35289),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4968_3_lut_4_lut_LC_1_23_6 .C_ON=1'b0;
    defparam \c0.tx2.i4968_3_lut_4_lut_LC_1_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4968_3_lut_4_lut_LC_1_23_6 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \c0.tx2.i4968_3_lut_4_lut_LC_1_23_6  (
            .in0(N__13804),
            .in1(N__13850),
            .in2(N__14397),
            .in3(N__14237),
            .lcout(),
            .ltout(\c0.tx2.n5312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i0_LC_1_23_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i0_LC_1_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i0_LC_1_23_7 .LUT_INIT=16'b1010000010100100;
    LogicCell40 \c0.tx2.r_Bit_Index_i0_LC_1_23_7  (
            .in0(N__15632),
            .in1(N__14386),
            .in2(N__12157),
            .in3(N__14318),
            .lcout(\c0.tx2.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35289),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i0_LC_1_24_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i0_LC_1_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i0_LC_1_24_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i0_LC_1_24_2  (
            .in0(N__14525),
            .in1(N__13045),
            .in2(N__12151),
            .in3(N__21532),
            .lcout(\c0.tx2.r_Tx_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35295),
            .ce(N__12982),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5450_LC_1_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5450_LC_1_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5450_LC_1_25_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5450_LC_1_25_0  (
            .in0(N__32524),
            .in1(N__16015),
            .in2(N__12295),
            .in3(N__33221),
            .lcout(),
            .ltout(\c0.n5815_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5815_bdd_4_lut_LC_1_25_1 .C_ON=1'b0;
    defparam \c0.n5815_bdd_4_lut_LC_1_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5815_bdd_4_lut_LC_1_25_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n5815_bdd_4_lut_LC_1_25_1  (
            .in0(N__29539),
            .in1(N__32525),
            .in2(N__12154),
            .in3(N__32026),
            .lcout(\c0.n5818 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5659_bdd_4_lut_LC_1_25_2 .C_ON=1'b0;
    defparam \c0.n5659_bdd_4_lut_LC_1_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.n5659_bdd_4_lut_LC_1_25_2 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n5659_bdd_4_lut_LC_1_25_2  (
            .in0(N__22060),
            .in1(N__34807),
            .in2(N__14443),
            .in3(N__12943),
            .lcout(\c0.n5662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n5929_bdd_4_lut_LC_1_25_3 .C_ON=1'b0;
    defparam \c0.tx2.n5929_bdd_4_lut_LC_1_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n5929_bdd_4_lut_LC_1_25_3 .LUT_INIT=16'b1111101000001100;
    LogicCell40 \c0.tx2.n5929_bdd_4_lut_LC_1_25_3  (
            .in0(N__12190),
            .in1(N__12898),
            .in2(N__15604),
            .in3(N__12202),
            .lcout(),
            .ltout(\c0.tx2.n5932_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i341524_i1_3_lut_LC_1_25_4 .C_ON=1'b0;
    defparam \c0.tx2.i341524_i1_3_lut_LC_1_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i341524_i1_3_lut_LC_1_25_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx2.i341524_i1_3_lut_LC_1_25_4  (
            .in0(_gnd_net_),
            .in1(N__15538),
            .in2(N__12142),
            .in3(N__12910),
            .lcout(\c0.tx2.o_Tx_Serial_N_1798 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5543_LC_1_26_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5543_LC_1_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5543_LC_1_26_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5543_LC_1_26_0  (
            .in0(N__14665),
            .in1(N__32522),
            .in2(N__14431),
            .in3(N__33222),
            .lcout(),
            .ltout(\c0.n5917_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5917_bdd_4_lut_LC_1_26_1 .C_ON=1'b0;
    defparam \c0.n5917_bdd_4_lut_LC_1_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5917_bdd_4_lut_LC_1_26_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5917_bdd_4_lut_LC_1_26_1  (
            .in0(N__32523),
            .in1(N__22627),
            .in2(N__12139),
            .in3(N__25677),
            .lcout(),
            .ltout(\c0.n5920_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i7_LC_1_26_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i7_LC_1_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i7_LC_1_26_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i7_LC_1_26_2  (
            .in0(N__14532),
            .in1(N__13060),
            .in2(N__12220),
            .in3(N__12217),
            .lcout(\c0.tx2.r_Tx_Data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35305),
            .ce(N__12992),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_5553_LC_1_26_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_5553_LC_1_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_5553_LC_1_26_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_5553_LC_1_26_3  (
            .in0(N__12196),
            .in1(N__15603),
            .in2(N__12211),
            .in3(N__15633),
            .lcout(\c0.tx2.n5929 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i6_LC_1_26_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i6_LC_1_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i6_LC_1_26_4 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx2.r_Tx_Data_i6_LC_1_26_4  (
            .in0(N__14531),
            .in1(N__34696),
            .in2(N__12937),
            .in3(N__13059),
            .lcout(\c0.tx2.r_Tx_Data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35305),
            .ce(N__12992),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i5_LC_1_26_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i5_LC_1_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i5_LC_1_26_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i5_LC_1_26_6  (
            .in0(N__14530),
            .in1(N__13058),
            .in2(N__14572),
            .in3(N__12175),
            .lcout(\c0.tx2.r_Tx_Data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35305),
            .ce(N__12992),
            .sr(_gnd_net_));
    defparam \c0.n5869_bdd_4_lut_LC_1_27_3 .C_ON=1'b0;
    defparam \c0.n5869_bdd_4_lut_LC_1_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5869_bdd_4_lut_LC_1_27_3 .LUT_INIT=16'b1010110110101000;
    LogicCell40 \c0.n5869_bdd_4_lut_LC_1_27_3  (
            .in0(N__13114),
            .in1(N__25459),
            .in2(N__32588),
            .in3(N__21631),
            .lcout(),
            .ltout(\c0.n5399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5505_LC_1_27_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5505_LC_1_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5505_LC_1_27_4 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5505_LC_1_27_4  (
            .in0(N__34821),
            .in1(N__32115),
            .in2(N__12181),
            .in3(N__12250),
            .lcout(),
            .ltout(\c0.n5857_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5857_bdd_4_lut_LC_1_27_5 .C_ON=1'b0;
    defparam \c0.n5857_bdd_4_lut_LC_1_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.n5857_bdd_4_lut_LC_1_27_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5857_bdd_4_lut_LC_1_27_5  (
            .in0(N__34806),
            .in1(N__25219),
            .in2(N__12178),
            .in3(N__21682),
            .lcout(\c0.n5860 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_1_27_6 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_1_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_1_27_6 .LUT_INIT=16'b1011101110011001;
    LogicCell40 \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_1_27_6  (
            .in0(N__14398),
            .in1(N__13861),
            .in2(_gnd_net_),
            .in3(N__12169),
            .lcout(),
            .ltout(n3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_45_LC_1_27_7 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_45_LC_1_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.o_Tx_Serial_45_LC_1_27_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.tx2.o_Tx_Serial_45_LC_1_27_7  (
            .in0(N__14253),
            .in1(_gnd_net_),
            .in2(N__12160),
            .in3(N__12277),
            .lcout(tx2_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35309),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i153_LC_1_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i153_LC_1_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i153_LC_1_28_2 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0___i153_LC_1_28_2  (
            .in0(N__36175),
            .in1(N__12291),
            .in2(N__37268),
            .in3(N__21462),
            .lcout(\c0.data_in_frame_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_28_3 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_28_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_1_28_3  (
            .in0(N__12275),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx2_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5863_bdd_4_lut_LC_1_28_5 .C_ON=1'b0;
    defparam \c0.n5863_bdd_4_lut_LC_1_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.n5863_bdd_4_lut_LC_1_28_5 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n5863_bdd_4_lut_LC_1_28_5  (
            .in0(N__12229),
            .in1(N__17566),
            .in2(N__15967),
            .in3(N__32518),
            .lcout(\c0.n5402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i34_LC_1_29_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i34_LC_1_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i34_LC_1_29_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i34_LC_1_29_0  (
            .in0(N__29324),
            .in1(N__13422),
            .in2(_gnd_net_),
            .in3(N__34147),
            .lcout(data_in_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i156_LC_1_29_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i156_LC_1_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i156_LC_1_29_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i156_LC_1_29_2  (
            .in0(N__12243),
            .in1(N__15857),
            .in2(N__37228),
            .in3(N__36289),
            .lcout(\c0.data_in_frame_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5568_LC_1_29_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5568_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5568_LC_1_29_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5568_LC_1_29_3  (
            .in0(N__13084),
            .in1(N__32586),
            .in2(N__12244),
            .in3(N__33273),
            .lcout(\c0.n5959 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5490_LC_1_29_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5490_LC_1_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5490_LC_1_29_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5490_LC_1_29_4  (
            .in0(N__33272),
            .in1(N__23068),
            .in2(N__32629),
            .in3(N__28809),
            .lcout(\c0.n5863 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_1_29_5 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_1_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_1_29_5 .LUT_INIT=16'b0011010000110000;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_1_29_5  (
            .in0(N__13513),
            .in1(N__13180),
            .in2(N__18177),
            .in3(N__18283),
            .lcout(\c0.rx.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_2_lut_LC_1_30_0 .C_ON=1'b1;
    defparam \c0.rx.add_62_2_lut_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_2_lut_LC_1_30_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_2_lut_LC_1_30_0  (
            .in0(N__12301),
            .in1(N__14911),
            .in2(_gnd_net_),
            .in3(N__12223),
            .lcout(n5491),
            .ltout(),
            .carryin(bfn_1_30_0_),
            .carryout(\c0.rx.n4422 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_3_lut_LC_1_30_1 .C_ON=1'b1;
    defparam \c0.rx.add_62_3_lut_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_3_lut_LC_1_30_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_3_lut_LC_1_30_1  (
            .in0(N__13448),
            .in1(N__13345),
            .in2(_gnd_net_),
            .in3(N__12325),
            .lcout(\c0.rx.n5537 ),
            .ltout(),
            .carryin(\c0.rx.n4422 ),
            .carryout(\c0.rx.n4423 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_4_lut_LC_1_30_2 .C_ON=1'b1;
    defparam \c0.rx.add_62_4_lut_LC_1_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_4_lut_LC_1_30_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_4_lut_LC_1_30_2  (
            .in0(N__13440),
            .in1(N__14730),
            .in2(_gnd_net_),
            .in3(N__12322),
            .lcout(\c0.rx.n5536 ),
            .ltout(),
            .carryin(\c0.rx.n4423 ),
            .carryout(\c0.rx.n4424 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_5_lut_LC_1_30_3 .C_ON=1'b1;
    defparam \c0.rx.add_62_5_lut_LC_1_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_5_lut_LC_1_30_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_5_lut_LC_1_30_3  (
            .in0(N__13449),
            .in1(N__13308),
            .in2(_gnd_net_),
            .in3(N__12319),
            .lcout(\c0.rx.n5539 ),
            .ltout(),
            .carryin(\c0.rx.n4424 ),
            .carryout(\c0.rx.n4425 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_6_lut_LC_1_30_4 .C_ON=1'b1;
    defparam \c0.rx.add_62_6_lut_LC_1_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_6_lut_LC_1_30_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_6_lut_LC_1_30_4  (
            .in0(N__13439),
            .in1(N__13374),
            .in2(_gnd_net_),
            .in3(N__12316),
            .lcout(\c0.rx.n5535 ),
            .ltout(),
            .carryin(\c0.rx.n4425 ),
            .carryout(\c0.rx.n4426 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_7_lut_LC_1_30_5 .C_ON=1'b1;
    defparam \c0.rx.add_62_7_lut_LC_1_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_7_lut_LC_1_30_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_7_lut_LC_1_30_5  (
            .in0(N__13450),
            .in1(N__13398),
            .in2(_gnd_net_),
            .in3(N__12313),
            .lcout(\c0.rx.n5538 ),
            .ltout(),
            .carryin(\c0.rx.n4426 ),
            .carryout(\c0.rx.n4427 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_8_lut_LC_1_30_6 .C_ON=1'b1;
    defparam \c0.rx.add_62_8_lut_LC_1_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_8_lut_LC_1_30_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_8_lut_LC_1_30_6  (
            .in0(N__12355),
            .in1(N__14881),
            .in2(_gnd_net_),
            .in3(N__12310),
            .lcout(n5051),
            .ltout(),
            .carryin(\c0.rx.n4427 ),
            .carryout(\c0.rx.n4428 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_9_lut_LC_1_30_7 .C_ON=1'b0;
    defparam \c0.rx.add_62_9_lut_LC_1_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_9_lut_LC_1_30_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.rx.add_62_9_lut_LC_1_30_7  (
            .in0(_gnd_net_),
            .in1(N__12354),
            .in2(N__14767),
            .in3(N__12307),
            .lcout(n5050),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i59_3_lut_LC_1_31_0 .C_ON=1'b0;
    defparam \c0.rx.i59_3_lut_LC_1_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i59_3_lut_LC_1_31_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \c0.rx.i59_3_lut_LC_1_31_0  (
            .in0(N__14724),
            .in1(N__13338),
            .in2(_gnd_net_),
            .in3(N__13305),
            .lcout(\c0.rx.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_791_LC_1_31_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_791_LC_1_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_791_LC_1_31_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.rx.i1_2_lut_adj_791_LC_1_31_1  (
            .in0(N__18109),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18269),
            .lcout(n2156),
            .ltout(n2156_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4941_1_lut_4_lut_LC_1_31_2.C_ON=1'b0;
    defparam i4941_1_lut_4_lut_LC_1_31_2.SEQ_MODE=4'b0000;
    defparam i4941_1_lut_4_lut_LC_1_31_2.LUT_INIT=16'b0000010011111111;
    LogicCell40 i4941_1_lut_4_lut_LC_1_31_2 (
            .in0(N__18330),
            .in1(N__13282),
            .in2(N__12304),
            .in3(N__13153),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4954_2_lut_LC_1_31_3 .C_ON=1'b0;
    defparam \c0.rx.i4954_2_lut_LC_1_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4954_2_lut_LC_1_31_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i4954_2_lut_LC_1_31_3  (
            .in0(_gnd_net_),
            .in1(N__14760),
            .in2(_gnd_net_),
            .in3(N__13397),
            .lcout(),
            .ltout(\c0.rx.n5298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4972_4_lut_LC_1_31_4 .C_ON=1'b0;
    defparam \c0.rx.i4972_4_lut_LC_1_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4972_4_lut_LC_1_31_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.rx.i4972_4_lut_LC_1_31_4  (
            .in0(N__13339),
            .in1(N__13306),
            .in2(N__12364),
            .in3(N__13373),
            .lcout(n5316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i2_LC_1_31_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i2_LC_1_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_1_31_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_1_31_5  (
            .in0(N__13224),
            .in1(N__14725),
            .in2(_gnd_net_),
            .in3(N__12361),
            .lcout(\c0.rx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_4_lut_LC_1_31_6 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_4_lut_LC_1_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_4_lut_LC_1_31_6 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \c0.rx.i2_4_lut_4_lut_LC_1_31_6  (
            .in0(N__12379),
            .in1(N__18046),
            .in2(N__18282),
            .in3(N__13223),
            .lcout(\c0.rx.n5049 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i7_LC_1_31_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_1_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_1_31_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_1_31_7  (
            .in0(N__13225),
            .in1(N__14761),
            .in2(_gnd_net_),
            .in3(N__12346),
            .lcout(r_Clock_Count_7_adj_2004),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_4_lut_LC_1_32_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_4_lut_LC_1_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_4_lut_LC_1_32_0 .LUT_INIT=16'b0110001010101010;
    LogicCell40 \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_4_lut_LC_1_32_0  (
            .in0(N__18130),
            .in1(N__18266),
            .in2(N__13509),
            .in3(N__18047),
            .lcout(),
            .ltout(\c0.rx.n5923_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.n5923_bdd_4_lut_4_lut_LC_1_32_1 .C_ON=1'b0;
    defparam \c0.rx.n5923_bdd_4_lut_4_lut_LC_1_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.n5923_bdd_4_lut_4_lut_LC_1_32_1 .LUT_INIT=16'b1110000011100011;
    LogicCell40 \c0.rx.n5923_bdd_4_lut_4_lut_LC_1_32_1  (
            .in0(N__13280),
            .in1(N__18267),
            .in2(N__12340),
            .in3(N__20899),
            .lcout(),
            .ltout(\c0.rx.n5926_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_1_32_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_1_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_1_32_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_1_32_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12337),
            .in3(N__18363),
            .lcout(r_SM_Main_0_adj_2006),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i1_LC_1_32_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i1_LC_1_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_1_32_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_1_32_3  (
            .in0(N__13238),
            .in1(N__13344),
            .in2(_gnd_net_),
            .in3(N__12334),
            .lcout(\c0.rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(_gnd_net_));
    defparam i5253_2_lut_LC_1_32_4.C_ON=1'b0;
    defparam i5253_2_lut_LC_1_32_4.SEQ_MODE=4'b0000;
    defparam i5253_2_lut_LC_1_32_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 i5253_2_lut_LC_1_32_4 (
            .in0(_gnd_net_),
            .in1(N__18112),
            .in2(_gnd_net_),
            .in3(N__13278),
            .lcout(n5490),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5269_3_lut_LC_1_32_5 .C_ON=1'b0;
    defparam \c0.rx.i5269_3_lut_LC_1_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5269_3_lut_LC_1_32_5 .LUT_INIT=16'b1111111110101111;
    LogicCell40 \c0.rx.i5269_3_lut_LC_1_32_5  (
            .in0(N__13279),
            .in1(_gnd_net_),
            .in2(N__18131),
            .in3(N__20898),
            .lcout(\c0.rx.n5532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_795_LC_1_32_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_795_LC_1_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_795_LC_1_32_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_795_LC_1_32_6  (
            .in0(_gnd_net_),
            .in1(N__18116),
            .in2(_gnd_net_),
            .in3(N__18048),
            .lcout(),
            .ltout(\c0.rx.n3980_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_1_32_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_1_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_1_32_7 .LUT_INIT=16'b0000010000010101;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_1_32_7  (
            .in0(N__18362),
            .in1(N__18268),
            .in2(N__12373),
            .in3(N__12370),
            .lcout(\c0.rx.r_SM_Main_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i2_LC_2_16_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i2_LC_2_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i2_LC_2_16_0 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \c0.byte_transmit_counter__i2_LC_2_16_0  (
            .in0(N__13580),
            .in1(N__13542),
            .in2(N__13485),
            .in3(N__12433),
            .lcout(\c0.byte_transmit_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35271),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i7_LC_2_16_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i7_LC_2_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i7_LC_2_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter__i7_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__13478),
            .in2(_gnd_net_),
            .in3(N__13594),
            .lcout(\c0.byte_transmit_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35271),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_908_LC_2_16_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_908_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_908_LC_2_16_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_908_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__12432),
            .in2(_gnd_net_),
            .in3(N__12420),
            .lcout(\c0.n103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_968_LC_2_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_968_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_968_LC_2_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_968_LC_2_16_3  (
            .in0(N__20610),
            .in1(N__20718),
            .in2(_gnd_net_),
            .in3(N__16431),
            .lcout(n1525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i5_LC_2_16_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i5_LC_2_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i5_LC_2_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter__i5_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(N__13476),
            .in2(_gnd_net_),
            .in3(N__13618),
            .lcout(\c0.byte_transmit_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35271),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i3_LC_2_16_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i3_LC_2_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i3_LC_2_16_6 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \c0.byte_transmit_counter__i3_LC_2_16_6  (
            .in0(N__13581),
            .in1(N__13543),
            .in2(N__13486),
            .in3(N__12421),
            .lcout(\c0.byte_transmit_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35271),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i6_LC_2_16_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i6_LC_2_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i6_LC_2_16_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter__i6_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(N__13477),
            .in2(_gnd_net_),
            .in3(N__13606),
            .lcout(\c0.byte_transmit_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35271),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i0_LC_2_17_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter__i0_LC_2_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i0_LC_2_17_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \c0.byte_transmit_counter__i0_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__12457),
            .in2(N__20354),
            .in3(N__16663),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\c0.n4378 ),
            .clk(N__35269),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i1_LC_2_17_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter__i1_LC_2_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i1_LC_2_17_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.byte_transmit_counter__i1_LC_2_17_1  (
            .in0(N__16664),
            .in1(N__20508),
            .in2(_gnd_net_),
            .in3(N__12436),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(\c0.n4378 ),
            .carryout(\c0.n4379 ),
            .clk(N__35269),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_4_lut_LC_2_17_2 .C_ON=1'b1;
    defparam \c0.add_1824_4_lut_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_4_lut_LC_2_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_4_lut_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__21261),
            .in2(_gnd_net_),
            .in3(N__12424),
            .lcout(\c0.tx_transmit_N_568_2 ),
            .ltout(),
            .carryin(\c0.n4379 ),
            .carryout(\c0.n4380 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_5_lut_LC_2_17_3 .C_ON=1'b1;
    defparam \c0.add_1824_5_lut_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_5_lut_LC_2_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_5_lut_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__21345),
            .in2(_gnd_net_),
            .in3(N__12412),
            .lcout(\c0.tx_transmit_N_568_3 ),
            .ltout(),
            .carryin(\c0.n4380 ),
            .carryout(\c0.n4381 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_6_lut_LC_2_17_4 .C_ON=1'b1;
    defparam \c0.add_1824_6_lut_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_6_lut_LC_2_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_6_lut_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__21148),
            .in2(_gnd_net_),
            .in3(N__12409),
            .lcout(\c0.tx_transmit_N_568_4 ),
            .ltout(),
            .carryin(\c0.n4381 ),
            .carryout(\c0.n4382 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_7_lut_LC_2_17_5 .C_ON=1'b1;
    defparam \c0.add_1824_7_lut_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_7_lut_LC_2_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_7_lut_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__12406),
            .in2(_gnd_net_),
            .in3(N__12400),
            .lcout(\c0.tx_transmit_N_568_5 ),
            .ltout(),
            .carryin(\c0.n4382 ),
            .carryout(\c0.n4383 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_8_lut_LC_2_17_6 .C_ON=1'b1;
    defparam \c0.add_1824_8_lut_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_8_lut_LC_2_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_8_lut_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__12397),
            .in2(_gnd_net_),
            .in3(N__12391),
            .lcout(\c0.tx_transmit_N_568_6 ),
            .ltout(),
            .carryin(\c0.n4383 ),
            .carryout(\c0.n4384 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_9_lut_LC_2_17_7 .C_ON=1'b0;
    defparam \c0.add_1824_9_lut_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_9_lut_LC_2_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_9_lut_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__12388),
            .in2(_gnd_net_),
            .in3(N__12382),
            .lcout(\c0.tx_transmit_N_568_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i23_LC_2_18_1 .C_ON=1'b0;
    defparam \c0.data_out_0___i23_LC_2_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i23_LC_2_18_1 .LUT_INIT=16'b1010101011000011;
    LogicCell40 \c0.data_out_0___i23_LC_2_18_1  (
            .in0(N__20763),
            .in1(N__13671),
            .in2(N__16291),
            .in3(N__16672),
            .lcout(data_out_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35272),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_985_LC_2_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_985_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_985_LC_2_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_985_LC_2_18_2  (
            .in0(N__18967),
            .in1(N__18735),
            .in2(_gnd_net_),
            .in3(N__19297),
            .lcout(n5077),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_959_LC_2_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_959_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_959_LC_2_18_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i1_2_lut_adj_959_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__12451),
            .in2(_gnd_net_),
            .in3(N__13641),
            .lcout(\c0.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_prev_1793_LC_2_18_4 .C_ON=1'b0;
    defparam \c0.tx_active_prev_1793_LC_2_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx_active_prev_1793_LC_2_18_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.tx_active_prev_1793_LC_2_18_4  (
            .in0(N__13642),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.tx_active_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35272),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5277_4_lut_LC_2_18_5 .C_ON=1'b0;
    defparam \c0.i5277_4_lut_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5277_4_lut_LC_2_18_5 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.i5277_4_lut_LC_2_18_5  (
            .in0(N__21006),
            .in1(N__20324),
            .in2(N__16566),
            .in3(N__20509),
            .lcout(),
            .ltout(\c0.n5540_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_2_18_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_2_18_6 .LUT_INIT=16'b0111011111000000;
    LogicCell40 \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_2_18_6  (
            .in0(N__20510),
            .in1(N__21379),
            .in2(N__12445),
            .in3(N__21288),
            .lcout(),
            .ltout(\c0.n5977_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5977_bdd_4_lut_4_lut_LC_2_18_7 .C_ON=1'b0;
    defparam \c0.n5977_bdd_4_lut_4_lut_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.n5977_bdd_4_lut_4_lut_LC_2_18_7 .LUT_INIT=16'b1111000110100101;
    LogicCell40 \c0.n5977_bdd_4_lut_4_lut_LC_2_18_7  (
            .in0(N__21380),
            .in1(N__20325),
            .in2(N__12442),
            .in3(N__20511),
            .lcout(\c0.n5980 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_843_LC_2_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_843_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_843_LC_2_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_843_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__21075),
            .in2(_gnd_net_),
            .in3(N__21007),
            .lcout(n1760),
            .ltout(n1760_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i18_LC_2_19_1 .C_ON=1'b0;
    defparam \c0.data_out_0___i18_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i18_LC_2_19_1 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \c0.data_out_0___i18_LC_2_19_1  (
            .in0(N__15288),
            .in1(N__16444),
            .in2(N__12439),
            .in3(N__16677),
            .lcout(data_out_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35274),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_2_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_2_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_2_19_2  (
            .in0(N__19283),
            .in1(N__16284),
            .in2(_gnd_net_),
            .in3(N__20392),
            .lcout(\c0.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_935_LC_2_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_935_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_935_LC_2_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_935_LC_2_19_3  (
            .in0(N__16570),
            .in1(N__18805),
            .in2(_gnd_net_),
            .in3(N__15155),
            .lcout(),
            .ltout(\c0.n1529_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_835_LC_2_19_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_835_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_835_LC_2_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_835_LC_2_19_4  (
            .in0(N__15021),
            .in1(N__12496),
            .in2(N__12490),
            .in3(N__12487),
            .lcout(n5079),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_2_19_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_2_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_2_19_6  (
            .in0(N__20470),
            .in1(N__18979),
            .in2(_gnd_net_),
            .in3(N__21008),
            .lcout(n7_adj_2002),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_874_LC_2_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_874_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_874_LC_2_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_874_LC_2_19_7  (
            .in0(_gnd_net_),
            .in1(N__16283),
            .in2(_gnd_net_),
            .in3(N__16371),
            .lcout(\c0.n1801 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i6_LC_2_20_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i6_LC_2_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_2_20_1 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_2_20_1  (
            .in0(N__12481),
            .in1(N__13978),
            .in2(N__16999),
            .in3(N__12613),
            .lcout(\c0.tx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35278),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_2_20_2 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_2_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_2_20_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_2_20_2  (
            .in0(N__19342),
            .in1(N__15264),
            .in2(_gnd_net_),
            .in3(N__15415),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35278),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i2_LC_2_20_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i2_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_2_20_3 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_2_20_3  (
            .in0(N__16979),
            .in1(N__13977),
            .in2(N__12634),
            .in3(N__12475),
            .lcout(r_Clock_Count_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35278),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i1_LC_2_20_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i1_LC_2_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_2_20_4 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_2_20_4  (
            .in0(N__13976),
            .in1(N__16978),
            .in2(N__12595),
            .in3(N__12469),
            .lcout(\c0.tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35278),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_2_20_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i0_LC_2_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_2_20_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_2_20_7  (
            .in0(N__16977),
            .in1(N__12463),
            .in2(N__12676),
            .in3(N__13979),
            .lcout(\c0.tx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35278),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i8_LC_2_21_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_2_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_2_21_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_2_21_0  (
            .in0(N__12661),
            .in1(N__14025),
            .in2(N__17001),
            .in3(N__13983),
            .lcout(r_Clock_Count_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35284),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i5_LC_2_21_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i5_LC_2_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_2_21_1 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_2_21_1  (
            .in0(N__12570),
            .in1(N__12655),
            .in2(N__16998),
            .in3(N__13981),
            .lcout(r_Clock_Count_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35284),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i7_LC_2_21_2 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i7_LC_2_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_2_21_2 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_2_21_2  (
            .in0(N__12537),
            .in1(N__12649),
            .in2(N__17000),
            .in3(N__13982),
            .lcout(r_Clock_Count_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35284),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i4_LC_2_21_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i4_LC_2_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_2_21_3 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_2_21_3  (
            .in0(N__16973),
            .in1(N__13980),
            .in2(N__12643),
            .in3(N__12555),
            .lcout(r_Clock_Count_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35284),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_adj_805_LC_2_21_4 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_adj_805_LC_2_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_adj_805_LC_2_21_4 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \c0.tx.i1_4_lut_adj_805_LC_2_21_4  (
            .in0(N__12629),
            .in1(N__12611),
            .in2(N__12594),
            .in3(N__12509),
            .lcout(),
            .ltout(\c0.tx.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i3351_4_lut_LC_2_21_5 .C_ON=1'b0;
    defparam \c0.tx.i3351_4_lut_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i3351_4_lut_LC_2_21_5 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.tx.i3351_4_lut_LC_2_21_5  (
            .in0(N__12569),
            .in1(N__12554),
            .in2(N__12541),
            .in3(N__12536),
            .lcout(n3595),
            .ltout(n3595_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_2_21_6.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_2_21_6.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_2_21_6.LUT_INIT=16'b0100010001000000;
    LogicCell40 i2_3_lut_4_lut_LC_2_21_6 (
            .in0(N__16984),
            .in1(N__17051),
            .in2(N__12523),
            .in3(N__14024),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i3_LC_2_21_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i3_LC_2_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_2_21_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_2_21_7  (
            .in0(N__12510),
            .in1(_gnd_net_),
            .in2(N__12520),
            .in3(N__16985),
            .lcout(\c0.tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35284),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_LC_2_22_0 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_LC_2_22_0 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \c0.tx2.i1_4_lut_LC_2_22_0  (
            .in0(N__13877),
            .in1(N__12788),
            .in2(N__12886),
            .in3(N__14054),
            .lcout(),
            .ltout(\c0.tx2.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i3348_4_lut_LC_2_22_1 .C_ON=1'b0;
    defparam \c0.tx2.i3348_4_lut_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i3348_4_lut_LC_2_22_1 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \c0.tx2.i3348_4_lut_LC_2_22_1  (
            .in0(N__12818),
            .in1(N__12848),
            .in2(N__12718),
            .in3(N__13901),
            .lcout(\c0.tx2.n3591 ),
            .ltout(\c0.tx2.n3591_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i3380_2_lut_LC_2_22_2 .C_ON=1'b0;
    defparam \c0.tx2.i3380_2_lut_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i3380_2_lut_LC_2_22_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.tx2.i3380_2_lut_LC_2_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12709),
            .in3(N__12748),
            .lcout(r_SM_Main_2_N_1767_1),
            .ltout(r_SM_Main_2_N_1767_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i1_LC_2_22_3 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_22_3 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \c0.tx2.r_SM_Main_i1_LC_2_22_3  (
            .in0(N__14388),
            .in1(N__13860),
            .in2(N__12706),
            .in3(N__14248),
            .lcout(r_SM_Main_1_adj_2010),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i6_LC_2_22_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i6_LC_2_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i6_LC_2_22_4 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i6_LC_2_22_4  (
            .in0(N__14087),
            .in1(_gnd_net_),
            .in2(N__14263),
            .in3(N__12772),
            .lcout(\c0.tx2.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i4_LC_2_22_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i4_LC_2_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i4_LC_2_22_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i4_LC_2_22_5  (
            .in0(N__12832),
            .in1(N__14241),
            .in2(_gnd_net_),
            .in3(N__14085),
            .lcout(\c0.tx2.r_Clock_Count_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i5_LC_2_22_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i5_LC_2_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i5_LC_2_22_6 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i5_LC_2_22_6  (
            .in0(N__14086),
            .in1(_gnd_net_),
            .in2(N__14262),
            .in3(N__12802),
            .lcout(\c0.tx2.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_22_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_22_7 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i1_LC_2_22_7  (
            .in0(N__12865),
            .in1(N__14240),
            .in2(_gnd_net_),
            .in3(N__14084),
            .lcout(\c0.tx2.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_2_lut_LC_2_23_0 .C_ON=1'b1;
    defparam \c0.tx2.add_59_2_lut_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_2_lut_LC_2_23_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_2_lut_LC_2_23_0  (
            .in0(N__12703),
            .in1(N__12702),
            .in2(N__14254),
            .in3(N__12679),
            .lcout(n2460),
            .ltout(),
            .carryin(bfn_2_23_0_),
            .carryout(\c0.tx2.n4429 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_3_lut_LC_2_23_1 .C_ON=1'b1;
    defparam \c0.tx2.add_59_3_lut_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_3_lut_LC_2_23_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_3_lut_LC_2_23_1  (
            .in0(N__12885),
            .in1(N__12884),
            .in2(N__14258),
            .in3(N__12859),
            .lcout(n2399),
            .ltout(),
            .carryin(\c0.tx2.n4429 ),
            .carryout(\c0.tx2.n4430 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_4_lut_LC_2_23_2 .C_ON=1'b1;
    defparam \c0.tx2.add_59_4_lut_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_4_lut_LC_2_23_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_4_lut_LC_2_23_2  (
            .in0(N__13879),
            .in1(N__13878),
            .in2(N__14255),
            .in3(N__12856),
            .lcout(n2395),
            .ltout(),
            .carryin(\c0.tx2.n4430 ),
            .carryout(\c0.tx2.n4431 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_5_lut_LC_2_23_3 .C_ON=1'b1;
    defparam \c0.tx2.add_59_5_lut_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_5_lut_LC_2_23_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_5_lut_LC_2_23_3  (
            .in0(N__14056),
            .in1(N__14055),
            .in2(N__14259),
            .in3(N__12853),
            .lcout(n2392),
            .ltout(),
            .carryin(\c0.tx2.n4431 ),
            .carryout(\c0.tx2.n4432 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_6_lut_LC_2_23_4 .C_ON=1'b1;
    defparam \c0.tx2.add_59_6_lut_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_6_lut_LC_2_23_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_6_lut_LC_2_23_4  (
            .in0(N__12850),
            .in1(N__12849),
            .in2(N__14256),
            .in3(N__12823),
            .lcout(n2382),
            .ltout(),
            .carryin(\c0.tx2.n4432 ),
            .carryout(\c0.tx2.n4433 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_7_lut_LC_2_23_5 .C_ON=1'b1;
    defparam \c0.tx2.add_59_7_lut_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_7_lut_LC_2_23_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_7_lut_LC_2_23_5  (
            .in0(N__12820),
            .in1(N__12819),
            .in2(N__14260),
            .in3(N__12793),
            .lcout(n2379),
            .ltout(),
            .carryin(\c0.tx2.n4433 ),
            .carryout(\c0.tx2.n4434 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_8_lut_LC_2_23_6 .C_ON=1'b1;
    defparam \c0.tx2.add_59_8_lut_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_8_lut_LC_2_23_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_8_lut_LC_2_23_6  (
            .in0(N__12790),
            .in1(N__12789),
            .in2(N__14257),
            .in3(N__12763),
            .lcout(n2376),
            .ltout(),
            .carryin(\c0.tx2.n4434 ),
            .carryout(\c0.tx2.n4435 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_9_lut_LC_2_23_7 .C_ON=1'b1;
    defparam \c0.tx2.add_59_9_lut_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_9_lut_LC_2_23_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_9_lut_LC_2_23_7  (
            .in0(N__13903),
            .in1(N__13902),
            .in2(N__14261),
            .in3(N__12760),
            .lcout(n2372),
            .ltout(),
            .carryin(\c0.tx2.n4435 ),
            .carryout(\c0.tx2.n4436 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_10_lut_LC_2_24_0 .C_ON=1'b0;
    defparam \c0.tx2.add_59_10_lut_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_10_lut_LC_2_24_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx2.add_59_10_lut_LC_2_24_0  (
            .in0(N__12756),
            .in1(N__12757),
            .in2(N__14252),
            .in3(N__12730),
            .lcout(n2369),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i0_LC_2_24_1 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i0_LC_2_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i0_LC_2_24_1 .LUT_INIT=16'b0000011100000100;
    LogicCell40 \c0.tx2.r_SM_Main_i0_LC_2_24_1  (
            .in0(N__13807),
            .in1(N__13854),
            .in2(N__14250),
            .in3(N__12904),
            .lcout(r_SM_Main_0_adj_2011),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_24_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_24_2 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_24_2  (
            .in0(N__12955),
            .in1(N__12892),
            .in2(N__15602),
            .in3(N__15624),
            .lcout(\c0.tx2.n5947 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n5947_bdd_4_lut_LC_2_24_3 .C_ON=1'b0;
    defparam \c0.tx2.n5947_bdd_4_lut_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n5947_bdd_4_lut_LC_2_24_3 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.tx2.n5947_bdd_4_lut_LC_2_24_3  (
            .in0(N__13003),
            .in1(N__15594),
            .in2(N__12925),
            .in3(N__12916),
            .lcout(\c0.tx2.n5950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1104_4_lut_LC_2_24_4 .C_ON=1'b0;
    defparam \c0.tx2.i1104_4_lut_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1104_4_lut_LC_2_24_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \c0.tx2.i1104_4_lut_LC_2_24_4  (
            .in0(N__14391),
            .in1(N__15783),
            .in2(N__14322),
            .in3(N__13805),
            .lcout(n1345),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_3_lut_4_lut_LC_2_24_5 .C_ON=1'b0;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_2_24_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx2.i2_3_lut_4_lut_LC_2_24_5  (
            .in0(N__15782),
            .in1(N__13852),
            .in2(N__14249),
            .in3(N__14392),
            .lcout(\c0.tx2.n1592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i817_2_lut_LC_2_24_6 .C_ON=1'b0;
    defparam \c0.i817_2_lut_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i817_2_lut_LC_2_24_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i817_2_lut_LC_2_24_6  (
            .in0(_gnd_net_),
            .in1(N__34747),
            .in2(_gnd_net_),
            .in3(N__32079),
            .lcout(\c0.n1058 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i2_LC_2_24_7 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i2_LC_2_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i2_LC_2_24_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.tx2.r_SM_Main_i2_LC_2_24_7  (
            .in0(N__13806),
            .in1(N__13853),
            .in2(N__14251),
            .in3(N__14393),
            .lcout(r_SM_Main_2_adj_2009),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5563_LC_2_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5563_LC_2_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5563_LC_2_25_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5563_LC_2_25_0  (
            .in0(N__15997),
            .in1(N__32316),
            .in2(N__35440),
            .in3(N__33115),
            .lcout(\c0.n5953 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i4_LC_2_25_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i4_LC_2_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i4_LC_2_25_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.tx2.r_Tx_Data_i4_LC_2_25_2  (
            .in0(N__13048),
            .in1(N__14511),
            .in2(N__14284),
            .in3(N__18916),
            .lcout(\c0.tx2.r_Tx_Data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35306),
            .ce(N__12993),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i2_LC_2_25_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i2_LC_2_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i2_LC_2_25_5 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i2_LC_2_25_5  (
            .in0(N__14509),
            .in1(N__13046),
            .in2(N__14452),
            .in3(N__22882),
            .lcout(\c0.tx2.r_Tx_Data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35306),
            .ce(N__12993),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i3_LC_2_25_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i3_LC_2_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i3_LC_2_25_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i3_LC_2_25_7  (
            .in0(N__14510),
            .in1(N__13047),
            .in2(N__13096),
            .in3(N__14458),
            .lcout(\c0.tx2.r_Tx_Data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35306),
            .ce(N__12993),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5326_LC_2_26_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5326_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5326_LC_2_26_0 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5326_LC_2_26_0  (
            .in0(N__17732),
            .in1(N__33287),
            .in2(N__32544),
            .in3(N__27661),
            .lcout(),
            .ltout(\c0.n5665_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5665_bdd_4_lut_LC_2_26_1 .C_ON=1'b0;
    defparam \c0.n5665_bdd_4_lut_LC_2_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5665_bdd_4_lut_LC_2_26_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n5665_bdd_4_lut_LC_2_26_1  (
            .in0(N__25702),
            .in1(N__24756),
            .in2(N__12949),
            .in3(N__32444),
            .lcout(),
            .ltout(\c0.n5372_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5331_LC_2_26_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5331_LC_2_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5331_LC_2_26_2 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5331_LC_2_26_2  (
            .in0(N__32099),
            .in1(N__34805),
            .in2(N__12946),
            .in3(N__13123),
            .lcout(\c0.n5659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5310_4_lut_LC_2_26_3 .C_ON=1'b0;
    defparam \c0.i5310_4_lut_LC_2_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5310_4_lut_LC_2_26_3 .LUT_INIT=16'b0001111100111111;
    LogicCell40 \c0.i5310_4_lut_LC_2_26_3  (
            .in0(N__33288),
            .in1(N__13056),
            .in2(N__14533),
            .in3(N__32443),
            .lcout(\c0.FRAME_MATCHER_wait_for_transmission_N_909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5935_bdd_4_lut_LC_2_26_4 .C_ON=1'b0;
    defparam \c0.n5935_bdd_4_lut_LC_2_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.n5935_bdd_4_lut_LC_2_26_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5935_bdd_4_lut_LC_2_26_4  (
            .in0(N__32445),
            .in1(N__27139),
            .in2(N__14407),
            .in3(N__19681),
            .lcout(\c0.n5938 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i140_LC_2_26_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i140_LC_2_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i140_LC_2_26_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \c0.data_in_0___i140_LC_2_26_6  (
            .in0(N__34362),
            .in1(N__14639),
            .in2(N__17534),
            .in3(_gnd_net_),
            .lcout(data_in_17_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35310),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i148_LC_2_26_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i148_LC_2_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i148_LC_2_26_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.data_in_0___i148_LC_2_26_7  (
            .in0(_gnd_net_),
            .in1(N__15861),
            .in2(N__14646),
            .in3(N__34361),
            .lcout(data_in_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35310),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_27_0 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_27_0  (
            .in0(N__33246),
            .in1(N__13138),
            .in2(N__14593),
            .in3(N__32526),
            .lcout(),
            .ltout(\c0.n5971_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5971_bdd_4_lut_LC_2_27_1 .C_ON=1'b0;
    defparam \c0.n5971_bdd_4_lut_LC_2_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5971_bdd_4_lut_LC_2_27_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5971_bdd_4_lut_LC_2_27_1  (
            .in0(N__32527),
            .in1(N__30872),
            .in2(N__12928),
            .in3(N__19939),
            .lcout(\c0.n5974 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5395_LC_2_27_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5395_LC_2_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5395_LC_2_27_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5395_LC_2_27_2  (
            .in0(N__32108),
            .in1(N__16051),
            .in2(N__34827),
            .in3(N__14608),
            .lcout(),
            .ltout(\c0.n5725_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5725_bdd_4_lut_LC_2_27_3 .C_ON=1'b0;
    defparam \c0.n5725_bdd_4_lut_LC_2_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5725_bdd_4_lut_LC_2_27_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n5725_bdd_4_lut_LC_2_27_3  (
            .in0(N__25822),
            .in1(N__34811),
            .in2(N__13063),
            .in3(N__14542),
            .lcout(),
            .ltout(\c0.n5728_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i1_LC_2_27_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i1_LC_2_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i1_LC_2_27_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.tx2.r_Tx_Data_i1_LC_2_27_4  (
            .in0(N__14526),
            .in1(N__13057),
            .in2(N__13012),
            .in3(N__13009),
            .lcout(\c0.tx2.r_Tx_Data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35314),
            .ce(N__12994),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i132_LC_2_28_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i132_LC_2_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i132_LC_2_28_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i132_LC_2_28_0  (
            .in0(N__26831),
            .in1(N__17535),
            .in2(_gnd_net_),
            .in3(N__34294),
            .lcout(data_in_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i42_LC_2_28_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i42_LC_2_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i42_LC_2_28_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i42_LC_2_28_1  (
            .in0(N__36787),
            .in1(N__36041),
            .in2(N__17436),
            .in3(N__13423),
            .lcout(\c0.data_in_field_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5440_LC_2_28_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5440_LC_2_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5440_LC_2_28_2 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5440_LC_2_28_2  (
            .in0(N__33274),
            .in1(N__26271),
            .in2(N__24964),
            .in3(N__32516),
            .lcout(),
            .ltout(\c0.n5803_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5803_bdd_4_lut_LC_2_28_3 .C_ON=1'b0;
    defparam \c0.n5803_bdd_4_lut_LC_2_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5803_bdd_4_lut_LC_2_28_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5803_bdd_4_lut_LC_2_28_3  (
            .in0(N__32517),
            .in1(N__25057),
            .in2(N__12958),
            .in3(N__19984),
            .lcout(\c0.n5426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i22_LC_2_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i22_LC_2_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i22_LC_2_28_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i22_LC_2_28_5  (
            .in0(N__16111),
            .in1(N__36040),
            .in2(N__37000),
            .in3(N__23739),
            .lcout(\c0.data_in_field_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i149_LC_2_28_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i149_LC_2_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i149_LC_2_28_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i149_LC_2_28_6  (
            .in0(N__26795),
            .in1(N__37334),
            .in2(_gnd_net_),
            .in3(N__34295),
            .lcout(data_in_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_909_LC_2_28_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_909_LC_2_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_909_LC_2_28_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_909_LC_2_28_7  (
            .in0(N__32022),
            .in1(N__29535),
            .in2(_gnd_net_),
            .in3(N__22245),
            .lcout(\c0.n16_adj_1922 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i146_LC_2_29_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i146_LC_2_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i146_LC_2_29_0 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0___i146_LC_2_29_0  (
            .in0(N__13137),
            .in1(N__37124),
            .in2(N__36261),
            .in3(N__20086),
            .lcout(\c0.data_in_frame_18_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i156_LC_2_29_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i156_LC_2_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i156_LC_2_29_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i156_LC_2_29_1  (
            .in0(N__34151),
            .in1(N__14797),
            .in2(_gnd_net_),
            .in3(N__15853),
            .lcout(data_in_19_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5671_bdd_4_lut_LC_2_29_2 .C_ON=1'b0;
    defparam \c0.n5671_bdd_4_lut_LC_2_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.n5671_bdd_4_lut_LC_2_29_2 .LUT_INIT=16'b1010111010100100;
    LogicCell40 \c0.n5671_bdd_4_lut_LC_2_29_2  (
            .in0(N__14803),
            .in1(N__17509),
            .in2(N__32593),
            .in3(N__25501),
            .lcout(\c0.n5369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5495_LC_2_29_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5495_LC_2_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5495_LC_2_29_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5495_LC_2_29_4  (
            .in0(N__33236),
            .in1(N__23623),
            .in2(N__32594),
            .in3(N__26953),
            .lcout(\c0.n5869 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5959_bdd_4_lut_LC_2_29_5 .C_ON=1'b0;
    defparam \c0.n5959_bdd_4_lut_LC_2_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.n5959_bdd_4_lut_LC_2_29_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5959_bdd_4_lut_LC_2_29_5  (
            .in0(N__32587),
            .in1(N__14692),
            .in2(N__13105),
            .in3(N__25009),
            .lcout(\c0.n5962 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i148_LC_2_29_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i148_LC_2_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i148_LC_2_29_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0___i148_LC_2_29_6  (
            .in0(N__13083),
            .in1(N__37125),
            .in2(N__36262),
            .in3(N__14647),
            .lcout(\c0.data_in_frame_18_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i6_LC_2_30_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i6_LC_2_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_2_30_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_2_30_0  (
            .in0(N__13240),
            .in1(N__14882),
            .in2(_gnd_net_),
            .in3(N__13069),
            .lcout(r_Clock_Count_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_2_30_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_2_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_2_30_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_2_30_1  (
            .in0(N__18056),
            .in1(N__18138),
            .in2(N__18355),
            .in3(N__18281),
            .lcout(r_SM_Main_2_adj_2005),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_878_LC_2_30_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_878_LC_2_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_878_LC_2_30_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_878_LC_2_30_2  (
            .in0(N__19800),
            .in1(N__22573),
            .in2(N__24434),
            .in3(N__28030),
            .lcout(\c0.n15_adj_1894 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_2_30_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i0_LC_2_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_2_30_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_2_30_3  (
            .in0(N__14912),
            .in1(N__13192),
            .in2(_gnd_net_),
            .in3(N__13241),
            .lcout(r_Clock_Count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i4_LC_2_30_4 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i4_LC_2_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_2_30_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_2_30_4  (
            .in0(N__13186),
            .in1(N__13243),
            .in2(_gnd_net_),
            .in3(N__13375),
            .lcout(\c0.rx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_4_lut_LC_2_30_5 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_4_lut_LC_2_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_4_lut_LC_2_30_5 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \c0.rx.i1_4_lut_4_lut_LC_2_30_5  (
            .in0(N__18055),
            .in1(N__18137),
            .in2(N__18354),
            .in3(N__18280),
            .lcout(\c0.rx.n2157 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i5_LC_2_30_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i5_LC_2_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_2_30_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_2_30_6  (
            .in0(N__13239),
            .in1(N__13399),
            .in2(_gnd_net_),
            .in3(N__13174),
            .lcout(\c0.rx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i3_LC_2_30_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i3_LC_2_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_2_30_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_2_30_7  (
            .in0(N__13242),
            .in1(N__13309),
            .in2(_gnd_net_),
            .in3(N__13168),
            .lcout(\c0.rx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35329),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_794_LC_2_31_0 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_794_LC_2_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_794_LC_2_31_0 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \c0.rx.i1_4_lut_adj_794_LC_2_31_0  (
            .in0(N__14766),
            .in1(N__13162),
            .in2(N__14884),
            .in3(N__13351),
            .lcout(\c0.rx.r_SM_Main_2_N_1824_2 ),
            .ltout(\c0.rx.r_SM_Main_2_N_1824_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_3_lut_LC_2_31_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_3_lut_LC_2_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_3_lut_LC_2_31_1 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \c0.rx.i1_2_lut_3_lut_LC_2_31_1  (
            .in0(_gnd_net_),
            .in1(N__18328),
            .in2(N__13156),
            .in3(N__18276),
            .lcout(n4474),
            .ltout(n4474_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_796_LC_2_31_2 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_796_LC_2_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_796_LC_2_31_2 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \c0.rx.i1_4_lut_adj_796_LC_2_31_2  (
            .in0(N__18329),
            .in1(N__13147),
            .in2(N__13141),
            .in3(N__13281),
            .lcout(),
            .ltout(\c0.rx.n4_adj_1866_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3748_2_lut_LC_2_31_3 .C_ON=1'b0;
    defparam \c0.rx.i3748_2_lut_LC_2_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3748_2_lut_LC_2_31_3 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \c0.rx.i3748_2_lut_LC_2_31_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13453),
            .in3(N__13222),
            .lcout(\c0.rx.n4011 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i42_LC_2_31_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i42_LC_2_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i42_LC_2_31_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i42_LC_2_31_5  (
            .in0(N__23956),
            .in1(_gnd_net_),
            .in2(N__34363),
            .in3(N__13410),
            .lcout(data_in_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35337),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_793_LC_2_31_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_793_LC_2_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_793_LC_2_31_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_adj_793_LC_2_31_6  (
            .in0(_gnd_net_),
            .in1(N__13396),
            .in2(_gnd_net_),
            .in3(N__13372),
            .lcout(\c0.rx.n37 ),
            .ltout(\c0.rx.n37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i4_4_lut_LC_2_31_7 .C_ON=1'b0;
    defparam \c0.rx.i4_4_lut_LC_2_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i4_4_lut_LC_2_31_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.rx.i4_4_lut_LC_2_31_7  (
            .in0(N__14701),
            .in1(N__13340),
            .in2(N__13312),
            .in3(N__13307),
            .lcout(r_SM_Main_2_N_1830_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_LC_2_32_0 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_LC_2_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_LC_2_32_0 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \c0.rx.i2_4_lut_LC_2_32_0  (
            .in0(N__18247),
            .in1(N__18111),
            .in2(N__18356),
            .in3(N__18049),
            .lcout(\c0.rx.n2213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_2_32_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_2_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_2_32_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_2_32_1  (
            .in0(N__13258),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35344),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_29_i4_2_lut_LC_2_32_2 .C_ON=1'b0;
    defparam \c0.rx.equal_29_i4_2_lut_LC_2_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_29_i4_2_lut_LC_2_32_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.equal_29_i4_2_lut_LC_2_32_2  (
            .in0(N__14963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14934),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5_4_lut_LC_2_32_3 .C_ON=1'b0;
    defparam \c0.rx.i5_4_lut_LC_2_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5_4_lut_LC_2_32_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.rx.i5_4_lut_LC_2_32_3  (
            .in0(N__18110),
            .in1(N__18246),
            .in2(N__20915),
            .in3(N__14729),
            .lcout(),
            .ltout(n12_adj_1995_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_1012_LC_2_32_4.C_ON=1'b0;
    defparam i1_4_lut_adj_1012_LC_2_32_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_1012_LC_2_32_4.LUT_INIT=16'b1010101011101010;
    LogicCell40 i1_4_lut_adj_1012_LC_2_32_4 (
            .in0(N__18337),
            .in1(N__14848),
            .in2(N__13252),
            .in3(N__13249),
            .lcout(n16_adj_1993),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_3_lut_LC_2_32_5 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_3_lut_LC_2_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_3_lut_LC_2_32_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i2_2_lut_3_lut_LC_2_32_5  (
            .in0(N__14933),
            .in1(N__18176),
            .in2(_gnd_net_),
            .in3(N__14962),
            .lcout(\c0.rx.n3573 ),
            .ltout(\c0.rx.n3573_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2073_2_lut_3_lut_LC_2_32_6 .C_ON=1'b0;
    defparam \c0.rx.i2073_2_lut_3_lut_LC_2_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2073_2_lut_3_lut_LC_2_32_6 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \c0.rx.i2073_2_lut_3_lut_LC_2_32_6  (
            .in0(N__18248),
            .in1(_gnd_net_),
            .in2(N__13492),
            .in3(N__14988),
            .lcout(\c0.rx.n2317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i36_LC_2_32_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i36_LC_2_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i36_LC_2_32_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i36_LC_2_32_7  (
            .in0(N__34152),
            .in1(N__26584),
            .in2(_gnd_net_),
            .in3(N__17669),
            .lcout(data_in_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35344),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_3_15_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_3_15_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_3_15_2  (
            .in0(N__20639),
            .in1(N__20739),
            .in2(N__18817),
            .in3(N__16430),
            .lcout(n4_adj_1988),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_1794_LC_3_16_0 .C_ON=1'b0;
    defparam \c0.tx_transmit_1794_LC_3_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_1794_LC_3_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.tx_transmit_1794_LC_3_16_0  (
            .in0(N__13549),
            .in1(N__13541),
            .in2(N__13723),
            .in3(N__13656),
            .lcout(\c0.tx_transmit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35275),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_902_LC_3_16_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_902_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_902_LC_3_16_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_902_LC_3_16_1  (
            .in0(N__14818),
            .in1(N__15036),
            .in2(N__15082),
            .in3(N__15181),
            .lcout(),
            .ltout(\c0.n20_adj_1918_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_906_LC_3_16_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_906_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_906_LC_3_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_906_LC_3_16_2  (
            .in0(N__15057),
            .in1(N__15111),
            .in2(N__13489),
            .in3(N__13459),
            .lcout(n21_adj_1999),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_939_LC_3_16_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_939_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_939_LC_3_16_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_939_LC_3_16_4  (
            .in0(N__13710),
            .in1(N__19167),
            .in2(_gnd_net_),
            .in3(N__13655),
            .lcout(\c0.n87 ),
            .ltout(\c0.n87_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i4_LC_3_16_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i4_LC_3_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i4_LC_3_16_5 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \c0.byte_transmit_counter__i4_LC_3_16_5  (
            .in0(N__13540),
            .in1(N__13582),
            .in2(N__13462),
            .in3(N__13561),
            .lcout(\c0.byte_transmit_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35275),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_LC_3_16_7 .C_ON=1'b0;
    defparam \c0.i5_2_lut_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_LC_3_16_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i5_2_lut_LC_3_16_7  (
            .in0(_gnd_net_),
            .in1(N__15096),
            .in2(_gnd_net_),
            .in3(N__14835),
            .lcout(\c0.n16_adj_1909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i14_LC_3_17_0 .C_ON=1'b0;
    defparam \c0.data_out_0___i14_LC_3_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i14_LC_3_17_0 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.data_out_0___i14_LC_3_17_0  (
            .in0(N__19174),
            .in1(N__20730),
            .in2(N__18406),
            .in3(N__19033),
            .lcout(data_out_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35270),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_913_LC_3_17_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_913_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_913_LC_3_17_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_913_LC_3_17_2  (
            .in0(N__13617),
            .in1(N__13605),
            .in2(_gnd_net_),
            .in3(N__13593),
            .lcout(\c0.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i119_2_lut_LC_3_17_3 .C_ON=1'b0;
    defparam \c0.i119_2_lut_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i119_2_lut_LC_3_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i119_2_lut_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__13579),
            .in2(_gnd_net_),
            .in3(N__13560),
            .lcout(\c0.n109 ),
            .ltout(\c0.n109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5298_3_lut_4_lut_LC_3_17_4 .C_ON=1'b0;
    defparam \c0.i5298_3_lut_4_lut_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5298_3_lut_4_lut_LC_3_17_4 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \c0.i5298_3_lut_4_lut_LC_3_17_4  (
            .in0(N__13702),
            .in1(N__13539),
            .in2(N__13519),
            .in3(N__13654),
            .lcout(n4315),
            .ltout(n4315_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i12_LC_3_17_5 .C_ON=1'b0;
    defparam \c0.data_out_0___i12_LC_3_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i12_LC_3_17_5 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \c0.data_out_0___i12_LC_3_17_5  (
            .in0(N__18427),
            .in1(N__16565),
            .in2(N__13516),
            .in3(N__19175),
            .lcout(data_out_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35270),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i29_LC_3_17_6 .C_ON=1'b0;
    defparam \c0.data_out_0___i29_LC_3_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i29_LC_3_17_6 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \c0.data_out_0___i29_LC_3_17_6  (
            .in0(N__16711),
            .in1(N__13777),
            .in2(N__16144),
            .in3(N__16673),
            .lcout(data_out_19_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35270),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i15_LC_3_17_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i15_LC_3_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i15_LC_3_17_7 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_out_0___i15_LC_3_17_7  (
            .in0(N__19034),
            .in1(N__18382),
            .in2(N__20640),
            .in3(N__19176),
            .lcout(data_out_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35270),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i10_LC_3_18_0 .C_ON=1'b0;
    defparam \c0.data_out_0___i10_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i10_LC_3_18_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0___i10_LC_3_18_0  (
            .in0(N__19029),
            .in1(N__16807),
            .in2(N__18472),
            .in3(N__19179),
            .lcout(data_out_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i6_LC_3_18_1 .C_ON=1'b0;
    defparam \c0.data_out_0___i6_LC_3_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i6_LC_3_18_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.data_out_0___i6_LC_3_18_1  (
            .in0(N__19178),
            .in1(N__21109),
            .in2(N__18535),
            .in3(N__19032),
            .lcout(data_out_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i5_LC_3_18_2 .C_ON=1'b0;
    defparam \c0.data_out_0___i5_LC_3_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i5_LC_3_18_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_out_0___i5_LC_3_18_2  (
            .in0(N__19031),
            .in1(N__18553),
            .in2(N__18749),
            .in3(N__19181),
            .lcout(data_out_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i27_LC_3_18_3 .C_ON=1'b0;
    defparam \c0.data_out_0___i27_LC_3_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i27_LC_3_18_3 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \c0.data_out_0___i27_LC_3_18_3  (
            .in0(N__16227),
            .in1(N__16186),
            .in2(N__15493),
            .in3(N__16666),
            .lcout(data_out_19_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i4_LC_3_18_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i4_LC_3_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i4_LC_3_18_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0___i4_LC_3_18_4  (
            .in0(N__19030),
            .in1(N__21012),
            .in2(N__18574),
            .in3(N__19180),
            .lcout(data_out_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_943_LC_3_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_943_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_943_LC_3_18_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.i1_2_lut_adj_943_LC_3_18_5  (
            .in0(N__19177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19028),
            .lcout(n4316),
            .ltout(n4316_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i20_LC_3_18_6 .C_ON=1'b0;
    defparam \c0.data_out_0___i20_LC_3_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i20_LC_3_18_6 .LUT_INIT=16'b1100101011000101;
    LogicCell40 \c0.data_out_0___i20_LC_3_18_6  (
            .in0(N__20979),
            .in1(N__15357),
            .in2(N__13684),
            .in3(N__15163),
            .lcout(data_out_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i25_LC_3_18_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i25_LC_3_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i25_LC_3_18_7 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \c0.data_out_0___i25_LC_3_18_7  (
            .in0(N__15249),
            .in1(N__13747),
            .in2(N__13681),
            .in3(N__16665),
            .lcout(data_out_19_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_4_lut_LC_3_19_0 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_4_lut_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_4_lut_LC_3_19_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx.i2_3_lut_4_lut_LC_3_19_0  (
            .in0(N__13724),
            .in1(N__17121),
            .in2(N__17002),
            .in3(N__17062),
            .lcout(n1442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i21_LC_3_19_2 .C_ON=1'b0;
    defparam \c0.data_out_0___i21_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i21_LC_3_19_2 .LUT_INIT=16'b1100110010100101;
    LogicCell40 \c0.data_out_0___i21_LC_3_19_2  (
            .in0(N__13672),
            .in1(N__13762),
            .in2(N__15274),
            .in3(N__16671),
            .lcout(data_out_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35279),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_3_19_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_3_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_3_19_3 .LUT_INIT=16'b1111000001110100;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_3_19_3  (
            .in0(N__17122),
            .in1(N__13735),
            .in2(N__13657),
            .in3(N__16996),
            .lcout(tx_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35279),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_3_19_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_3_19_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_3_19_4  (
            .in0(N__13776),
            .in1(N__20393),
            .in2(_gnd_net_),
            .in3(N__13761),
            .lcout(),
            .ltout(\c0.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_3_19_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_3_19_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_3_19_5  (
            .in0(N__21186),
            .in1(N__18706),
            .in2(N__13753),
            .in3(N__20683),
            .lcout(),
            .ltout(tx_data_4_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_3_19_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_3_19_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_3_19_6  (
            .in0(N__16827),
            .in1(_gnd_net_),
            .in2(N__13750),
            .in3(N__19340),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35279),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i16_LC_3_20_0 .C_ON=1'b0;
    defparam \c0.data_out_0___i16_LC_3_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i16_LC_3_20_0 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i16_LC_3_20_0  (
            .in0(N__16416),
            .in1(N__19220),
            .in2(N__18628),
            .in3(N__19058),
            .lcout(data_out_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35285),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_LC_3_20_3 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_LC_3_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_LC_3_20_3  (
            .in0(N__16474),
            .in1(N__19300),
            .in2(N__16378),
            .in3(N__21079),
            .lcout(n8_adj_2001),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_3_20_4 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_3_20_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i1_2_lut_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__14022),
            .in2(_gnd_net_),
            .in3(N__13995),
            .lcout(\c0.tx.r_SM_Main_2_N_1767_1 ),
            .ltout(\c0.tx.r_SM_Main_2_N_1767_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5288_3_lut_4_lut_4_lut_LC_3_20_5 .C_ON=1'b0;
    defparam \c0.tx.i5288_3_lut_4_lut_4_lut_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5288_3_lut_4_lut_4_lut_LC_3_20_5 .LUT_INIT=16'b1100000000100010;
    LogicCell40 \c0.tx.i5288_3_lut_4_lut_4_lut_LC_3_20_5  (
            .in0(N__13725),
            .in1(N__17116),
            .in2(N__13738),
            .in3(N__17058),
            .lcout(n5041),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_3_21_0 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_3_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_3_21_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_3_21_0  (
            .in0(N__17120),
            .in1(N__17049),
            .in2(N__16997),
            .in3(N__15405),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_3_21_1 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_3_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_3_21_1 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_3_21_1  (
            .in0(N__15404),
            .in1(N__16972),
            .in2(N__17060),
            .in3(N__17119),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i29_4_lut_LC_3_21_2 .C_ON=1'b0;
    defparam \c0.tx.i29_4_lut_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i29_4_lut_LC_3_21_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \c0.tx.i29_4_lut_LC_3_21_2  (
            .in0(N__13729),
            .in1(N__17098),
            .in2(N__15385),
            .in3(N__15403),
            .lcout(),
            .ltout(\c0.tx.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_3_21_3 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_3_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_3_21_3 .LUT_INIT=16'b0001000100110000;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_3_21_3  (
            .in0(N__15406),
            .in1(N__16967),
            .in2(N__14029),
            .in3(N__17059),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1066_2_lut_LC_3_21_4 .C_ON=1'b0;
    defparam \c0.tx.i1066_2_lut_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1066_2_lut_LC_3_21_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i1066_2_lut_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(N__17097),
            .in2(_gnd_net_),
            .in3(N__17044),
            .lcout(n1307),
            .ltout(n1307_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_adj_802_LC_3_21_5 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_adj_802_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_adj_802_LC_3_21_5 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \c0.tx.i1_4_lut_adj_802_LC_3_21_5  (
            .in0(N__16949),
            .in1(N__14023),
            .in2(N__13999),
            .in3(N__13996),
            .lcout(n4221),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_3_21_6.C_ON=1'b0;
    defparam i1_4_lut_LC_3_21_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_3_21_6.LUT_INIT=16'b1110101011100000;
    LogicCell40 i1_4_lut_LC_3_21_6 (
            .in0(N__17118),
            .in1(N__17045),
            .in2(N__13927),
            .in3(N__13942),
            .lcout(),
            .ltout(n4_adj_2003_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Done_44_LC_3_21_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Done_44_LC_3_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Done_44_LC_3_21_7 .LUT_INIT=16'b1111101111110000;
    LogicCell40 \c0.tx.r_Tx_Done_44_LC_3_21_7  (
            .in0(N__13926),
            .in1(N__13936),
            .in2(N__13930),
            .in3(N__16968),
            .lcout(n4155),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i7_LC_3_22_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i7_LC_3_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i7_LC_3_22_0 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \c0.tx2.r_Clock_Count__i7_LC_3_22_0  (
            .in0(N__14097),
            .in1(_gnd_net_),
            .in2(N__13912),
            .in3(N__14234),
            .lcout(\c0.tx2.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i2_LC_3_22_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i2_LC_3_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i2_LC_3_22_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i2_LC_3_22_3  (
            .in0(N__14233),
            .in1(N__13885),
            .in2(_gnd_net_),
            .in3(N__14096),
            .lcout(\c0.tx2.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_3_lut_4_lut_LC_3_22_4 .C_ON=1'b0;
    defparam \c0.tx2.i1_3_lut_4_lut_LC_3_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_3_lut_4_lut_LC_3_22_4 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.tx2.i1_3_lut_4_lut_LC_3_22_4  (
            .in0(N__13855),
            .in1(N__14232),
            .in2(N__14389),
            .in3(N__13795),
            .lcout(\c0.tx2.n2218 ),
            .ltout(\c0.tx2.n2218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2075_2_lut_3_lut_LC_3_22_5 .C_ON=1'b0;
    defparam \c0.tx2.i2075_2_lut_3_lut_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2075_2_lut_3_lut_LC_3_22_5 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \c0.tx2.i2075_2_lut_3_lut_LC_3_22_5  (
            .in0(_gnd_net_),
            .in1(N__14368),
            .in2(N__14326),
            .in3(N__14323),
            .lcout(\c0.tx2.n2319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5953_bdd_4_lut_LC_3_23_1 .C_ON=1'b0;
    defparam \c0.n5953_bdd_4_lut_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5953_bdd_4_lut_LC_3_23_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5953_bdd_4_lut_LC_3_23_1  (
            .in0(N__32319),
            .in1(N__28861),
            .in2(N__14296),
            .in3(N__27433),
            .lcout(\c0.n5956 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i3_LC_3_23_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i3_LC_3_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i3_LC_3_23_3 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i3_LC_3_23_3  (
            .in0(N__14269),
            .in1(N__14207),
            .in2(_gnd_net_),
            .in3(N__14101),
            .lcout(\c0.tx2.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i15_LC_3_23_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i15_LC_3_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i15_LC_3_23_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i15_LC_3_23_5  (
            .in0(N__23864),
            .in1(N__34283),
            .in2(_gnd_net_),
            .in3(N__27892),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i93_LC_3_23_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i93_LC_3_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i93_LC_3_23_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i93_LC_3_23_6  (
            .in0(N__34282),
            .in1(N__28708),
            .in2(_gnd_net_),
            .in3(N__27038),
            .lcout(data_in_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_525_526__i1_LC_3_24_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_525_526__i1_LC_3_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i1_LC_3_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i1_LC_3_24_0  (
            .in0(_gnd_net_),
            .in1(N__33116),
            .in2(N__15823),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter2_0 ),
            .ltout(),
            .carryin(bfn_3_24_0_),
            .carryout(\c0.n4400 ),
            .clk(N__35307),
            .ce(N__15733),
            .sr(N__15721));
    defparam \c0.byte_transmit_counter2_525_526__i2_LC_3_24_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_525_526__i2_LC_3_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i2_LC_3_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i2_LC_3_24_1  (
            .in0(_gnd_net_),
            .in1(N__32320),
            .in2(_gnd_net_),
            .in3(N__14038),
            .lcout(\c0.byte_transmit_counter2_1 ),
            .ltout(),
            .carryin(\c0.n4400 ),
            .carryout(\c0.n4401 ),
            .clk(N__35307),
            .ce(N__15733),
            .sr(N__15721));
    defparam \c0.byte_transmit_counter2_525_526__i3_LC_3_24_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_525_526__i3_LC_3_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i3_LC_3_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i3_LC_3_24_2  (
            .in0(_gnd_net_),
            .in1(N__32098),
            .in2(_gnd_net_),
            .in3(N__14035),
            .lcout(\c0.byte_transmit_counter2_2 ),
            .ltout(),
            .carryin(\c0.n4401 ),
            .carryout(\c0.n4402 ),
            .clk(N__35307),
            .ce(N__15733),
            .sr(N__15721));
    defparam \c0.byte_transmit_counter2_525_526__i4_LC_3_24_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_525_526__i4_LC_3_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i4_LC_3_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i4_LC_3_24_3  (
            .in0(_gnd_net_),
            .in1(N__34762),
            .in2(_gnd_net_),
            .in3(N__14032),
            .lcout(\c0.byte_transmit_counter2_3 ),
            .ltout(),
            .carryin(\c0.n4402 ),
            .carryout(\c0.n4403 ),
            .clk(N__35307),
            .ce(N__15733),
            .sr(N__15721));
    defparam \c0.byte_transmit_counter2_525_526__i5_LC_3_24_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_525_526__i5_LC_3_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i5_LC_3_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i5_LC_3_24_4  (
            .in0(_gnd_net_),
            .in1(N__14505),
            .in2(_gnd_net_),
            .in3(N__14536),
            .lcout(\c0.byte_transmit_counter2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35307),
            .ce(N__15733),
            .sr(N__15721));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5455_LC_3_25_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5455_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5455_LC_3_25_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5455_LC_3_25_1  (
            .in0(N__32097),
            .in1(N__21751),
            .in2(N__34800),
            .in3(N__21775),
            .lcout(),
            .ltout(\c0.n5785_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5785_bdd_4_lut_LC_3_25_2 .C_ON=1'b0;
    defparam \c0.n5785_bdd_4_lut_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.n5785_bdd_4_lut_LC_3_25_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n5785_bdd_4_lut_LC_3_25_2  (
            .in0(N__21853),
            .in1(N__34761),
            .in2(N__14470),
            .in3(N__14467),
            .lcout(\c0.n5788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5965_bdd_4_lut_LC_3_25_3 .C_ON=1'b0;
    defparam \c0.n5965_bdd_4_lut_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5965_bdd_4_lut_LC_3_25_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5965_bdd_4_lut_LC_3_25_3  (
            .in0(N__32318),
            .in1(N__28396),
            .in2(N__17386),
            .in3(N__28438),
            .lcout(\c0.n5968 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i28_LC_3_25_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i28_LC_3_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i28_LC_3_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i28_LC_3_25_6  (
            .in0(N__34219),
            .in1(N__17686),
            .in2(_gnd_net_),
            .in3(N__23305),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35311),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5809_bdd_4_lut_LC_3_25_7 .C_ON=1'b0;
    defparam \c0.n5809_bdd_4_lut_LC_3_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.n5809_bdd_4_lut_LC_3_25_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5809_bdd_4_lut_LC_3_25_7  (
            .in0(N__32317),
            .in1(N__30358),
            .in2(N__19417),
            .in3(N__20119),
            .lcout(\c0.n5363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i160_LC_3_26_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i160_LC_3_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i160_LC_3_26_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i160_LC_3_26_0  (
            .in0(N__14427),
            .in1(N__20164),
            .in2(N__37003),
            .in3(N__36199),
            .lcout(\c0.data_in_frame_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5548_LC_3_26_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5548_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5548_LC_3_26_1 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5548_LC_3_26_1  (
            .in0(N__16129),
            .in1(N__33181),
            .in2(N__14559),
            .in3(N__32446),
            .lcout(\c0.n5935 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i102_LC_3_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i102_LC_3_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i102_LC_3_26_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i102_LC_3_26_2  (
            .in0(N__36798),
            .in1(N__36198),
            .in2(N__16039),
            .in3(N__15963),
            .lcout(\c0.data_in_field_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i158_LC_3_26_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i158_LC_3_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i158_LC_3_26_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i158_LC_3_26_3  (
            .in0(N__34215),
            .in1(N__14782),
            .in2(_gnd_net_),
            .in3(N__24505),
            .lcout(data_in_19_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i94_LC_3_26_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i94_LC_3_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i94_LC_3_26_4 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \c0.data_in_0___i94_LC_3_26_4  (
            .in0(N__16035),
            .in1(N__34216),
            .in2(N__26983),
            .in3(_gnd_net_),
            .lcout(data_in_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5941_bdd_4_lut_LC_3_26_5 .C_ON=1'b0;
    defparam \c0.n5941_bdd_4_lut_LC_3_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.n5941_bdd_4_lut_LC_3_26_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5941_bdd_4_lut_LC_3_26_5  (
            .in0(N__32447),
            .in1(N__23932),
            .in2(N__18904),
            .in3(N__20050),
            .lcout(\c0.n5944 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i86_LC_3_26_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i86_LC_3_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i86_LC_3_26_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i86_LC_3_26_6  (
            .in0(N__26978),
            .in1(N__34217),
            .in2(_gnd_net_),
            .in3(N__27528),
            .lcout(data_in_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_3_lut_4_lut_LC_3_26_7 .C_ON=1'b0;
    defparam \c0.i10_3_lut_4_lut_LC_3_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10_3_lut_4_lut_LC_3_26_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_3_lut_4_lut_LC_3_26_7  (
            .in0(N__14614),
            .in1(N__22198),
            .in2(N__22399),
            .in3(N__22165),
            .lcout(\c0.n23_adj_1931 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i14_LC_3_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i14_LC_3_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i14_LC_3_27_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i14_LC_3_27_0  (
            .in0(N__24154),
            .in1(N__36272),
            .in2(N__37002),
            .in3(N__21707),
            .lcout(\c0.data_in_field_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i12_LC_3_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i12_LC_3_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i12_LC_3_27_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i12_LC_3_27_2  (
            .in0(N__21875),
            .in1(N__22375),
            .in2(N__37001),
            .in3(N__36273),
            .lcout(\c0.data_in_field_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i159_LC_3_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i159_LC_3_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i159_LC_3_27_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i159_LC_3_27_3  (
            .in0(N__36271),
            .in1(N__36791),
            .in2(N__14560),
            .in3(N__17370),
            .lcout(\c0.data_in_frame_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5743_bdd_4_lut_LC_3_27_4 .C_ON=1'b0;
    defparam \c0.n5743_bdd_4_lut_LC_3_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.n5743_bdd_4_lut_LC_3_27_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5743_bdd_4_lut_LC_3_27_4  (
            .in0(N__32543),
            .in1(N__17422),
            .in2(N__19852),
            .in3(N__29302),
            .lcout(\c0.n5456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_975_LC_3_27_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_975_LC_3_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_975_LC_3_27_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_975_LC_3_27_5  (
            .in0(N__23618),
            .in1(N__21579),
            .in2(_gnd_net_),
            .in3(N__19935),
            .lcout(\c0.n1893 ),
            .ltout(\c0.n1893_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_907_LC_3_27_6 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_907_LC_3_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_907_LC_3_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_907_LC_3_27_6  (
            .in0(N__19503),
            .in1(N__14635),
            .in2(N__14617),
            .in3(N__28395),
            .lcout(\c0.n20_adj_1921 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_849_LC_3_27_7 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_849_LC_3_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_849_LC_3_27_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_849_LC_3_27_7  (
            .in0(N__17421),
            .in1(N__21874),
            .in2(N__17508),
            .in3(N__17277),
            .lcout(\c0.n1821 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_846_LC_3_28_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_846_LC_3_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_846_LC_3_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_846_LC_3_28_1  (
            .in0(N__15958),
            .in1(N__31344),
            .in2(_gnd_net_),
            .in3(N__14689),
            .lcout(\c0.n5072 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_891_LC_3_28_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_891_LC_3_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_891_LC_3_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_891_LC_3_28_2  (
            .in0(N__19518),
            .in1(N__23638),
            .in2(N__19804),
            .in3(N__25810),
            .lcout(\c0.n24_adj_1907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i132_LC_3_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i132_LC_3_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i132_LC_3_28_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i132_LC_3_28_3  (
            .in0(N__36786),
            .in1(N__36013),
            .in2(N__26835),
            .in3(N__14690),
            .lcout(\c0.data_in_field_131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35323),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5737_bdd_4_lut_LC_3_28_6 .C_ON=1'b0;
    defparam \c0.n5737_bdd_4_lut_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.n5737_bdd_4_lut_LC_3_28_6 .LUT_INIT=16'b1010111010100100;
    LogicCell40 \c0.n5737_bdd_4_lut_LC_3_28_6  (
            .in0(N__14602),
            .in1(N__30271),
            .in2(N__32595),
            .in3(N__20017),
            .lcout(\c0.n5459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_3_28_7 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_3_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_3_28_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_LC_3_28_7  (
            .in0(N__24640),
            .in1(N__17435),
            .in2(N__24223),
            .in3(N__28437),
            .lcout(\c0.n22_adj_1881 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5385_LC_3_29_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5385_LC_3_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5385_LC_3_29_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5385_LC_3_29_0  (
            .in0(N__33237),
            .in1(N__23554),
            .in2(N__32545),
            .in3(N__15701),
            .lcout(\c0.n5737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i82_LC_3_29_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i82_LC_3_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i82_LC_3_29_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i82_LC_3_29_1  (
            .in0(N__15702),
            .in1(N__28573),
            .in2(N__36200),
            .in3(N__37123),
            .lcout(\c0.data_in_field_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i154_LC_3_29_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i154_LC_3_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i154_LC_3_29_2 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0___i154_LC_3_29_2  (
            .in0(N__14586),
            .in1(N__36006),
            .in2(N__37226),
            .in3(N__17878),
            .lcout(\c0.data_in_frame_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i120_LC_3_29_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i120_LC_3_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i120_LC_3_29_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i120_LC_3_29_3  (
            .in0(N__36005),
            .in1(N__37116),
            .in2(N__21667),
            .in3(N__17725),
            .lcout(\c0.data_in_field_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i20_LC_3_29_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i20_LC_3_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i20_LC_3_29_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i20_LC_3_29_4  (
            .in0(N__23354),
            .in1(N__17845),
            .in2(N__37227),
            .in3(N__36010),
            .lcout(\c0.data_in_field_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_832_LC_3_29_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_832_LC_3_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_832_LC_3_29_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_832_LC_3_29_5  (
            .in0(N__15700),
            .in1(N__23353),
            .in2(N__23740),
            .in3(N__14691),
            .lcout(\c0.n2036 ),
            .ltout(\c0.n2036_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_834_LC_3_29_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_834_LC_3_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_834_LC_3_29_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_834_LC_3_29_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14671),
            .in3(N__24956),
            .lcout(),
            .ltout(\c0.n5273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_3_29_7 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_3_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_3_29_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_LC_3_29_7  (
            .in0(N__19470),
            .in1(N__24579),
            .in2(N__14668),
            .in3(N__25939),
            .lcout(\c0.n42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i4_LC_3_30_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i4_LC_3_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i4_LC_3_30_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i4_LC_3_30_0  (
            .in0(N__34030),
            .in1(N__31731),
            .in2(_gnd_net_),
            .in3(N__22371),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i152_LC_3_30_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i152_LC_3_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i152_LC_3_30_1 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0___i152_LC_3_30_1  (
            .in0(N__14661),
            .in1(N__36146),
            .in2(N__37203),
            .in3(N__26043),
            .lcout(\c0.data_in_frame_18_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i151_LC_3_30_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i151_LC_3_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i151_LC_3_30_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i151_LC_3_30_2  (
            .in0(N__34029),
            .in1(N__17359),
            .in2(_gnd_net_),
            .in3(N__24211),
            .lcout(data_in_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i127_LC_3_30_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i127_LC_3_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i127_LC_3_30_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i127_LC_3_30_5  (
            .in0(N__23672),
            .in1(N__34031),
            .in2(_gnd_net_),
            .in3(N__17934),
            .lcout(data_in_15_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5336_LC_3_30_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5336_LC_3_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5336_LC_3_30_7 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5336_LC_3_30_7  (
            .in0(N__33117),
            .in1(N__19834),
            .in2(N__32589),
            .in3(N__23007),
            .lcout(\c0.n5671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i17_LC_3_31_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i17_LC_3_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i17_LC_3_31_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i17_LC_3_31_0  (
            .in0(N__31439),
            .in1(N__31528),
            .in2(_gnd_net_),
            .in3(N__33881),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35345),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_3_31_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_3_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_3_31_1 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_3_31_1  (
            .in0(N__14793),
            .in1(N__20859),
            .in2(N__20930),
            .in3(N__17964),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35345),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i138_LC_3_31_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i138_LC_3_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i138_LC_3_31_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i138_LC_3_31_3  (
            .in0(N__33880),
            .in1(N__20798),
            .in2(_gnd_net_),
            .in3(N__20084),
            .lcout(data_in_17_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35345),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i22_LC_3_31_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i22_LC_3_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i22_LC_3_31_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i22_LC_3_31_4  (
            .in0(N__33885),
            .in1(N__16107),
            .in2(_gnd_net_),
            .in3(N__27967),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35345),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i20_LC_3_31_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i20_LC_3_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i20_LC_3_31_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i20_LC_3_31_5  (
            .in0(N__33882),
            .in1(N__23312),
            .in2(_gnd_net_),
            .in3(N__17837),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35345),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_3_31_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_3_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_3_31_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_3_31_6  (
            .in0(N__20911),
            .in1(N__14778),
            .in2(N__20863),
            .in3(N__16170),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35345),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_LC_3_31_7 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_LC_3_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_LC_3_31_7 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \c0.rx.i1_4_lut_LC_3_31_7  (
            .in0(N__14874),
            .in1(N__14765),
            .in2(N__14913),
            .in3(N__14731),
            .lcout(\c0.rx.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_26_i4_2_lut_LC_3_32_0 .C_ON=1'b0;
    defparam \c0.rx.equal_26_i4_2_lut_LC_3_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_26_i4_2_lut_LC_3_32_0 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \c0.rx.equal_26_i4_2_lut_LC_3_32_0  (
            .in0(N__14965),
            .in1(N__14938),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n4_adj_1990),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_3_32_1 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_3_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_3_32_1 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_3_32_1  (
            .in0(N__14940),
            .in1(_gnd_net_),
            .in2(N__18184),
            .in3(N__14967),
            .lcout(\c0.rx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35352),
            .ce(N__14992),
            .sr(N__14977));
    defparam \c0.rx.r_Bit_Index_i1_LC_3_32_2 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_3_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_3_32_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_3_32_2  (
            .in0(N__14968),
            .in1(N__18180),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.rx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35352),
            .ce(N__14992),
            .sr(N__14977));
    defparam \c0.rx.equal_27_i4_2_lut_LC_3_32_3 .C_ON=1'b0;
    defparam \c0.rx.equal_27_i4_2_lut_LC_3_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_27_i4_2_lut_LC_3_32_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \c0.rx.equal_27_i4_2_lut_LC_3_32_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14941),
            .in3(N__14964),
            .lcout(n4_adj_1986),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3101_2_lut_LC_3_32_4 .C_ON=1'b0;
    defparam \c0.rx.i3101_2_lut_LC_3_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3101_2_lut_LC_3_32_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.rx.i3101_2_lut_LC_3_32_4  (
            .in0(N__14966),
            .in1(N__14939),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n3342),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_797_LC_3_32_5 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_797_LC_3_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_797_LC_3_32_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i1_2_lut_adj_797_LC_3_32_5  (
            .in0(_gnd_net_),
            .in1(N__14914),
            .in2(_gnd_net_),
            .in3(N__14883),
            .lcout(n8_adj_1996),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4002_1_lut_LC_3_32_6 .C_ON=1'b0;
    defparam \c0.tx.i4002_1_lut_LC_3_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4002_1_lut_LC_3_32_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.i4002_1_lut_LC_3_32_6  (
            .in0(N__16891),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i0_LC_4_16_0 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i0_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i0_LC_4_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i0_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__19027),
            .in2(N__15211),
            .in3(_gnd_net_),
            .lcout(\c0.delay_counter_0 ),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\c0.n4404 ),
            .clk(N__35280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i1_LC_4_16_1 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i1_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i1_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i1_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__14836),
            .in2(_gnd_net_),
            .in3(N__14824),
            .lcout(\c0.delay_counter_1 ),
            .ltout(),
            .carryin(\c0.n4404 ),
            .carryout(\c0.n4405 ),
            .clk(N__35280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i2_LC_4_16_2 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i2_LC_4_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i2_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i2_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__15223),
            .in2(_gnd_net_),
            .in3(N__14821),
            .lcout(\c0.delay_counter_2 ),
            .ltout(),
            .carryin(\c0.n4405 ),
            .carryout(\c0.n4406 ),
            .clk(N__35280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i3_LC_4_16_3 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i3_LC_4_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i3_LC_4_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i3_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__14817),
            .in2(_gnd_net_),
            .in3(N__15115),
            .lcout(\c0.delay_counter_3 ),
            .ltout(),
            .carryin(\c0.n4406 ),
            .carryout(\c0.n4407 ),
            .clk(N__35280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i4_LC_4_16_4 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i4_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i4_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i4_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__15112),
            .in2(_gnd_net_),
            .in3(N__15100),
            .lcout(\c0.delay_counter_4 ),
            .ltout(),
            .carryin(\c0.n4407 ),
            .carryout(\c0.n4408 ),
            .clk(N__35280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i5_LC_4_16_5 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i5_LC_4_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i5_LC_4_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i5_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(N__15097),
            .in2(_gnd_net_),
            .in3(N__15085),
            .lcout(\c0.delay_counter_5 ),
            .ltout(),
            .carryin(\c0.n4408 ),
            .carryout(\c0.n4409 ),
            .clk(N__35280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i6_LC_4_16_6 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i6_LC_4_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i6_LC_4_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i6_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__15081),
            .in2(_gnd_net_),
            .in3(N__15067),
            .lcout(\c0.delay_counter_6 ),
            .ltout(),
            .carryin(\c0.n4409 ),
            .carryout(\c0.n4410 ),
            .clk(N__35280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i7_LC_4_16_7 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i7_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i7_LC_4_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i7_LC_4_16_7  (
            .in0(_gnd_net_),
            .in1(N__15193),
            .in2(_gnd_net_),
            .in3(N__15064),
            .lcout(\c0.delay_counter_7 ),
            .ltout(),
            .carryin(\c0.n4410 ),
            .carryout(\c0.n4411 ),
            .clk(N__35280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i8_LC_4_17_0 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i8_LC_4_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i8_LC_4_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i8_LC_4_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15061),
            .in3(N__15046),
            .lcout(\c0.delay_counter_8 ),
            .ltout(),
            .carryin(bfn_4_17_0_),
            .carryout(\c0.n4412 ),
            .clk(N__35273),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i9_LC_4_17_1 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i9_LC_4_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i9_LC_4_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i9_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15235),
            .in3(N__15043),
            .lcout(\c0.delay_counter_9 ),
            .ltout(),
            .carryin(\c0.n4412 ),
            .carryout(\c0.n4413 ),
            .clk(N__35273),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i10_LC_4_17_2 .C_ON=1'b0;
    defparam \c0.delay_counter_528__i10_LC_4_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i10_LC_4_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i10_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(N__15037),
            .in2(_gnd_net_),
            .in3(N__15040),
            .lcout(\c0.delay_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35273),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i19_LC_4_17_3 .C_ON=1'b0;
    defparam \c0.data_out_0___i19_LC_4_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i19_LC_4_17_3 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \c0.data_out_0___i19_LC_4_17_3  (
            .in0(N__15025),
            .in1(N__16246),
            .in2(N__15004),
            .in3(N__16678),
            .lcout(data_out_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35273),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_944_LC_4_17_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_944_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_944_LC_4_17_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_944_LC_4_17_4  (
            .in0(N__16796),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16273),
            .lcout(n4_adj_2000),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_894_LC_4_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_894_LC_4_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_894_LC_4_17_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_894_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(N__16797),
            .in2(_gnd_net_),
            .in3(N__21077),
            .lcout(n5063),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5267_4_lut_LC_4_17_6 .C_ON=1'b0;
    defparam \c0.i5267_4_lut_LC_4_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5267_4_lut_LC_4_17_6 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \c0.i5267_4_lut_LC_4_17_6  (
            .in0(N__15126),
            .in1(N__20679),
            .in2(N__15250),
            .in3(N__20391),
            .lcout(\c0.n5501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_893_LC_4_17_7 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_893_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_893_LC_4_17_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_893_LC_4_17_7  (
            .in0(N__15231),
            .in1(N__15222),
            .in2(N__15210),
            .in3(N__15192),
            .lcout(\c0.n18_adj_1908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_942_LC_4_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_942_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_942_LC_4_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_942_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__16469),
            .in2(_gnd_net_),
            .in3(N__19299),
            .lcout(),
            .ltout(n5086_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i31_LC_4_18_1 .C_ON=1'b0;
    defparam \c0.data_out_0___i31_LC_4_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i31_LC_4_18_1 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \c0.data_out_0___i31_LC_4_18_1  (
            .in0(N__16669),
            .in1(N__15175),
            .in2(N__15166),
            .in3(N__20784),
            .lcout(data_out_19_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35281),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i22_LC_4_18_2 .C_ON=1'b0;
    defparam \c0.data_out_0___i22_LC_4_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i22_LC_4_18_2 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \c0.data_out_0___i22_LC_4_18_2  (
            .in0(N__16204),
            .in1(N__16198),
            .in2(N__20983),
            .in3(N__16668),
            .lcout(data_out_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35281),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_967_LC_4_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_967_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_967_LC_4_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_967_LC_4_18_3  (
            .in0(N__18806),
            .in1(N__15162),
            .in2(N__16513),
            .in3(N__16558),
            .lcout(n5156),
            .ltout(n5156_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i17_LC_4_18_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i17_LC_4_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i17_LC_4_18_4 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \c0.data_out_0___i17_LC_4_18_4  (
            .in0(N__19240),
            .in1(N__15127),
            .in2(N__15130),
            .in3(N__16667),
            .lcout(data_out_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35281),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_LC_4_18_6 .C_ON=1'b0;
    defparam \c0.i3_3_lut_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_LC_4_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_LC_4_18_6  (
            .in0(N__15376),
            .in1(N__21108),
            .in2(_gnd_net_),
            .in3(N__19298),
            .lcout(n8_adj_1997),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i32_LC_4_18_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i32_LC_4_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i32_LC_4_18_7 .LUT_INIT=16'b1110101101000001;
    LogicCell40 \c0.data_out_0___i32_LC_4_18_7  (
            .in0(N__16670),
            .in1(N__16470),
            .in2(N__15370),
            .in3(N__15342),
            .lcout(data_out_19_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35281),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5254_4_lut_4_lut_LC_4_19_1 .C_ON=1'b0;
    defparam \c0.i5254_4_lut_4_lut_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5254_4_lut_4_lut_LC_4_19_1 .LUT_INIT=16'b1101100011111111;
    LogicCell40 \c0.i5254_4_lut_4_lut_LC_4_19_1  (
            .in0(N__20409),
            .in1(N__15297),
            .in2(N__15358),
            .in3(N__20572),
            .lcout(\c0.n5519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_4_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_4_19_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_4_19_2  (
            .in0(N__15343),
            .in1(N__20407),
            .in2(_gnd_net_),
            .in3(N__15309),
            .lcout(\c0.n17_adj_1961 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i24_LC_4_19_3 .C_ON=1'b0;
    defparam \c0.data_out_0___i24_LC_4_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i24_LC_4_19_3 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \c0.data_out_0___i24_LC_4_19_3  (
            .in0(N__15310),
            .in1(N__15328),
            .in2(N__15319),
            .in3(N__16679),
            .lcout(data_out_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35286),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i28_LC_4_19_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i28_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i28_LC_4_19_4 .LUT_INIT=16'b1110010010110001;
    LogicCell40 \c0.data_out_0___i28_LC_4_19_4  (
            .in0(N__16680),
            .in1(N__15486),
            .in2(N__15301),
            .in3(N__16690),
            .lcout(data_out_19_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35286),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5227_4_lut_4_lut_LC_4_19_5 .C_ON=1'b0;
    defparam \c0.i5227_4_lut_4_lut_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5227_4_lut_4_lut_LC_4_19_5 .LUT_INIT=16'b1110010011111111;
    LogicCell40 \c0.i5227_4_lut_4_lut_LC_4_19_5  (
            .in0(N__20408),
            .in1(N__15289),
            .in2(N__16308),
            .in3(N__20571),
            .lcout(\c0.n5531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_934_LC_4_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_934_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_934_LC_4_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_934_LC_4_19_6  (
            .in0(N__20638),
            .in1(N__19296),
            .in2(_gnd_net_),
            .in3(N__16415),
            .lcout(n4_adj_2007),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n5719_bdd_4_lut_LC_4_20_0 .C_ON=1'b0;
    defparam \c0.tx.n5719_bdd_4_lut_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n5719_bdd_4_lut_LC_4_20_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.tx.n5719_bdd_4_lut_LC_4_20_0  (
            .in0(N__15265),
            .in1(N__17234),
            .in2(N__15436),
            .in3(N__17158),
            .lcout(\c0.tx.n5722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i932_4_lut_LC_4_20_2 .C_ON=1'b0;
    defparam \c0.i932_4_lut_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i932_4_lut_LC_4_20_2 .LUT_INIT=16'b1101000100100010;
    LogicCell40 \c0.i932_4_lut_LC_4_20_2  (
            .in0(N__20412),
            .in1(N__21408),
            .in2(N__15466),
            .in3(N__20580),
            .lcout(),
            .ltout(\c0.n1173_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_4_20_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_4_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_4_20_3 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_4_20_3  (
            .in0(N__21189),
            .in1(N__15451),
            .in2(N__15442),
            .in3(N__21313),
            .lcout(),
            .ltout(tx_data_0_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_4_20_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_4_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_4_20_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_4_20_4  (
            .in0(N__15435),
            .in1(_gnd_net_),
            .in2(N__15439),
            .in3(N__19341),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35292),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_4_lut_LC_4_20_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_4_lut_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_4_lut_LC_4_20_5 .LUT_INIT=16'b0110010010011001;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_4_lut_LC_4_20_5  (
            .in0(N__21407),
            .in1(N__21312),
            .in2(N__16765),
            .in3(N__20579),
            .lcout(),
            .ltout(\c0.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_4_20_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_4_20_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_4_20_6  (
            .in0(N__21230),
            .in1(N__15424),
            .in2(N__15418),
            .in3(N__21188),
            .lcout(tx_data_1_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_4_21_1 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_4_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_4_21_1 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_4_21_1  (
            .in0(N__15676),
            .in1(N__17237),
            .in2(N__17191),
            .in3(N__15666),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35297),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_4_21_2 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_4_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_4_21_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_4_21_2  (
            .in0(N__15665),
            .in1(N__17186),
            .in2(_gnd_net_),
            .in3(N__15675),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35297),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_adj_799_LC_4_21_3 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_adj_799_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_adj_799_LC_4_21_3 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \c0.tx.i1_4_lut_adj_799_LC_4_21_3  (
            .in0(N__17050),
            .in1(N__17099),
            .in2(N__16983),
            .in3(N__15402),
            .lcout(n2200),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_3_lut_LC_4_21_4 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_3_lut_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_3_lut_LC_4_21_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i2_2_lut_3_lut_LC_4_21_4  (
            .in0(N__17150),
            .in1(N__17235),
            .in2(_gnd_net_),
            .in3(N__17185),
            .lcout(\c0.tx.n3507 ),
            .ltout(\c0.tx.n3507_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2063_3_lut_LC_4_21_5 .C_ON=1'b0;
    defparam \c0.tx.i2063_3_lut_LC_4_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2063_3_lut_LC_4_21_5 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \c0.tx.i2063_3_lut_LC_4_21_5  (
            .in0(_gnd_net_),
            .in1(N__17100),
            .in2(N__15679),
            .in3(N__15664),
            .lcout(n2307),
            .ltout(n2307_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_4_21_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_4_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_4_21_6 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_4_21_6  (
            .in0(N__15667),
            .in1(N__15649),
            .in2(N__15652),
            .in3(N__17152),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35297),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i573_2_lut_LC_4_22_1 .C_ON=1'b0;
    defparam \c0.tx.i573_2_lut_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i573_2_lut_LC_4_22_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx.i573_2_lut_LC_4_22_1  (
            .in0(_gnd_net_),
            .in1(N__17236),
            .in2(_gnd_net_),
            .in3(N__17190),
            .lcout(n805),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i1_LC_4_22_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i1_LC_4_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i1_LC_4_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.tx2.r_Bit_Index_i1_LC_4_22_3  (
            .in0(_gnd_net_),
            .in1(N__15572),
            .in2(_gnd_net_),
            .in3(N__15639),
            .lcout(\c0.tx2.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35302),
            .ce(N__15508),
            .sr(N__15499));
    defparam \c0.tx2.r_Bit_Index_i2_LC_4_22_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i2_LC_4_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i2_LC_4_22_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \c0.tx2.r_Bit_Index_i2_LC_4_22_4  (
            .in0(N__15640),
            .in1(_gnd_net_),
            .in2(N__15590),
            .in3(N__15530),
            .lcout(\c0.tx2.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35302),
            .ce(N__15508),
            .sr(N__15499));
    defparam \c0.i1_2_lut_adj_847_LC_4_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_847_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_847_LC_4_22_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_847_LC_4_22_6  (
            .in0(_gnd_net_),
            .in1(N__20471),
            .in2(_gnd_net_),
            .in3(N__21123),
            .lcout(n5153),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3173_2_lut_LC_4_24_0 .C_ON=1'b0;
    defparam \c0.i3173_2_lut_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3173_2_lut_LC_4_24_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i3173_2_lut_LC_4_24_0  (
            .in0(_gnd_net_),
            .in1(N__15756),
            .in2(_gnd_net_),
            .in3(N__15781),
            .lcout(\c0.n3414 ),
            .ltout(\c0.n3414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_1801_LC_4_24_1 .C_ON=1'b0;
    defparam \c0.tx2_transmit_1801_LC_4_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2_transmit_1801_LC_4_24_1 .LUT_INIT=16'b0000100001011101;
    LogicCell40 \c0.tx2_transmit_1801_LC_4_24_1  (
            .in0(N__36482),
            .in1(N__15822),
            .in2(N__15469),
            .in3(N__17320),
            .lcout(\c0.r_SM_Main_2_N_1770_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5430_LC_4_24_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5430_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5430_LC_4_24_2 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5430_LC_4_24_2  (
            .in0(N__33138),
            .in1(N__26101),
            .in2(N__32506),
            .in3(N__31348),
            .lcout(\c0.n5791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_4_24_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_4_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_4_24_3 .LUT_INIT=16'b1110000011101111;
    LogicCell40 \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_4_24_3  (
            .in0(N__15829),
            .in1(N__15821),
            .in2(N__36636),
            .in3(N__17319),
            .lcout(\c0.FRAME_MATCHER_wait_for_transmission ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i489_3_lut_4_lut_LC_4_24_5 .C_ON=1'b0;
    defparam \c0.i489_3_lut_4_lut_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i489_3_lut_4_lut_LC_4_24_5 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \c0.i489_3_lut_4_lut_LC_4_24_5  (
            .in0(N__15780),
            .in1(N__15757),
            .in2(N__36635),
            .in3(N__17318),
            .lcout(\c0.n195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5475_LC_4_24_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5475_LC_4_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5475_LC_4_24_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5475_LC_4_24_6  (
            .in0(N__33139),
            .in1(N__28024),
            .in2(N__32507),
            .in3(N__31069),
            .lcout(),
            .ltout(\c0.n5845_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5845_bdd_4_lut_LC_4_24_7 .C_ON=1'b0;
    defparam \c0.n5845_bdd_4_lut_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.n5845_bdd_4_lut_LC_4_24_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5845_bdd_4_lut_LC_4_24_7  (
            .in0(N__32315),
            .in1(N__31585),
            .in2(N__15724),
            .in3(N__21997),
            .lcout(\c0.n5411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i118_LC_4_25_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i118_LC_4_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i118_LC_4_25_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i118_LC_4_25_0  (
            .in0(N__34075),
            .in1(N__20218),
            .in2(_gnd_net_),
            .in3(N__19433),
            .lcout(data_in_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35316),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5293_2_lut_LC_4_25_1 .C_ON=1'b0;
    defparam \c0.i5293_2_lut_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5293_2_lut_LC_4_25_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \c0.i5293_2_lut_LC_4_25_1  (
            .in0(N__36437),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17317),
            .lcout(\c0.n2275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_810_LC_4_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_810_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_810_LC_4_25_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_810_LC_4_25_2  (
            .in0(_gnd_net_),
            .in1(N__23432),
            .in2(_gnd_net_),
            .in3(N__15709),
            .lcout(\c0.n1918 ),
            .ltout(\c0.n1918_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_995_LC_4_25_3 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_995_LC_4_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_995_LC_4_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_995_LC_4_25_3  (
            .in0(N__22622),
            .in1(N__17754),
            .in2(N__15685),
            .in3(N__31954),
            .lcout(\c0.n5192 ),
            .ltout(\c0.n5192_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_3_lut_adj_881_LC_4_25_4 .C_ON=1'b0;
    defparam \c0.i9_3_lut_adj_881_LC_4_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_3_lut_adj_881_LC_4_25_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i9_3_lut_adj_881_LC_4_25_4  (
            .in0(_gnd_net_),
            .in1(N__23750),
            .in2(N__15682),
            .in3(N__23372),
            .lcout(),
            .ltout(\c0.n30_adj_1897_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_923_LC_4_25_5 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_923_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_923_LC_4_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_923_LC_4_25_5  (
            .in0(N__17578),
            .in1(N__25774),
            .in2(N__15919),
            .in3(N__25809),
            .lcout(),
            .ltout(\c0.n36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_LC_4_25_6 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_4_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_LC_4_25_6  (
            .in0(N__26284),
            .in1(N__19387),
            .in2(N__15916),
            .in3(N__22009),
            .lcout(\c0.n5277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_917_LC_4_26_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_917_LC_4_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_917_LC_4_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_917_LC_4_26_0  (
            .in0(N__15910),
            .in1(N__21624),
            .in2(N__26113),
            .in3(N__30511),
            .lcout(\c0.n21_adj_1928 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_4_26_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_4_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_4_26_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_4_26_1  (
            .in0(N__25885),
            .in1(N__25381),
            .in2(N__23023),
            .in3(N__24081),
            .lcout(\c0.n5080 ),
            .ltout(\c0.n5080_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_911_LC_4_26_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_911_LC_4_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_911_LC_4_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_911_LC_4_26_2  (
            .in0(N__29890),
            .in1(N__19669),
            .in2(N__15913),
            .in3(N__21993),
            .lcout(\c0.n24_adj_1924 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_853_LC_4_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_853_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_853_LC_4_26_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_853_LC_4_26_3  (
            .in0(_gnd_net_),
            .in1(N__32913),
            .in2(_gnd_net_),
            .in3(N__22830),
            .lcout(\c0.n1990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_916_LC_4_26_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_916_LC_4_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_916_LC_4_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_916_LC_4_26_4  (
            .in0(N__24913),
            .in1(N__15904),
            .in2(N__30267),
            .in3(N__15895),
            .lcout(),
            .ltout(\c0.n22_adj_1927_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_921_LC_4_26_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_921_LC_4_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_921_LC_4_26_5 .LUT_INIT=16'b1111111110010110;
    LogicCell40 \c0.i7_4_lut_adj_921_LC_4_26_5  (
            .in0(N__15889),
            .in1(N__15883),
            .in2(N__15877),
            .in3(N__15973),
            .lcout(\c0.n23_adj_1932 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_904_LC_4_27_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_904_LC_4_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_904_LC_4_27_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_904_LC_4_27_0  (
            .in0(N__15874),
            .in1(N__24580),
            .in2(N__15865),
            .in3(N__27225),
            .lcout(\c0.n27_adj_1919 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i72_LC_4_27_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i72_LC_4_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i72_LC_4_27_1 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i72_LC_4_27_1  (
            .in0(N__36058),
            .in1(N__22468),
            .in2(N__36650),
            .in3(N__17499),
            .lcout(\c0.data_in_field_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i83_LC_4_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i83_LC_4_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i83_LC_4_27_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i83_LC_4_27_2  (
            .in0(N__22769),
            .in1(N__36501),
            .in2(N__31639),
            .in3(N__36061),
            .lcout(\c0.data_in_field_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i145_LC_4_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i145_LC_4_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i145_LC_4_27_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0___i145_LC_4_27_3  (
            .in0(N__36057),
            .in1(N__16011),
            .in2(N__36649),
            .in3(N__33477),
            .lcout(\c0.data_in_frame_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i100_LC_4_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i100_LC_4_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i100_LC_4_27_4 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i100_LC_4_27_4  (
            .in0(N__21581),
            .in1(N__36500),
            .in2(N__31840),
            .in3(N__36060),
            .lcout(\c0.data_in_field_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_851_LC_4_27_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_851_LC_4_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_851_LC_4_27_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_851_LC_4_27_5  (
            .in0(_gnd_net_),
            .in1(N__21580),
            .in2(_gnd_net_),
            .in3(N__22768),
            .lcout(\c0.n5225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i149_LC_4_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i149_LC_4_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i149_LC_4_27_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i149_LC_4_27_6  (
            .in0(N__15993),
            .in1(N__36059),
            .in2(N__26808),
            .in3(N__36508),
            .lcout(\c0.data_in_frame_18_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_918_LC_4_27_7 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_918_LC_4_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_918_LC_4_27_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_918_LC_4_27_7  (
            .in0(N__15979),
            .in1(N__22078),
            .in2(N__17896),
            .in3(N__15925),
            .lcout(\c0.n5266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i104_LC_4_28_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i104_LC_4_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i104_LC_4_28_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i104_LC_4_28_0  (
            .in0(N__34074),
            .in1(N__24779),
            .in2(_gnd_net_),
            .in3(N__25725),
            .lcout(data_in_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35331),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_4_lut_LC_4_28_1 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_4_lut_LC_4_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_4_lut_LC_4_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_2_lut_3_lut_4_lut_LC_4_28_1  (
            .in0(N__32990),
            .in1(N__29367),
            .in2(N__24757),
            .in3(N__22946),
            .lcout(),
            .ltout(\c0.n18_adj_1882_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_866_LC_4_28_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_866_LC_4_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_866_LC_4_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_866_LC_4_28_2  (
            .in0(N__24709),
            .in1(N__15959),
            .in2(N__15928),
            .in3(N__25018),
            .lcout(\c0.n26_adj_1883 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_120_2_lut_3_lut_4_lut_LC_4_28_3 .C_ON=1'b0;
    defparam \c0.i1_rep_120_2_lut_3_lut_4_lut_LC_4_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_120_2_lut_3_lut_4_lut_LC_4_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_rep_120_2_lut_3_lut_4_lut_LC_4_28_3  (
            .in0(N__22823),
            .in1(N__32985),
            .in2(N__32914),
            .in3(N__29366),
            .lcout(\c0.n6103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i87_LC_4_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i87_LC_4_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i87_LC_4_28_4 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i87_LC_4_28_4  (
            .in0(N__29977),
            .in1(N__36011),
            .in2(N__32994),
            .in3(N__36638),
            .lcout(\c0.data_in_field_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35331),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_859_LC_4_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_859_LC_4_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_859_LC_4_28_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_859_LC_4_28_5  (
            .in0(_gnd_net_),
            .in1(N__21733),
            .in2(_gnd_net_),
            .in3(N__32986),
            .lcout(\c0.n5201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i31_LC_4_28_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i31_LC_4_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i31_LC_4_28_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i31_LC_4_28_6  (
            .in0(N__21734),
            .in1(N__36637),
            .in2(N__27850),
            .in3(N__36012),
            .lcout(\c0.data_in_field_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35331),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i110_LC_4_28_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i110_LC_4_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i110_LC_4_28_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i110_LC_4_28_7  (
            .in0(N__34218),
            .in1(N__19440),
            .in2(_gnd_net_),
            .in3(N__17594),
            .lcout(data_in_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35331),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5731_bdd_4_lut_LC_4_29_0 .C_ON=1'b0;
    defparam \c0.n5731_bdd_4_lut_LC_4_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.n5731_bdd_4_lut_LC_4_29_0 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n5731_bdd_4_lut_LC_4_29_0  (
            .in0(N__21947),
            .in1(N__32791),
            .in2(N__17905),
            .in3(N__29800),
            .lcout(\c0.n5462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i102_LC_4_29_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i102_LC_4_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i102_LC_4_29_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i102_LC_4_29_1  (
            .in0(N__17595),
            .in1(N__34073),
            .in2(_gnd_net_),
            .in3(N__16029),
            .lcout(data_in_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i84_LC_4_29_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i84_LC_4_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i84_LC_4_29_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i84_LC_4_29_2  (
            .in0(N__35991),
            .in1(N__37127),
            .in2(N__26473),
            .in3(N__23422),
            .lcout(\c0.data_in_field_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i106_LC_4_29_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i106_LC_4_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i106_LC_4_29_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i106_LC_4_29_3  (
            .in0(N__37126),
            .in1(N__35992),
            .in2(N__21954),
            .in3(N__30979),
            .lcout(\c0.data_in_field_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i121_LC_4_29_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i121_LC_4_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i121_LC_4_29_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i121_LC_4_29_4  (
            .in0(N__23468),
            .in1(N__19629),
            .in2(N__36196),
            .in3(N__37128),
            .lcout(\c0.data_in_field_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_986_LC_4_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_986_LC_4_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_986_LC_4_29_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_986_LC_4_29_5  (
            .in0(N__22161),
            .in1(N__21946),
            .in2(_gnd_net_),
            .in3(N__23467),
            .lcout(\c0.n5222 ),
            .ltout(\c0.n5222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_3_lut_LC_4_29_6 .C_ON=1'b0;
    defparam \c0.i9_3_lut_LC_4_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_3_lut_LC_4_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i9_3_lut_LC_4_29_6  (
            .in0(_gnd_net_),
            .in1(N__17506),
            .in2(N__16069),
            .in3(N__21882),
            .lcout(),
            .ltout(\c0.n33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_LC_4_29_7 .C_ON=1'b0;
    defparam \c0.i21_4_lut_LC_4_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_LC_4_29_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_LC_4_29_7  (
            .in0(N__28333),
            .in1(N__16066),
            .in2(N__16060),
            .in3(N__25414),
            .lcout(\c0.n45_adj_1885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i96_LC_4_30_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i96_LC_4_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i96_LC_4_30_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i96_LC_4_30_0  (
            .in0(N__24789),
            .in1(N__34082),
            .in2(_gnd_net_),
            .in3(N__22721),
            .lcout(data_in_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35346),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i152_LC_4_30_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i152_LC_4_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i152_LC_4_30_1 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \c0.data_in_0___i152_LC_4_30_1  (
            .in0(N__26039),
            .in1(N__20159),
            .in2(N__34284),
            .in3(_gnd_net_),
            .lcout(data_in_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35346),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_825_LC_4_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_825_LC_4_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_825_LC_4_30_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_825_LC_4_30_2  (
            .in0(_gnd_net_),
            .in1(N__20185),
            .in2(_gnd_net_),
            .in3(N__24841),
            .lcout(\c0.n2008 ),
            .ltout(\c0.n2008_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_867_LC_4_30_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_867_LC_4_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_867_LC_4_30_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_867_LC_4_30_3  (
            .in0(N__24635),
            .in1(N__23553),
            .in2(N__16057),
            .in3(N__22870),
            .lcout(),
            .ltout(\c0.n38_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_4_30_4 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_4_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_4_30_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_LC_4_30_4  (
            .in0(N__24853),
            .in1(N__26038),
            .in2(N__16054),
            .in3(N__26264),
            .lcout(\c0.n43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i112_LC_4_30_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i112_LC_4_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i112_LC_4_30_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i112_LC_4_30_5  (
            .in0(N__34076),
            .in1(N__21663),
            .in2(_gnd_net_),
            .in3(N__25718),
            .lcout(data_in_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35346),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i121_LC_4_30_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i121_LC_4_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i121_LC_4_30_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i121_LC_4_30_6  (
            .in0(N__27613),
            .in1(N__34081),
            .in2(_gnd_net_),
            .in3(N__19614),
            .lcout(data_in_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35346),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i159_LC_4_30_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i159_LC_4_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i159_LC_4_30_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i159_LC_4_30_7  (
            .in0(N__34077),
            .in1(N__16084),
            .in2(_gnd_net_),
            .in3(N__17360),
            .lcout(data_in_19_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35346),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_124_2_lut_LC_4_31_0 .C_ON=1'b0;
    defparam \c0.i1_rep_124_2_lut_LC_4_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_124_2_lut_LC_4_31_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_rep_124_2_lut_LC_4_31_0  (
            .in0(_gnd_net_),
            .in1(N__28789),
            .in2(_gnd_net_),
            .in3(N__20042),
            .lcout(\c0.n6107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i14_LC_4_31_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i14_LC_4_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i14_LC_4_31_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i14_LC_4_31_1  (
            .in0(N__34035),
            .in1(N__16103),
            .in2(_gnd_net_),
            .in3(N__24146),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35353),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i151_LC_4_31_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i151_LC_4_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i151_LC_4_31_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i151_LC_4_31_2  (
            .in0(N__16125),
            .in1(N__24212),
            .in2(N__36193),
            .in3(N__36639),
            .lcout(\c0.data_in_frame_18_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35353),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_949_LC_4_31_3 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_949_LC_4_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_949_LC_4_31_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10_4_lut_adj_949_LC_4_31_3  (
            .in0(N__31730),
            .in1(N__16102),
            .in2(N__31440),
            .in3(N__17836),
            .lcout(\c0.n26_adj_1955 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i62_LC_4_31_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i62_LC_4_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i62_LC_4_31_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i62_LC_4_31_5  (
            .in0(N__34036),
            .in1(N__22497),
            .in2(_gnd_net_),
            .in3(N__24234),
            .lcout(data_in_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35353),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i157_LC_4_31_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i157_LC_4_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i157_LC_4_31_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i157_LC_4_31_6  (
            .in0(N__16156),
            .in1(N__34037),
            .in2(_gnd_net_),
            .in3(N__37315),
            .lcout(data_in_19_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35353),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_4_32_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_4_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_4_32_0 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_4_32_0  (
            .in0(N__16080),
            .in1(N__20935),
            .in2(N__17953),
            .in3(N__20835),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i72_LC_4_32_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i72_LC_4_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i72_LC_4_32_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i72_LC_4_32_1  (
            .in0(N__23845),
            .in1(N__33874),
            .in2(_gnd_net_),
            .in3(N__22457),
            .lcout(data_in_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i16_LC_4_32_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i16_LC_4_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i16_LC_4_32_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i16_LC_4_32_2  (
            .in0(N__33872),
            .in1(N__22671),
            .in2(_gnd_net_),
            .in3(N__27577),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13_4_lut_4_lut_LC_4_32_3 .C_ON=1'b0;
    defparam \c0.rx.i13_4_lut_4_lut_LC_4_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13_4_lut_4_lut_LC_4_32_3 .LUT_INIT=16'b0001100100010001;
    LogicCell40 \c0.rx.i13_4_lut_4_lut_LC_4_32_3  (
            .in0(N__18136),
            .in1(N__18278),
            .in2(N__18364),
            .in3(N__18066),
            .lcout(),
            .ltout(\c0.rx.n2151_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_4_32_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_4_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_4_32_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_4_32_4  (
            .in0(N__33873),
            .in1(N__18279),
            .in2(N__16177),
            .in3(N__18361),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_4_lut_4_lut_adj_792_LC_4_32_5 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_4_lut_4_lut_adj_792_LC_4_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_4_lut_4_lut_adj_792_LC_4_32_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.rx.i1_2_lut_4_lut_4_lut_adj_792_LC_4_32_5  (
            .in0(N__18179),
            .in1(N__18190),
            .in2(N__18139),
            .in3(N__18065),
            .lcout(n1709),
            .ltout(n1709_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_4_32_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_4_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_4_32_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_4_32_6  (
            .in0(N__20933),
            .in1(N__16155),
            .in2(N__16174),
            .in3(N__16171),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_4_32_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_4_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_4_32_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_4_32_7  (
            .in0(N__18015),
            .in1(N__17948),
            .in2(N__21480),
            .in3(N__20934),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i8_LC_5_16_2 .C_ON=1'b0;
    defparam \c0.data_out_0___i8_LC_5_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i8_LC_5_16_2 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i8_LC_5_16_2  (
            .in0(N__16354),
            .in1(N__19207),
            .in2(N__18508),
            .in3(N__19078),
            .lcout(data_out_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35287),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_973_LC_5_16_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_973_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_973_LC_5_16_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_973_LC_5_16_3  (
            .in0(N__20468),
            .in1(N__20748),
            .in2(N__18813),
            .in3(N__16582),
            .lcout(n4_adj_1992),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i972_2_lut_LC_5_16_5 .C_ON=1'b0;
    defparam \c0.i972_2_lut_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i972_2_lut_LC_5_16_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i972_2_lut_LC_5_16_5  (
            .in0(_gnd_net_),
            .in1(N__21318),
            .in2(_gnd_net_),
            .in3(N__20586),
            .lcout(\c0.n1227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2006_4_lut_LC_5_17_1 .C_ON=1'b0;
    defparam \c0.i2006_4_lut_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2006_4_lut_LC_5_17_1 .LUT_INIT=16'b1100000010111011;
    LogicCell40 \c0.i2006_4_lut_LC_5_17_1  (
            .in0(N__18976),
            .in1(N__21417),
            .in2(N__16514),
            .in3(N__20403),
            .lcout(\c0.n2249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i11_LC_5_17_2 .C_ON=1'b0;
    defparam \c0.data_out_0___i11_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i11_LC_5_17_2 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i11_LC_5_17_2  (
            .in0(N__16512),
            .in1(N__19221),
            .in2(N__18448),
            .in3(N__19056),
            .lcout(data_out_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35277),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_971_LC_5_17_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_971_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_971_LC_5_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_971_LC_5_17_3  (
            .in0(N__16809),
            .in1(N__16344),
            .in2(N__16515),
            .in3(N__16271),
            .lcout(n5135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i9_LC_5_17_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i9_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i9_LC_5_17_4 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i9_LC_5_17_4  (
            .in0(N__16272),
            .in1(N__19222),
            .in2(N__18490),
            .in3(N__19057),
            .lcout(data_out_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35277),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5249_4_lut_LC_5_17_5 .C_ON=1'b0;
    defparam \c0.i5249_4_lut_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5249_4_lut_LC_5_17_5 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \c0.i5249_4_lut_LC_5_17_5  (
            .in0(N__16245),
            .in1(N__20678),
            .in2(N__16234),
            .in3(N__20404),
            .lcout(),
            .ltout(\c0.n5522_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_5_17_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_5_17_6 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_5_17_6  (
            .in0(N__18657),
            .in1(N__16213),
            .in2(N__16207),
            .in3(N__21187),
            .lcout(tx_data_2_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_845_LC_5_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_845_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_845_LC_5_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_845_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(N__16363),
            .in2(_gnd_net_),
            .in3(N__16435),
            .lcout(n4_adj_1991),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5257_4_lut_LC_5_18_1 .C_ON=1'b0;
    defparam \c0.i5257_4_lut_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5257_4_lut_LC_5_18_1 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \c0.i5257_4_lut_LC_5_18_1  (
            .in0(N__16197),
            .in1(N__20677),
            .in2(N__16600),
            .in3(N__20413),
            .lcout(\c0.n5489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_940_LC_5_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_940_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_940_LC_5_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_940_LC_5_18_2  (
            .in0(N__16703),
            .in1(N__18748),
            .in2(_gnd_net_),
            .in3(N__16580),
            .lcout(n4_adj_1994),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_941_LC_5_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_941_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_941_LC_5_18_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_941_LC_5_18_4  (
            .in0(N__18792),
            .in1(_gnd_net_),
            .in2(N__16710),
            .in3(N__16581),
            .lcout(n5117),
            .ltout(n5117_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i30_LC_5_18_5 .C_ON=1'b0;
    defparam \c0.data_out_0___i30_LC_5_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i30_LC_5_18_5 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \c0.data_out_0___i30_LC_5_18_5  (
            .in0(N__16599),
            .in1(N__20692),
            .in2(N__16684),
            .in3(N__16681),
            .lcout(data_out_19_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35288),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_5_18_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_5_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_5_18_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_5_18_6  (
            .in0(N__19368),
            .in1(N__16588),
            .in2(_gnd_net_),
            .in3(N__17256),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35288),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_936_LC_5_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_936_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_936_LC_5_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_936_LC_5_19_0  (
            .in0(N__18781),
            .in1(N__20744),
            .in2(_gnd_net_),
            .in3(N__16579),
            .lcout(\c0.n1805 ),
            .ltout(\c0.n1805_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_965_LC_5_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_965_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_965_LC_5_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_965_LC_5_19_1  (
            .in0(N__16519),
            .in1(N__20641),
            .in2(N__16477),
            .in3(N__16433),
            .lcout(n135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_5_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_5_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_5_19_2  (
            .in0(N__21119),
            .in1(N__20743),
            .in2(_gnd_net_),
            .in3(N__20410),
            .lcout(\c0.n9_adj_1890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_933_LC_5_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_933_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_933_LC_5_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_933_LC_5_19_3  (
            .in0(N__16450),
            .in1(N__20642),
            .in2(_gnd_net_),
            .in3(N__16434),
            .lcout(n5173),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2004_4_lut_LC_5_19_4 .C_ON=1'b0;
    defparam \c0.i2004_4_lut_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2004_4_lut_LC_5_19_4 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \c0.i2004_4_lut_LC_5_19_4  (
            .in0(N__16432),
            .in1(N__21415),
            .in2(N__16370),
            .in3(N__20411),
            .lcout(\c0.n2247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i26_LC_5_19_5 .C_ON=1'b0;
    defparam \c0.data_out_0___i26_LC_5_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i26_LC_5_19_5 .LUT_INIT=16'b1011000111110000;
    LogicCell40 \c0.data_out_0___i26_LC_5_19_5  (
            .in0(N__19208),
            .in1(N__16318),
            .in2(N__16309),
            .in3(N__19079),
            .lcout(data_out_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_5_19_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_5_19_6 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_5_19_6  (
            .in0(N__16849),
            .in1(N__16843),
            .in2(N__21238),
            .in3(N__21190),
            .lcout(tx_data_3_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_5365_LC_5_20_1 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_5365_LC_5_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_5365_LC_5_20_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx.r_Bit_Index_0__bdd_4_lut_5365_LC_5_20_1  (
            .in0(N__18639),
            .in1(N__19311),
            .in2(N__17242),
            .in3(N__17184),
            .lcout(),
            .ltout(\c0.tx.n5713_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n5713_bdd_4_lut_LC_5_20_2 .C_ON=1'b0;
    defparam \c0.tx.n5713_bdd_4_lut_LC_5_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n5713_bdd_4_lut_LC_5_20_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.tx.n5713_bdd_4_lut_LC_5_20_2  (
            .in0(N__17233),
            .in1(N__16831),
            .in2(N__16813),
            .in3(N__16728),
            .lcout(\c0.tx.n5716 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_5_20_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_5_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_5_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_5_20_3  (
            .in0(N__16808),
            .in1(N__21044),
            .in2(_gnd_net_),
            .in3(N__20405),
            .lcout(\c0.n9_adj_1880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i750_4_lut_LC_5_20_4 .C_ON=1'b0;
    defparam \c0.i750_4_lut_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i750_4_lut_LC_5_20_4 .LUT_INIT=16'b1101000100100010;
    LogicCell40 \c0.i750_4_lut_LC_5_20_4  (
            .in0(N__20406),
            .in1(N__21416),
            .in2(N__16756),
            .in3(N__20587),
            .lcout(),
            .ltout(\c0.n991_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_5_20_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_5_20_5 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_5_20_5  (
            .in0(N__21191),
            .in1(N__16744),
            .in2(N__16735),
            .in3(N__21314),
            .lcout(),
            .ltout(tx_data_5_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_5_20_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_5_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_5_20_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_5_20_6  (
            .in0(_gnd_net_),
            .in1(N__19369),
            .in2(N__16732),
            .in3(N__16729),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35298),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i2_LC_5_21_1 .C_ON=1'b0;
    defparam \c0.data_out_0___i2_LC_5_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i2_LC_5_21_1 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i2_LC_5_21_1  (
            .in0(N__21059),
            .in1(N__19224),
            .in2(N__18601),
            .in3(N__19083),
            .lcout(data_out_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35303),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_5_21_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_5_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_5_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_5_21_3  (
            .in0(N__19370),
            .in1(N__16720),
            .in2(_gnd_net_),
            .in3(N__17266),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35303),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_21_4 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_21_4 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_5_21_4  (
            .in0(N__17265),
            .in1(N__17257),
            .in2(N__17238),
            .in3(N__17183),
            .lcout(\c0.tx.n5719 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i342127_i1_3_lut_LC_5_21_5 .C_ON=1'b0;
    defparam \c0.tx.i342127_i1_3_lut_LC_5_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i342127_i1_3_lut_LC_5_21_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.i342127_i1_3_lut_LC_5_21_5  (
            .in0(N__17151),
            .in1(N__17134),
            .in2(_gnd_net_),
            .in3(N__17128),
            .lcout(),
            .ltout(\c0.tx.o_Tx_Serial_N_1798_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_21_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_21_6 .LUT_INIT=16'b1100110011110011;
    LogicCell40 \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_5_21_6  (
            .in0(_gnd_net_),
            .in1(N__17117),
            .in2(N__17065),
            .in3(N__17061),
            .lcout(),
            .ltout(\c0.tx.n3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_5_21_7 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_5_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_5_21_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_5_21_7  (
            .in0(N__16992),
            .in1(_gnd_net_),
            .in2(N__16894),
            .in3(N__16869),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35303),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_811_LC_5_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_811_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_811_LC_5_23_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_811_LC_5_23_0  (
            .in0(_gnd_net_),
            .in1(N__29030),
            .in2(_gnd_net_),
            .in3(N__25998),
            .lcout(\c0.n2018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_870_LC_5_24_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_870_LC_5_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_870_LC_5_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_870_LC_5_24_1  (
            .in0(N__19746),
            .in1(N__29534),
            .in2(N__16858),
            .in3(N__23757),
            .lcout(\c0.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i147_LC_5_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i147_LC_5_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i147_LC_5_24_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i147_LC_5_24_2  (
            .in0(N__17398),
            .in1(N__36496),
            .in2(N__31251),
            .in3(N__36321),
            .lcout(\c0.data_in_frame_18_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_857_LC_5_24_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_857_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_857_LC_5_24_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_857_LC_5_24_3  (
            .in0(_gnd_net_),
            .in1(N__30381),
            .in2(_gnd_net_),
            .in3(N__30849),
            .lcout(\c0.n5147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i108_LC_5_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i108_LC_5_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i108_LC_5_24_4 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i108_LC_5_24_4  (
            .in0(N__30382),
            .in1(N__36494),
            .in2(N__31870),
            .in3(N__36319),
            .lcout(\c0.data_in_field_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i130_LC_5_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i130_LC_5_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i130_LC_5_24_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i130_LC_5_24_6  (
            .in0(N__30850),
            .in1(N__36495),
            .in2(N__30223),
            .in3(N__36320),
            .lcout(\c0.data_in_field_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5573_LC_5_24_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5573_LC_5_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5573_LC_5_24_7 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5573_LC_5_24_7  (
            .in0(N__17397),
            .in1(N__32412),
            .in2(N__18889),
            .in3(N__33212),
            .lcout(\c0.n5965 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_885_LC_5_25_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_885_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_885_LC_5_25_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_885_LC_5_25_0  (
            .in0(N__19378),
            .in1(N__28029),
            .in2(N__17371),
            .in3(N__28756),
            .lcout(),
            .ltout(\c0.n22_adj_1901_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_928_LC_5_25_1 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_928_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_928_LC_5_25_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_928_LC_5_25_1  (
            .in0(N__19951),
            .in1(N__23179),
            .in2(N__17332),
            .in3(N__34684),
            .lcout(\c0.n5280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_931_LC_5_25_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_931_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_931_LC_5_25_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_931_LC_5_25_2  (
            .in0(N__17635),
            .in1(N__17329),
            .in2(N__19549),
            .in3(N__17776),
            .lcout(),
            .ltout(\c0.n30_adj_1940_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3321_4_lut_LC_5_25_3 .C_ON=1'b0;
    defparam \c0.i3321_4_lut_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3321_4_lut_LC_5_25_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3321_4_lut_LC_5_25_3  (
            .in0(N__35838),
            .in1(N__17290),
            .in2(N__17323),
            .in3(N__17446),
            .lcout(\c0.n3563 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_932_LC_5_25_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_932_LC_5_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_932_LC_5_25_4 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \c0.i9_4_lut_adj_932_LC_5_25_4  (
            .in0(N__19690),
            .in1(N__17302),
            .in2(N__19402),
            .in3(N__17296),
            .lcout(\c0.n25_adj_1941 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_900_LC_5_26_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_900_LC_5_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_900_LC_5_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_900_LC_5_26_0  (
            .in0(N__23335),
            .in1(N__17284),
            .in2(N__17626),
            .in3(N__17695),
            .lcout(),
            .ltout(\c0.n26_adj_1915_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_903_LC_5_26_1 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_903_LC_5_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_903_LC_5_26_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_903_LC_5_26_1  (
            .in0(N__19603),
            .in1(N__24484),
            .in2(N__17542),
            .in3(N__22441),
            .lcout(\c0.n5250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i140_LC_5_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i140_LC_5_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i140_LC_5_26_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i140_LC_5_26_2  (
            .in0(N__17539),
            .in1(N__36314),
            .in2(N__25008),
            .in3(N__36509),
            .lcout(\c0.data_in_field_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_3_lut_LC_5_26_3 .C_ON=1'b0;
    defparam \c0.i11_3_lut_LC_5_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11_3_lut_LC_5_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i11_3_lut_LC_5_26_3  (
            .in0(N__19602),
            .in1(N__22522),
            .in2(_gnd_net_),
            .in3(N__17608),
            .lcout(),
            .ltout(\c0.n26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_901_LC_5_26_4 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_901_LC_5_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_901_LC_5_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_901_LC_5_26_4  (
            .in0(N__30316),
            .in1(N__17507),
            .in2(N__17464),
            .in3(N__22315),
            .lcout(),
            .ltout(\c0.n28_adj_1917_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_930_LC_5_26_5 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_930_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_930_LC_5_26_5 .LUT_INIT=16'b1111111111101101;
    LogicCell40 \c0.i10_4_lut_adj_930_LC_5_26_5  (
            .in0(N__17461),
            .in1(N__17455),
            .in2(N__17449),
            .in3(N__19717),
            .lcout(\c0.n26_adj_1939 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_886_LC_5_27_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_886_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_886_LC_5_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_886_LC_5_27_1  (
            .in0(N__17440),
            .in1(N__31203),
            .in2(N__17877),
            .in3(N__25161),
            .lcout(\c0.n28_adj_1902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i127_LC_5_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i127_LC_5_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i127_LC_5_27_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i127_LC_5_27_2  (
            .in0(N__23692),
            .in1(N__36315),
            .in2(N__33360),
            .in3(N__36951),
            .lcout(\c0.data_in_field_126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i135_LC_5_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i135_LC_5_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i135_LC_5_27_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0___i135_LC_5_27_3  (
            .in0(N__36950),
            .in1(N__19680),
            .in2(N__36330),
            .in3(N__17935),
            .lcout(\c0.data_in_field_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_873_LC_5_27_4 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_873_LC_5_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_873_LC_5_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_873_LC_5_27_4  (
            .in0(N__23492),
            .in1(N__19670),
            .in2(N__19584),
            .in3(N__33346),
            .lcout(),
            .ltout(\c0.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_LC_5_27_5 .C_ON=1'b0;
    defparam \c0.i7_3_lut_LC_5_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_LC_5_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i7_3_lut_LC_5_27_5  (
            .in0(_gnd_net_),
            .in1(N__24280),
            .in2(N__17401),
            .in3(N__23575),
            .lcout(),
            .ltout(\c0.n16_adj_1893_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_920_LC_5_27_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_920_LC_5_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_920_LC_5_27_6 .LUT_INIT=16'b1101111001111011;
    LogicCell40 \c0.i6_4_lut_adj_920_LC_5_27_6  (
            .in0(N__17653),
            .in1(N__19891),
            .in2(N__17638),
            .in3(N__23161),
            .lcout(\c0.n22_adj_1930 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_830_LC_5_27_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_830_LC_5_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_830_LC_5_27_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_830_LC_5_27_7  (
            .in0(_gnd_net_),
            .in1(N__29608),
            .in2(_gnd_net_),
            .in3(N__28025),
            .lcout(\c0.n2058 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_5_28_0 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_5_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_LC_5_28_0  (
            .in0(N__21735),
            .in1(N__17561),
            .in2(N__22623),
            .in3(N__26901),
            .lcout(\c0.n39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_858_LC_5_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_858_LC_5_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_858_LC_5_28_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_858_LC_5_28_1  (
            .in0(_gnd_net_),
            .in1(N__27296),
            .in2(_gnd_net_),
            .in3(N__23546),
            .lcout(),
            .ltout(\c0.n5096_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_861_LC_5_28_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_861_LC_5_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_861_LC_5_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_861_LC_5_28_2  (
            .in0(N__19825),
            .in1(N__20284),
            .in2(N__17614),
            .in3(N__22023),
            .lcout(\c0.n1785 ),
            .ltout(\c0.n1785_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_862_LC_5_28_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_862_LC_5_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_862_LC_5_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_862_LC_5_28_3  (
            .in0(N__30673),
            .in1(N__28304),
            .in2(N__17611),
            .in3(N__25052),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i110_LC_5_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i110_LC_5_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i110_LC_5_28_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i110_LC_5_28_4  (
            .in0(N__36937),
            .in1(N__35996),
            .in2(N__17599),
            .in3(N__17562),
            .lcout(\c0.data_in_field_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_981_LC_5_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_981_LC_5_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_981_LC_5_28_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_981_LC_5_28_5  (
            .in0(N__17560),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19826),
            .lcout(\c0.n5150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_962_LC_5_28_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_962_LC_5_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_962_LC_5_28_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_962_LC_5_28_6  (
            .in0(N__19824),
            .in1(N__17559),
            .in2(_gnd_net_),
            .in3(N__25004),
            .lcout(\c0.n2033 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_896_LC_5_28_7 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_896_LC_5_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_896_LC_5_28_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_896_LC_5_28_7  (
            .in0(N__29739),
            .in1(N__24328),
            .in2(N__33476),
            .in3(N__17764),
            .lcout(\c0.n12_adj_1911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_LC_5_29_0 .C_ON=1'b0;
    defparam \c0.i23_4_lut_LC_5_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_LC_5_29_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_4_lut_LC_5_29_0  (
            .in0(N__17815),
            .in1(N__17809),
            .in2(N__17803),
            .in3(N__17740),
            .lcout(),
            .ltout(\c0.n5275_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_919_LC_5_29_1 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_919_LC_5_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_919_LC_5_29_1 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i8_4_lut_adj_919_LC_5_29_1  (
            .in0(N__17701),
            .in1(N__17791),
            .in2(N__17779),
            .in3(N__20227),
            .lcout(\c0.n24_adj_1929 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_998_LC_5_29_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_998_LC_5_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_998_LC_5_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_998_LC_5_29_2  (
            .in0(N__27657),
            .in1(N__27297),
            .in2(N__17733),
            .in3(N__19641),
            .lcout(\c0.n5182 ),
            .ltout(\c0.n5182_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_LC_5_29_3 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_5_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_LC_5_29_3  (
            .in0(N__17758),
            .in1(N__31554),
            .in2(N__17743),
            .in3(N__23571),
            .lcout(\c0.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_872_LC_5_29_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_872_LC_5_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_872_LC_5_29_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_872_LC_5_29_4  (
            .in0(N__23928),
            .in1(N__30757),
            .in2(N__17734),
            .in3(N__26730),
            .lcout(\c0.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_LC_5_29_5 .C_ON=1'b0;
    defparam \c0.i6_3_lut_LC_5_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_LC_5_29_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i6_3_lut_LC_5_29_5  (
            .in0(N__26260),
            .in1(N__26111),
            .in2(_gnd_net_),
            .in3(N__19870),
            .lcout(\c0.n20_adj_1906 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i36_LC_5_30_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i36_LC_5_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i36_LC_5_30_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i36_LC_5_30_0  (
            .in0(N__35649),
            .in1(N__37132),
            .in2(N__19983),
            .in3(N__17685),
            .lcout(\c0.data_in_field_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35354),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i11_LC_5_30_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i11_LC_5_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i11_LC_5_30_1 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i11_LC_5_30_1  (
            .in0(N__27466),
            .in1(N__35650),
            .in2(N__37229),
            .in3(N__22822),
            .lcout(\c0.data_in_field_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35354),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i135_LC_5_30_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i135_LC_5_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i135_LC_5_30_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i135_LC_5_30_3  (
            .in0(N__24183),
            .in1(N__34220),
            .in2(_gnd_net_),
            .in3(N__17921),
            .lcout(data_in_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35354),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5380_LC_5_30_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5380_LC_5_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5380_LC_5_30_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5380_LC_5_30_4  (
            .in0(N__33286),
            .in1(N__22571),
            .in2(N__32630),
            .in3(N__24085),
            .lcout(\c0.n5731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i134_LC_5_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i134_LC_5_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i134_LC_5_30_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i134_LC_5_30_5  (
            .in0(N__20041),
            .in1(N__24475),
            .in2(N__37230),
            .in3(N__35651),
            .lcout(\c0.data_in_field_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35354),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_989_LC_5_30_6 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_989_LC_5_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_989_LC_5_30_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_989_LC_5_30_6  (
            .in0(N__20005),
            .in1(N__21711),
            .in2(N__28788),
            .in3(N__20040),
            .lcout(\c0.n5264 ),
            .ltout(\c0.n5264_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_990_LC_5_30_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_990_LC_5_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_990_LC_5_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_990_LC_5_30_7  (
            .in0(_gnd_net_),
            .in1(N__20186),
            .in2(N__17881),
            .in3(N__22821),
            .lcout(\c0.n14_adj_1967 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i154_LC_5_31_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i154_LC_5_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i154_LC_5_31_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i154_LC_5_31_0  (
            .in0(N__33884),
            .in1(N__17998),
            .in2(_gnd_net_),
            .in3(N__17866),
            .lcout(data_in_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i26_LC_5_31_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i26_LC_5_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i26_LC_5_31_1 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i26_LC_5_31_1  (
            .in0(N__23788),
            .in1(N__35645),
            .in2(N__37231),
            .in3(N__20188),
            .lcout(\c0.data_in_field_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i146_LC_5_31_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i146_LC_5_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i146_LC_5_31_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i146_LC_5_31_2  (
            .in0(N__33883),
            .in1(N__20085),
            .in2(_gnd_net_),
            .in3(N__17867),
            .lcout(data_in_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i12_LC_5_31_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i12_LC_5_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i12_LC_5_31_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i12_LC_5_31_3  (
            .in0(N__33878),
            .in1(N__17844),
            .in2(_gnd_net_),
            .in3(N__22363),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i8_LC_5_31_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i8_LC_5_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i8_LC_5_31_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i8_LC_5_31_4  (
            .in0(N__35644),
            .in1(N__17982),
            .in2(N__20115),
            .in3(N__37142),
            .lcout(\c0.data_in_field_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i126_LC_5_31_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i126_LC_5_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i126_LC_5_31_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i126_LC_5_31_5  (
            .in0(N__33877),
            .in1(N__24474),
            .in2(_gnd_net_),
            .in3(N__20207),
            .lcout(data_in_15_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_948_LC_5_31_6 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_948_LC_5_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_948_LC_5_31_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i12_4_lut_adj_948_LC_5_31_6  (
            .in0(N__23111),
            .in1(N__24139),
            .in2(N__27585),
            .in3(N__17981),
            .lcout(\c0.n28_adj_1954 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i7_LC_5_31_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i7_LC_5_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i7_LC_5_31_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i7_LC_5_31_7  (
            .in0(N__33879),
            .in1(N__23891),
            .in2(_gnd_net_),
            .in3(N__23112),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_798_LC_5_32_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_798_LC_5_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_798_LC_5_32_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.i1_2_lut_adj_798_LC_5_32_0  (
            .in0(_gnd_net_),
            .in1(N__18357),
            .in2(_gnd_net_),
            .in3(N__18277),
            .lcout(\c0.rx.n5058 ),
            .ltout(\c0.rx.n5058_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_4_lut_4_lut_LC_5_32_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_4_lut_4_lut_LC_5_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_4_lut_4_lut_LC_5_32_1 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \c0.rx.i1_2_lut_4_lut_4_lut_LC_5_32_1  (
            .in0(N__18178),
            .in1(N__18132),
            .in2(N__18070),
            .in3(N__18067),
            .lcout(n1714),
            .ltout(n1714_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_5_32_2 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_5_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_5_32_2 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_5_32_2  (
            .in0(N__17994),
            .in1(N__18016),
            .in2(N__18001),
            .in3(N__20931),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i8_LC_5_32_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i8_LC_5_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i8_LC_5_32_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i8_LC_5_32_3  (
            .in0(N__33876),
            .in1(N__17983),
            .in2(_gnd_net_),
            .in3(N__27578),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_5_32_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_5_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_5_32_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_5_32_4  (
            .in0(N__17968),
            .in1(N__17952),
            .in2(N__22416),
            .in3(N__20932),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i145_LC_5_32_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i145_LC_5_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i145_LC_5_32_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i145_LC_5_32_5  (
            .in0(N__33875),
            .in1(N__33454),
            .in2(_gnd_net_),
            .in3(N__21463),
            .lcout(data_in_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i0_LC_6_17_0 .C_ON=1'b1;
    defparam \c0.data_527__i0_LC_6_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i0_LC_6_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i0_LC_6_17_0  (
            .in0(_gnd_net_),
            .in1(N__18486),
            .in2(_gnd_net_),
            .in3(N__18475),
            .lcout(data_0),
            .ltout(),
            .carryin(bfn_6_17_0_),
            .carryout(\c0.n4385 ),
            .clk(N__35282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i1_LC_6_17_1 .C_ON=1'b1;
    defparam \c0.data_527__i1_LC_6_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i1_LC_6_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i1_LC_6_17_1  (
            .in0(_gnd_net_),
            .in1(N__18462),
            .in2(_gnd_net_),
            .in3(N__18451),
            .lcout(data_1),
            .ltout(),
            .carryin(\c0.n4385 ),
            .carryout(\c0.n4386 ),
            .clk(N__35282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i2_LC_6_17_2 .C_ON=1'b1;
    defparam \c0.data_527__i2_LC_6_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i2_LC_6_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i2_LC_6_17_2  (
            .in0(_gnd_net_),
            .in1(N__18441),
            .in2(_gnd_net_),
            .in3(N__18430),
            .lcout(data_2),
            .ltout(),
            .carryin(\c0.n4386 ),
            .carryout(\c0.n4387 ),
            .clk(N__35282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i3_LC_6_17_3 .C_ON=1'b1;
    defparam \c0.data_527__i3_LC_6_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i3_LC_6_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i3_LC_6_17_3  (
            .in0(_gnd_net_),
            .in1(N__18423),
            .in2(_gnd_net_),
            .in3(N__18412),
            .lcout(data_3),
            .ltout(),
            .carryin(\c0.n4387 ),
            .carryout(\c0.n4388 ),
            .clk(N__35282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i4_LC_6_17_4 .C_ON=1'b1;
    defparam \c0.data_527__i4_LC_6_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i4_LC_6_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i4_LC_6_17_4  (
            .in0(_gnd_net_),
            .in1(N__18843),
            .in2(_gnd_net_),
            .in3(N__18409),
            .lcout(data_4),
            .ltout(),
            .carryin(\c0.n4388 ),
            .carryout(\c0.n4389 ),
            .clk(N__35282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i5_LC_6_17_5 .C_ON=1'b1;
    defparam \c0.data_527__i5_LC_6_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i5_LC_6_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i5_LC_6_17_5  (
            .in0(_gnd_net_),
            .in1(N__18396),
            .in2(_gnd_net_),
            .in3(N__18385),
            .lcout(data_5),
            .ltout(),
            .carryin(\c0.n4389 ),
            .carryout(\c0.n4390 ),
            .clk(N__35282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i6_LC_6_17_6 .C_ON=1'b1;
    defparam \c0.data_527__i6_LC_6_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i6_LC_6_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i6_LC_6_17_6  (
            .in0(_gnd_net_),
            .in1(N__18378),
            .in2(_gnd_net_),
            .in3(N__18367),
            .lcout(data_6),
            .ltout(),
            .carryin(\c0.n4390 ),
            .carryout(\c0.n4391 ),
            .clk(N__35282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i7_LC_6_17_7 .C_ON=1'b1;
    defparam \c0.data_527__i7_LC_6_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i7_LC_6_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i7_LC_6_17_7  (
            .in0(_gnd_net_),
            .in1(N__18618),
            .in2(_gnd_net_),
            .in3(N__18607),
            .lcout(data_7),
            .ltout(),
            .carryin(\c0.n4391 ),
            .carryout(\c0.n4392 ),
            .clk(N__35282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i8_LC_6_18_0 .C_ON=1'b1;
    defparam \c0.data_527__i8_LC_6_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i8_LC_6_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i8_LC_6_18_0  (
            .in0(_gnd_net_),
            .in1(N__18696),
            .in2(_gnd_net_),
            .in3(N__18604),
            .lcout(data_8),
            .ltout(),
            .carryin(bfn_6_18_0_),
            .carryout(\c0.n4393 ),
            .clk(N__35294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i9_LC_6_18_1 .C_ON=1'b1;
    defparam \c0.data_527__i9_LC_6_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i9_LC_6_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i9_LC_6_18_1  (
            .in0(_gnd_net_),
            .in1(N__18591),
            .in2(_gnd_net_),
            .in3(N__18580),
            .lcout(data_9),
            .ltout(),
            .carryin(\c0.n4393 ),
            .carryout(\c0.n4394 ),
            .clk(N__35294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i10_LC_6_18_2 .C_ON=1'b1;
    defparam \c0.data_527__i10_LC_6_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i10_LC_6_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i10_LC_6_18_2  (
            .in0(_gnd_net_),
            .in1(N__19098),
            .in2(_gnd_net_),
            .in3(N__18577),
            .lcout(data_10),
            .ltout(),
            .carryin(\c0.n4394 ),
            .carryout(\c0.n4395 ),
            .clk(N__35294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i11_LC_6_18_3 .C_ON=1'b1;
    defparam \c0.data_527__i11_LC_6_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i11_LC_6_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i11_LC_6_18_3  (
            .in0(_gnd_net_),
            .in1(N__18567),
            .in2(_gnd_net_),
            .in3(N__18556),
            .lcout(data_11),
            .ltout(),
            .carryin(\c0.n4395 ),
            .carryout(\c0.n4396 ),
            .clk(N__35294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i12_LC_6_18_4 .C_ON=1'b1;
    defparam \c0.data_527__i12_LC_6_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i12_LC_6_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i12_LC_6_18_4  (
            .in0(_gnd_net_),
            .in1(N__18549),
            .in2(_gnd_net_),
            .in3(N__18538),
            .lcout(data_12),
            .ltout(),
            .carryin(\c0.n4396 ),
            .carryout(\c0.n4397 ),
            .clk(N__35294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i13_LC_6_18_5 .C_ON=1'b1;
    defparam \c0.data_527__i13_LC_6_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i13_LC_6_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i13_LC_6_18_5  (
            .in0(_gnd_net_),
            .in1(N__18528),
            .in2(_gnd_net_),
            .in3(N__18517),
            .lcout(data_13),
            .ltout(),
            .carryin(\c0.n4397 ),
            .carryout(\c0.n4398 ),
            .clk(N__35294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i14_LC_6_18_6 .C_ON=1'b1;
    defparam \c0.data_527__i14_LC_6_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i14_LC_6_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i14_LC_6_18_6  (
            .in0(_gnd_net_),
            .in1(N__18828),
            .in2(_gnd_net_),
            .in3(N__18514),
            .lcout(data_14),
            .ltout(),
            .carryin(\c0.n4398 ),
            .carryout(\c0.n4399 ),
            .clk(N__35294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i15_LC_6_18_7 .C_ON=1'b0;
    defparam \c0.data_527__i15_LC_6_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i15_LC_6_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i15_LC_6_18_7  (
            .in0(_gnd_net_),
            .in1(N__18504),
            .in2(_gnd_net_),
            .in3(N__18511),
            .lcout(data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i13_LC_6_19_0 .C_ON=1'b0;
    defparam \c0.data_out_0___i13_LC_6_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i13_LC_6_19_0 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i13_LC_6_19_0  (
            .in0(N__18780),
            .in1(N__19209),
            .in2(N__18850),
            .in3(N__19080),
            .lcout(data_out_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i7_LC_6_19_1 .C_ON=1'b0;
    defparam \c0.data_out_0___i7_LC_6_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i7_LC_6_19_1 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0___i7_LC_6_19_1  (
            .in0(N__19082),
            .in1(N__20459),
            .in2(N__18832),
            .in3(N__19213),
            .lcout(data_out_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_6_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_6_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_6_19_2  (
            .in0(N__18779),
            .in1(N__18750),
            .in2(_gnd_net_),
            .in3(N__20415),
            .lcout(),
            .ltout(\c0.n9_adj_1887_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i15_3_lut_3_lut_4_lut_LC_6_19_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i15_3_lut_3_lut_4_lut_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i15_3_lut_3_lut_4_lut_LC_6_19_3 .LUT_INIT=16'b1010100001110111;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i15_3_lut_3_lut_4_lut_LC_6_19_3  (
            .in0(N__21414),
            .in1(N__21321),
            .in2(N__18709),
            .in3(N__20584),
            .lcout(\c0.n15_adj_1889 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i1_LC_6_19_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i1_LC_6_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i1_LC_6_19_4 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.data_out_0___i1_LC_6_19_4  (
            .in0(N__19282),
            .in1(N__18697),
            .in2(N__19223),
            .in3(N__19081),
            .lcout(data_out_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i980_2_lut_LC_6_20_0 .C_ON=1'b0;
    defparam \c0.i980_2_lut_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i980_2_lut_LC_6_20_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i980_2_lut_LC_6_20_0  (
            .in0(_gnd_net_),
            .in1(N__21413),
            .in2(_gnd_net_),
            .in3(N__21320),
            .lcout(\c0.n1236 ),
            .ltout(\c0.n1236_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5231_3_lut_LC_6_20_1 .C_ON=1'b0;
    defparam \c0.i5231_3_lut_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5231_3_lut_LC_6_20_1 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \c0.i5231_3_lut_LC_6_20_1  (
            .in0(N__18685),
            .in1(_gnd_net_),
            .in2(N__18673),
            .in3(N__20585),
            .lcout(),
            .ltout(\c0.n5511_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_6_20_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_6_20_2 .LUT_INIT=16'b1111000010111011;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_6_20_2  (
            .in0(N__18670),
            .in1(N__18664),
            .in2(N__18646),
            .in3(N__21196),
            .lcout(),
            .ltout(tx_data_7_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_6_20_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_6_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_6_20_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_6_20_3  (
            .in0(N__19372),
            .in1(_gnd_net_),
            .in2(N__18643),
            .in3(N__18640),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35304),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_6_20_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_6_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_6_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_6_20_7  (
            .in0(N__19371),
            .in1(N__21130),
            .in2(_gnd_net_),
            .in3(N__19312),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35304),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_833_LC_6_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_833_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_833_LC_6_21_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_833_LC_6_21_4  (
            .in0(N__19292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18954),
            .lcout(n1748),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i3_LC_6_21_6 .C_ON=1'b0;
    defparam \c0.data_out_0___i3_LC_6_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i3_LC_6_21_6 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i3_LC_6_21_6  (
            .in0(N__18955),
            .in1(N__19225),
            .in2(N__19105),
            .in3(N__19087),
            .lcout(data_out_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5827_bdd_4_lut_LC_6_23_7 .C_ON=1'b0;
    defparam \c0.n5827_bdd_4_lut_LC_6_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.n5827_bdd_4_lut_LC_6_23_7 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n5827_bdd_4_lut_LC_6_23_7  (
            .in0(N__34820),
            .in1(N__18928),
            .in2(N__24595),
            .in3(N__20941),
            .lcout(\c0.n5830 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5558_LC_6_24_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5558_LC_6_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5558_LC_6_24_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5558_LC_6_24_0  (
            .in0(N__18870),
            .in1(N__32483),
            .in2(N__18862),
            .in3(N__33186),
            .lcout(\c0.n5941 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i155_LC_6_24_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i155_LC_6_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i155_LC_6_24_1 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i155_LC_6_24_1  (
            .in0(N__35857),
            .in1(N__18888),
            .in2(N__24442),
            .in3(N__36607),
            .lcout(\c0.data_in_frame_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i150_LC_6_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i150_LC_6_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i150_LC_6_24_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i150_LC_6_24_2  (
            .in0(N__36605),
            .in1(N__21523),
            .in2(N__18874),
            .in3(N__35861),
            .lcout(\c0.data_in_frame_18_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i158_LC_6_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i158_LC_6_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i158_LC_6_24_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i158_LC_6_24_3  (
            .in0(N__35858),
            .in1(N__18861),
            .in2(N__24529),
            .in3(N__36608),
            .lcout(\c0.data_in_frame_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i118_LC_6_24_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i118_LC_6_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i118_LC_6_24_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i118_LC_6_24_4  (
            .in0(N__36604),
            .in1(N__35859),
            .in2(N__19447),
            .in3(N__23047),
            .lcout(\c0.data_in_field_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_6_24_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_6_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_6_24_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_LC_6_24_5  (
            .in0(N__19793),
            .in1(N__21517),
            .in2(N__23054),
            .in3(N__23256),
            .lcout(\c0.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i55_LC_6_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i55_LC_6_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i55_LC_6_24_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i55_LC_6_24_6  (
            .in0(N__36606),
            .in1(N__35860),
            .in2(N__26218),
            .in3(N__22864),
            .lcout(\c0.data_in_field_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5445_LC_6_24_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5445_LC_6_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5445_LC_6_24_7 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5445_LC_6_24_7  (
            .in0(N__33185),
            .in1(N__22160),
            .in2(N__32572),
            .in3(N__20272),
            .lcout(\c0.n5809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i98_LC_6_25_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i98_LC_6_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i98_LC_6_25_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i98_LC_6_25_0  (
            .in0(N__34286),
            .in1(N__30975),
            .in2(_gnd_net_),
            .in3(N__25331),
            .lcout(data_in_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_927_LC_6_25_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_927_LC_6_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_927_LC_6_25_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_927_LC_6_25_1  (
            .in0(N__28305),
            .in1(N__19567),
            .in2(N__34636),
            .in3(N__21637),
            .lcout(\c0.n5241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_field_143__I_0_1808_2_lut_LC_6_25_2 .C_ON=1'b0;
    defparam \c0.data_in_field_143__I_0_1808_2_lut_LC_6_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_field_143__I_0_1808_2_lut_LC_6_25_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_in_field_143__I_0_1808_2_lut_LC_6_25_2  (
            .in0(_gnd_net_),
            .in1(N__27137),
            .in2(_gnd_net_),
            .in3(N__25678),
            .lcout(\c0.tx2_transmit_N_1031 ),
            .ltout(\c0.tx2_transmit_N_1031_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_LC_6_25_3 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_6_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_6_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_LC_6_25_3  (
            .in0(N__21496),
            .in1(N__21826),
            .in2(N__19390),
            .in3(N__21901),
            .lcout(\c0.n38_adj_1934 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i13_LC_6_25_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i13_LC_6_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i13_LC_6_25_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i13_LC_6_25_4  (
            .in0(N__34285),
            .in1(N__26155),
            .in2(_gnd_net_),
            .in3(N__22265),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_979_LC_6_25_5 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_979_LC_6_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_4_lut_adj_979_LC_6_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_2_lut_3_lut_4_lut_adj_979_LC_6_25_5  (
            .in0(N__29140),
            .in1(N__24675),
            .in2(N__29218),
            .in3(N__27426),
            .lcout(\c0.n14_adj_1900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i150_LC_6_25_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i150_LC_6_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i150_LC_6_25_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i150_LC_6_25_7  (
            .in0(N__24528),
            .in1(N__34287),
            .in2(_gnd_net_),
            .in3(N__21521),
            .lcout(data_in_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i113_LC_6_26_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i113_LC_6_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i113_LC_6_26_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i113_LC_6_26_0  (
            .in0(N__34460),
            .in1(N__19630),
            .in2(_gnd_net_),
            .in3(N__24351),
            .lcout(data_in_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35333),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_855_LC_6_26_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_855_LC_6_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_855_LC_6_26_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_855_LC_6_26_1  (
            .in0(_gnd_net_),
            .in1(N__20013),
            .in2(_gnd_net_),
            .in3(N__29139),
            .lcout(\c0.n5210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_883_LC_6_26_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_883_LC_6_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_883_LC_6_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_883_LC_6_26_4  (
            .in0(N__30664),
            .in1(N__19591),
            .in2(N__37338),
            .in3(N__19585),
            .lcout(\c0.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_914_LC_6_26_5 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_914_LC_6_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_914_LC_6_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_914_LC_6_26_5  (
            .in0(N__26416),
            .in1(N__30481),
            .in2(N__31030),
            .in3(N__19453),
            .lcout(),
            .ltout(\c0.n5259_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_922_LC_6_26_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_922_LC_6_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_922_LC_6_26_6 .LUT_INIT=16'b1111011011111001;
    LogicCell40 \c0.i5_4_lut_adj_922_LC_6_26_6  (
            .in0(N__23449),
            .in1(N__19561),
            .in2(N__19552),
            .in3(N__21781),
            .lcout(\c0.n21_adj_1933 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_895_LC_6_27_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_895_LC_6_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_895_LC_6_27_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_895_LC_6_27_0  (
            .in0(N__19540),
            .in1(N__21811),
            .in2(N__19531),
            .in3(N__19507),
            .lcout(\c0.n18_adj_1910 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_850_LC_6_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_850_LC_6_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_850_LC_6_27_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_850_LC_6_27_1  (
            .in0(N__22975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21918),
            .lcout(\c0.n5198 ),
            .ltout(\c0.n5198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_6_27_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_6_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_6_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_LC_6_27_2  (
            .in0(N__19486),
            .in1(N__23211),
            .in2(N__19477),
            .in3(N__19474),
            .lcout(\c0.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_888_LC_6_27_3 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_888_LC_6_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_888_LC_6_27_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_888_LC_6_27_3  (
            .in0(N__21810),
            .in1(N__21598),
            .in2(N__24279),
            .in3(N__26629),
            .lcout(\c0.n31_adj_1904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_897_LC_6_27_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_897_LC_6_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_897_LC_6_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_897_LC_6_27_4  (
            .in0(N__19762),
            .in1(N__19885),
            .in2(N__19756),
            .in3(N__27391),
            .lcout(),
            .ltout(\c0.n17_adj_1912_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_905_LC_6_27_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_905_LC_6_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_905_LC_6_27_5 .LUT_INIT=16'b1101011111101011;
    LogicCell40 \c0.i3_4_lut_adj_905_LC_6_27_5  (
            .in0(N__27064),
            .in1(N__19732),
            .in2(N__19726),
            .in3(N__19723),
            .lcout(\c0.n19_adj_1920 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_3_lut_4_lut_LC_6_28_0 .C_ON=1'b0;
    defparam \c0.i14_3_lut_4_lut_LC_6_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_3_lut_4_lut_LC_6_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_3_lut_4_lut_LC_6_28_0  (
            .in0(N__19905),
            .in1(N__22033),
            .in2(N__24960),
            .in3(N__19711),
            .lcout(\c0.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_889_LC_6_28_1 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_889_LC_6_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_889_LC_6_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_889_LC_6_28_1  (
            .in0(N__30404),
            .in1(N__25315),
            .in2(N__23437),
            .in3(N__19642),
            .lcout(),
            .ltout(\c0.n29_adj_1905_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_929_LC_6_28_2 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_929_LC_6_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_929_LC_6_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_929_LC_6_28_2  (
            .in0(N__19861),
            .in1(N__19705),
            .in2(N__19699),
            .in3(N__19696),
            .lcout(\c0.n5278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_LC_6_28_3 .C_ON=1'b0;
    defparam \c0.i4_3_lut_LC_6_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_LC_6_28_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_3_lut_LC_6_28_3  (
            .in0(N__19668),
            .in1(N__33339),
            .in2(_gnd_net_),
            .in3(N__26295),
            .lcout(),
            .ltout(\c0.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_6_28_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_6_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_6_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_6_28_4  (
            .in0(N__22778),
            .in1(N__29885),
            .in2(N__19645),
            .in3(N__23080),
            .lcout(\c0.n1880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_876_LC_6_28_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_876_LC_6_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_876_LC_6_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_876_LC_6_28_6  (
            .in0(N__22437),
            .in1(N__20163),
            .in2(N__19909),
            .in3(N__22102),
            .lcout(\c0.n20_adj_1892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_983_LC_6_29_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_983_LC_6_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_983_LC_6_29_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_983_LC_6_29_0  (
            .in0(N__30865),
            .in1(N__19884),
            .in2(N__28924),
            .in3(N__25957),
            .lcout(),
            .ltout(\c0.n10_adj_1963_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_960_LC_6_29_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_960_LC_6_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_960_LC_6_29_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_960_LC_6_29_1  (
            .in0(N__25676),
            .in1(N__29031),
            .in2(N__19873),
            .in3(N__26004),
            .lcout(\c0.n5114 ),
            .ltout(\c0.n5114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_887_LC_6_29_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_887_LC_6_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_887_LC_6_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_887_LC_6_29_2  (
            .in0(N__28351),
            .in1(N__21894),
            .in2(N__19864),
            .in3(N__25396),
            .lcout(\c0.n30_adj_1903 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i91_LC_6_29_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i91_LC_6_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i91_LC_6_29_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i91_LC_6_29_3  (
            .in0(N__36038),
            .in1(N__37089),
            .in2(N__27310),
            .in3(N__31672),
            .lcout(\c0.data_in_field_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35355),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5390_LC_6_29_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5390_LC_6_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5390_LC_6_29_4 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5390_LC_6_29_4  (
            .in0(N__26005),
            .in1(N__33289),
            .in2(N__32789),
            .in3(N__19791),
            .lcout(\c0.n5743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i88_LC_6_29_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i88_LC_6_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i88_LC_6_29_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i88_LC_6_29_5  (
            .in0(N__36037),
            .in1(N__37088),
            .in2(N__22705),
            .in3(N__19830),
            .lcout(\c0.data_in_field_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35355),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i58_LC_6_29_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i58_LC_6_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i58_LC_6_29_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i58_LC_6_29_6  (
            .in0(N__37087),
            .in1(N__36039),
            .in2(N__23986),
            .in3(N__19792),
            .lcout(\c0.data_in_field_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35355),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1000_LC_6_30_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1000_LC_6_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1000_LC_6_30_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1000_LC_6_30_0  (
            .in0(N__21976),
            .in1(N__19969),
            .in2(N__32950),
            .in3(N__22995),
            .lcout(\c0.n5162 ),
            .ltout(\c0.n5162_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_819_LC_6_30_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_819_LC_6_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_819_LC_6_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_819_LC_6_30_1  (
            .in0(_gnd_net_),
            .in1(N__20105),
            .in2(N__20089),
            .in3(N__25250),
            .lcout(\c0.n1825 ),
            .ltout(\c0.n1825_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_869_LC_6_30_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_869_LC_6_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_869_LC_6_30_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_869_LC_6_30_2  (
            .in0(N__20071),
            .in1(N__26380),
            .in2(N__20053),
            .in3(N__20043),
            .lcout(\c0.n28_adj_1886 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i95_LC_6_30_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i95_LC_6_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i95_LC_6_30_3 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i95_LC_6_30_3  (
            .in0(N__32938),
            .in1(N__36992),
            .in2(N__31288),
            .in3(N__35653),
            .lcout(\c0.data_in_field_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i96_LC_6_30_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i96_LC_6_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i96_LC_6_30_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i96_LC_6_30_4  (
            .in0(N__36990),
            .in1(N__35643),
            .in2(N__22735),
            .in3(N__22997),
            .lcout(\c0.data_in_field_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i74_LC_6_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i74_LC_6_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i74_LC_6_30_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i74_LC_6_30_5  (
            .in0(N__35641),
            .in1(N__36991),
            .in2(N__26554),
            .in3(N__20012),
            .lcout(\c0.data_in_field_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i23_LC_6_30_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i23_LC_6_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i23_LC_6_30_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i23_LC_6_30_6  (
            .in0(N__27891),
            .in1(N__35642),
            .in2(N__37161),
            .in3(N__22238),
            .lcout(\c0.data_in_field_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35363),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_LC_6_30_7 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_LC_6_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_LC_6_30_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_3_lut_4_lut_LC_6_30_7  (
            .in0(N__22996),
            .in1(N__25084),
            .in2(N__19979),
            .in3(N__31555),
            .lcout(\c0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i80_LC_6_31_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i80_LC_6_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i80_LC_6_31_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i80_LC_6_31_0  (
            .in0(N__23828),
            .in1(_gnd_net_),
            .in2(N__34296),
            .in3(N__22695),
            .lcout(data_in_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i138_LC_6_31_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i138_LC_6_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i138_LC_6_31_1 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i138_LC_6_31_1  (
            .in0(N__20812),
            .in1(N__37285),
            .in2(N__35837),
            .in3(N__19923),
            .lcout(\c0.data_in_field_137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_829_LC_6_31_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_829_LC_6_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_829_LC_6_31_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_829_LC_6_31_2  (
            .in0(N__19922),
            .in1(N__20263),
            .in2(_gnd_net_),
            .in3(N__22303),
            .lcout(\c0.n2043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_860_LC_6_31_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_860_LC_6_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_860_LC_6_31_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_860_LC_6_31_3  (
            .in0(N__20264),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25143),
            .lcout(\c0.n6_adj_1877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i32_LC_6_31_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i32_LC_6_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i32_LC_6_31_4 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i32_LC_6_31_4  (
            .in0(N__35768),
            .in1(N__24052),
            .in2(N__37290),
            .in3(N__20265),
            .lcout(\c0.data_in_field_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_871_LC_6_31_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_871_LC_6_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_871_LC_6_31_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_871_LC_6_31_5  (
            .in0(N__22389),
            .in1(N__20248),
            .in2(N__20242),
            .in3(N__22504),
            .lcout(\c0.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_956_LC_6_31_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_956_LC_6_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_956_LC_6_31_6 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i1_4_lut_adj_956_LC_6_31_6  (
            .in0(N__23275),
            .in1(N__27811),
            .in2(N__22639),
            .in3(N__22321),
            .lcout(\c0.n1686 ),
            .ltout(\c0.n1686_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i126_LC_6_31_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i126_LC_6_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i126_LC_6_31_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i126_LC_6_31_7  (
            .in0(N__20217),
            .in1(N__37281),
            .in2(N__20191),
            .in3(N__28810),
            .lcout(\c0.data_in_field_125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5400_LC_6_32_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5400_LC_6_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5400_LC_6_32_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5400_LC_6_32_0  (
            .in0(N__33309),
            .in1(N__20187),
            .in2(N__32735),
            .in3(N__22307),
            .lcout(\c0.n5749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i24_LC_6_32_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i24_LC_6_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i24_LC_6_32_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i24_LC_6_32_1  (
            .in0(N__34010),
            .in1(N__24048),
            .in2(_gnd_net_),
            .in3(N__22670),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i114_LC_6_32_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i114_LC_6_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i114_LC_6_32_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i114_LC_6_32_2  (
            .in0(N__37201),
            .in1(N__35640),
            .in2(N__31012),
            .in3(N__22567),
            .lcout(\c0.data_in_field_113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i160_LC_6_32_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i160_LC_6_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i160_LC_6_32_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i160_LC_6_32_3  (
            .in0(N__34009),
            .in1(N__20820),
            .in2(_gnd_net_),
            .in3(N__20149),
            .lcout(data_in_19_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_6_32_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_6_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_6_32_4 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_6_32_4  (
            .in0(N__20916),
            .in1(N__20850),
            .in2(N__20824),
            .in3(N__20839),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i130_LC_6_32_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i130_LC_6_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i130_LC_6_32_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i130_LC_6_32_6  (
            .in0(N__20811),
            .in1(N__34011),
            .in2(_gnd_net_),
            .in3(N__30203),
            .lcout(data_in_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i136_LC_6_32_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i136_LC_6_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i136_LC_6_32_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i136_LC_6_32_7  (
            .in0(N__35639),
            .in1(N__37202),
            .in2(N__25618),
            .in3(N__22603),
            .lcout(\c0.data_in_field_135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3325_2_lut_LC_7_17_7 .C_ON=1'b0;
    defparam \c0.i3325_2_lut_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3325_2_lut_LC_7_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i3325_2_lut_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__20530),
            .in2(_gnd_net_),
            .in3(N__20355),
            .lcout(\c0.n3567 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5247_4_lut_4_lut_LC_7_18_3 .C_ON=1'b0;
    defparam \c0.i5247_4_lut_4_lut_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5247_4_lut_4_lut_LC_7_18_3 .LUT_INIT=16'b1101110111110101;
    LogicCell40 \c0.i5247_4_lut_4_lut_LC_7_18_3  (
            .in0(N__20582),
            .in1(N__20785),
            .in2(N__20770),
            .in3(N__20416),
            .lcout(\c0.n5515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_892_LC_7_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_892_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_892_LC_7_18_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_892_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(N__20647),
            .in2(_gnd_net_),
            .in3(N__20749),
            .lcout(n5176),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_972_LC_7_18_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_972_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_972_LC_7_18_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_972_LC_7_18_6  (
            .in0(N__21412),
            .in1(N__21319),
            .in2(_gnd_net_),
            .in3(N__20581),
            .lcout(\c0.n1590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5259_4_lut_4_lut_LC_7_19_3 .C_ON=1'b0;
    defparam \c0.i5259_4_lut_4_lut_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5259_4_lut_4_lut_LC_7_19_3 .LUT_INIT=16'b1011101111110011;
    LogicCell40 \c0.i5259_4_lut_4_lut_LC_7_19_3  (
            .in0(N__20643),
            .in1(N__20583),
            .in2(N__20469),
            .in3(N__20414),
            .lcout(),
            .ltout(\c0.n5523_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5256_4_lut_LC_7_19_4 .C_ON=1'b0;
    defparam \c0.i5256_4_lut_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5256_4_lut_LC_7_19_4 .LUT_INIT=16'b1111111111010001;
    LogicCell40 \c0.i5256_4_lut_LC_7_19_4  (
            .in0(N__21427),
            .in1(N__21418),
            .in2(N__21325),
            .in3(N__21322),
            .lcout(),
            .ltout(\c0.n5513_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_7_19_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_7_19_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_7_19_5  (
            .in0(N__21231),
            .in1(N__21205),
            .in2(N__21199),
            .in3(N__21195),
            .lcout(tx_data_6_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_980_LC_7_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_980_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_980_LC_7_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_980_LC_7_22_6  (
            .in0(N__21124),
            .in1(N__21078),
            .in2(_gnd_net_),
            .in3(N__21016),
            .lcout(n5132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5470_LC_7_23_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5470_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5470_LC_7_23_0 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5470_LC_7_23_0  (
            .in0(N__33275),
            .in1(N__30546),
            .in2(N__32777),
            .in3(N__27016),
            .lcout(),
            .ltout(\c0.n5839_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5839_bdd_4_lut_LC_7_23_1 .C_ON=1'b0;
    defparam \c0.n5839_bdd_4_lut_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5839_bdd_4_lut_LC_7_23_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5839_bdd_4_lut_LC_7_23_1  (
            .in0(N__32775),
            .in1(N__26379),
            .in2(N__20956),
            .in3(N__29686),
            .lcout(\c0.n5414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5465_LC_7_23_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5465_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5465_LC_7_23_2 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5465_LC_7_23_2  (
            .in0(N__33276),
            .in1(N__31114),
            .in2(N__32778),
            .in3(N__25117),
            .lcout(),
            .ltout(\c0.n5833_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5833_bdd_4_lut_LC_7_23_3 .C_ON=1'b0;
    defparam \c0.n5833_bdd_4_lut_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5833_bdd_4_lut_LC_7_23_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5833_bdd_4_lut_LC_7_23_3  (
            .in0(N__32776),
            .in1(N__27187),
            .in2(N__20953),
            .in3(N__28669),
            .lcout(),
            .ltout(\c0.n5417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5480_LC_7_23_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5480_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5480_LC_7_23_4 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5480_LC_7_23_4  (
            .in0(N__34813),
            .in1(N__32122),
            .in2(N__20950),
            .in3(N__20947),
            .lcout(\c0.n5827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5351_LC_7_24_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5351_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5351_LC_7_24_0 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5351_LC_7_24_0  (
            .in0(N__33201),
            .in1(N__29889),
            .in2(N__32582),
            .in3(N__25162),
            .lcout(\c0.n5695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5341_LC_7_24_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5341_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5341_LC_7_24_1 .LUT_INIT=16'b1011100011001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5341_LC_7_24_1  (
            .in0(N__23500),
            .in1(N__33202),
            .in2(N__24327),
            .in3(N__32502),
            .lcout(),
            .ltout(\c0.n5683_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5683_bdd_4_lut_LC_7_24_2 .C_ON=1'b0;
    defparam \c0.n5683_bdd_4_lut_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.n5683_bdd_4_lut_LC_7_24_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5683_bdd_4_lut_LC_7_24_2  (
            .in0(N__32503),
            .in1(N__22950),
            .in2(N__21553),
            .in3(N__23149),
            .lcout(\c0.n5483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5695_bdd_4_lut_LC_7_24_3 .C_ON=1'b0;
    defparam \c0.n5695_bdd_4_lut_LC_7_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5695_bdd_4_lut_LC_7_24_3 .LUT_INIT=16'b1010101011100100;
    LogicCell40 \c0.n5695_bdd_4_lut_LC_7_24_3  (
            .in0(N__21550),
            .in1(N__29032),
            .in2(N__29467),
            .in3(N__32504),
            .lcout(),
            .ltout(\c0.n5480_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5370_LC_7_24_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5370_LC_7_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5370_LC_7_24_4 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5370_LC_7_24_4  (
            .in0(N__34804),
            .in1(N__32123),
            .in2(N__21544),
            .in3(N__21541),
            .lcout(),
            .ltout(\c0.n5677_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5677_bdd_4_lut_LC_7_24_5 .C_ON=1'b0;
    defparam \c0.n5677_bdd_4_lut_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n5677_bdd_4_lut_LC_7_24_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5677_bdd_4_lut_LC_7_24_5  (
            .in0(N__34812),
            .in1(N__24865),
            .in2(N__21535),
            .in3(N__28207),
            .lcout(\c0.n5680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i90_LC_7_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i90_LC_7_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i90_LC_7_24_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i90_LC_7_24_7  (
            .in0(N__34543),
            .in1(N__25332),
            .in2(_gnd_net_),
            .in3(N__28589),
            .lcout(data_in_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35327),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i142_LC_7_25_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i142_LC_7_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i142_LC_7_25_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i142_LC_7_25_0  (
            .in0(N__34367),
            .in1(N__24003),
            .in2(_gnd_net_),
            .in3(N__21522),
            .lcout(data_in_17_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_LC_7_25_1 .C_ON=1'b0;
    defparam \c0.i3_2_lut_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_LC_7_25_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_LC_7_25_1  (
            .in0(_gnd_net_),
            .in1(N__21445),
            .in2(_gnd_net_),
            .in3(N__25056),
            .lcout(\c0.n24_adj_1895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i153_LC_7_25_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i153_LC_7_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i153_LC_7_25_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i153_LC_7_25_2  (
            .in0(N__21446),
            .in1(_gnd_net_),
            .in2(N__34505),
            .in3(N__21490),
            .lcout(data_in_19_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5797_bdd_4_lut_LC_7_25_3 .C_ON=1'b0;
    defparam \c0.n5797_bdd_4_lut_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5797_bdd_4_lut_LC_7_25_3 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n5797_bdd_4_lut_LC_7_25_3  (
            .in0(N__23392),
            .in1(N__24898),
            .in2(N__23260),
            .in3(N__32454),
            .lcout(\c0.n5429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5791_bdd_4_lut_LC_7_25_5 .C_ON=1'b0;
    defparam \c0.n5791_bdd_4_lut_LC_7_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.n5791_bdd_4_lut_LC_7_25_5 .LUT_INIT=16'b1100111011000010;
    LogicCell40 \c0.n5791_bdd_4_lut_LC_7_25_5  (
            .in0(N__21592),
            .in1(N__21763),
            .in2(N__32571),
            .in3(N__30405),
            .lcout(\c0.n5432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5530_LC_7_25_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5530_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5530_LC_7_25_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5530_LC_7_25_6  (
            .in0(N__33285),
            .in1(N__21742),
            .in2(N__32546),
            .in3(N__22246),
            .lcout(\c0.n5911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5881_bdd_4_lut_LC_7_25_7 .C_ON=1'b0;
    defparam \c0.n5881_bdd_4_lut_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.n5881_bdd_4_lut_LC_7_25_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5881_bdd_4_lut_LC_7_25_7  (
            .in0(N__32476),
            .in1(N__21715),
            .in2(N__23707),
            .in3(N__25534),
            .lcout(\c0.n5393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i120_LC_7_26_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i120_LC_7_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i120_LC_7_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i120_LC_7_26_1  (
            .in0(N__34378),
            .in1(N__27688),
            .in2(_gnd_net_),
            .in3(N__21648),
            .lcout(data_in_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_882_LC_7_26_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_882_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_882_LC_7_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_882_LC_7_26_2  (
            .in0(N__27085),
            .in1(N__26112),
            .in2(N__26272),
            .in3(N__26905),
            .lcout(\c0.n10_adj_1898 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i70_LC_7_26_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i70_LC_7_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i70_LC_7_26_3 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i70_LC_7_26_3  (
            .in0(N__21617),
            .in1(N__36691),
            .in2(N__22498),
            .in3(N__36201),
            .lcout(\c0.data_in_field_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_997_LC_7_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_997_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_997_LC_7_26_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_997_LC_7_26_4  (
            .in0(_gnd_net_),
            .in1(N__21616),
            .in2(_gnd_net_),
            .in3(N__22865),
            .lcout(\c0.n5159 ),
            .ltout(\c0.n5159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1001_LC_7_26_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1001_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1001_LC_7_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1001_LC_7_26_5  (
            .in0(N__26365),
            .in1(N__21588),
            .in2(N__21556),
            .in3(N__22785),
            .lcout(\c0.n1978 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_827_LC_7_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_827_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_827_LC_7_26_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_827_LC_7_26_6  (
            .in0(_gnd_net_),
            .in1(N__21955),
            .in2(_gnd_net_),
            .in3(N__23491),
            .lcout(),
            .ltout(\c0.n2095_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_880_LC_7_26_7 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_880_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_880_LC_7_26_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_880_LC_7_26_7  (
            .in0(N__22089),
            .in1(N__22897),
            .in2(N__21925),
            .in3(N__21922),
            .lcout(\c0.n34_adj_1896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5460_LC_7_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5460_LC_7_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5460_LC_7_27_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5460_LC_7_27_0  (
            .in0(N__33290),
            .in1(N__21837),
            .in2(N__32790),
            .in3(N__23380),
            .lcout(),
            .ltout(\c0.n5821_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5821_bdd_4_lut_LC_7_27_1 .C_ON=1'b0;
    defparam \c0.n5821_bdd_4_lut_LC_7_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5821_bdd_4_lut_LC_7_27_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5821_bdd_4_lut_LC_7_27_1  (
            .in0(N__32755),
            .in1(N__21895),
            .in2(N__21856),
            .in3(N__31714),
            .lcout(\c0.n5423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i28_LC_7_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i28_LC_7_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i28_LC_7_27_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i28_LC_7_27_2  (
            .in0(N__36227),
            .in1(N__21838),
            .in2(N__23323),
            .in3(N__36785),
            .lcout(\c0.data_in_field_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i13_LC_7_27_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i13_LC_7_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i13_LC_7_27_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i13_LC_7_27_3  (
            .in0(N__24617),
            .in1(N__22272),
            .in2(N__36999),
            .in3(N__36228),
            .lcout(\c0.data_in_field_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_977_LC_7_27_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_977_LC_7_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_977_LC_7_27_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_977_LC_7_27_4  (
            .in0(_gnd_net_),
            .in1(N__21836),
            .in2(_gnd_net_),
            .in3(N__24616),
            .lcout(\c0.n2080 ),
            .ltout(\c0.n2080_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_978_LC_7_27_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_978_LC_7_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_978_LC_7_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_978_LC_7_27_5  (
            .in0(N__26375),
            .in1(N__26325),
            .in2(N__21814),
            .in3(N__32830),
            .lcout(\c0.n5243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_915_LC_7_27_6 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_915_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_915_LC_7_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_915_LC_7_27_6  (
            .in0(N__30826),
            .in1(N__28326),
            .in2(N__21802),
            .in3(N__22077),
            .lcout(\c0.n25_adj_1926 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_969_LC_7_27_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_969_LC_7_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_969_LC_7_27_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_969_LC_7_27_7  (
            .in0(_gnd_net_),
            .in1(N__24340),
            .in2(_gnd_net_),
            .in3(N__22090),
            .lcout(\c0.n5261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5346_LC_7_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5346_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5346_LC_7_28_0 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5346_LC_7_28_0  (
            .in0(N__33294),
            .in1(N__22193),
            .in2(N__26740),
            .in3(N__32785),
            .lcout(),
            .ltout(\c0.n5689_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5689_bdd_4_lut_LC_7_28_1 .C_ON=1'b0;
    defparam \c0.n5689_bdd_4_lut_LC_7_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5689_bdd_4_lut_LC_7_28_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5689_bdd_4_lut_LC_7_28_1  (
            .in0(N__32756),
            .in1(N__27721),
            .in2(N__22063),
            .in3(N__25564),
            .lcout(\c0.n5366 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i56_LC_7_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i56_LC_7_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i56_LC_7_28_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i56_LC_7_28_2  (
            .in0(N__36017),
            .in1(N__36881),
            .in2(N__23812),
            .in3(N__22194),
            .lcout(\c0.data_in_field_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35356),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i133_LC_7_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i133_LC_7_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i133_LC_7_28_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i133_LC_7_28_3  (
            .in0(N__36880),
            .in1(N__36018),
            .in2(N__28195),
            .in3(N__27424),
            .lcout(\c0.data_in_field_132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35356),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_993_LC_7_28_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_993_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_993_LC_7_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_993_LC_7_28_4  (
            .in0(N__22045),
            .in1(N__29422),
            .in2(N__29743),
            .in3(N__22171),
            .lcout(\c0.n5276 ),
            .ltout(\c0.n5276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_924_LC_7_28_5 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_924_LC_7_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_924_LC_7_28_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_adj_924_LC_7_28_5  (
            .in0(N__22027),
            .in1(N__27262),
            .in2(N__22012),
            .in3(N__25938),
            .lcout(\c0.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i37_LC_7_29_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i37_LC_7_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i37_LC_7_29_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i37_LC_7_29_0  (
            .in0(N__36030),
            .in1(N__37070),
            .in2(N__21992),
            .in3(N__30073),
            .lcout(\c0.data_in_field_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35364),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i86_LC_7_29_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i86_LC_7_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i86_LC_7_29_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i86_LC_7_29_1  (
            .in0(N__37069),
            .in1(N__36032),
            .in2(N__27550),
            .in3(N__23600),
            .lcout(\c0.data_in_field_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35364),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_818_LC_7_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_818_LC_7_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_818_LC_7_29_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_818_LC_7_29_2  (
            .in0(N__24661),
            .in1(N__27414),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n2005_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_820_LC_7_29_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_820_LC_7_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_820_LC_7_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_820_LC_7_29_3  (
            .in0(N__22231),
            .in1(N__31048),
            .in2(N__22210),
            .in3(N__23239),
            .lcout(),
            .ltout(\c0.n10_adj_1873_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_821_LC_7_29_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_821_LC_7_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_821_LC_7_29_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i5_3_lut_adj_821_LC_7_29_4  (
            .in0(N__28250),
            .in1(_gnd_net_),
            .in2(N__22207),
            .in3(N__22204),
            .lcout(\c0.n5111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i53_LC_7_29_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i53_LC_7_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i53_LC_7_29_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i53_LC_7_29_5  (
            .in0(N__37068),
            .in1(N__36031),
            .in2(N__30037),
            .in3(N__31049),
            .lcout(\c0.data_in_field_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35364),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_3_lut_LC_7_29_6 .C_ON=1'b0;
    defparam \c0.i4_2_lut_3_lut_LC_7_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_3_lut_LC_7_29_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_2_lut_3_lut_LC_7_29_6  (
            .in0(N__25410),
            .in1(N__22189),
            .in2(_gnd_net_),
            .in3(N__22141),
            .lcout(\c0.n13_adj_1951 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i21_LC_7_29_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i21_LC_7_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i21_LC_7_29_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i21_LC_7_29_7  (
            .in0(N__24668),
            .in1(N__26154),
            .in2(N__37200),
            .in3(N__36033),
            .lcout(\c0.data_in_field_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35364),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i24_LC_7_30_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i24_LC_7_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i24_LC_7_30_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i24_LC_7_30_0  (
            .in0(N__35646),
            .in1(N__22145),
            .in2(N__22678),
            .in3(N__36998),
            .lcout(\c0.data_in_field_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i54_LC_7_30_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i54_LC_7_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i54_LC_7_30_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i54_LC_7_30_1  (
            .in0(N__34167),
            .in1(N__24246),
            .in2(_gnd_net_),
            .in3(N__28100),
            .lcout(data_in_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_875_LC_7_30_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_875_LC_7_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_875_LC_7_30_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_875_LC_7_30_2  (
            .in0(N__23921),
            .in1(N__33403),
            .in2(N__22117),
            .in3(N__33359),
            .lcout(\c0.n18_adj_1891 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_945_LC_7_30_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_945_LC_7_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_945_LC_7_30_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_945_LC_7_30_3  (
            .in0(N__22534),
            .in1(N__26946),
            .in2(_gnd_net_),
            .in3(N__25493),
            .lcout(\c0.n5249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i68_LC_7_30_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i68_LC_7_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i68_LC_7_30_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i68_LC_7_30_4  (
            .in0(N__35647),
            .in1(N__36996),
            .in2(N__33535),
            .in3(N__23248),
            .lcout(\c0.data_in_field_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i155_LC_7_30_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i155_LC_7_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i155_LC_7_30_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i155_LC_7_30_5  (
            .in0(N__34166),
            .in1(N__22423),
            .in2(_gnd_net_),
            .in3(N__24416),
            .lcout(data_in_19_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i89_LC_7_30_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i89_LC_7_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i89_LC_7_30_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i89_LC_7_30_6  (
            .in0(N__35648),
            .in1(N__36997),
            .in2(N__28543),
            .in3(N__25150),
            .lcout(\c0.data_in_field_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35372),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_946_LC_7_30_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_946_LC_7_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_946_LC_7_30_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_946_LC_7_30_7  (
            .in0(N__25668),
            .in1(N__26945),
            .in2(_gnd_net_),
            .in3(N__25492),
            .lcout(\c0.n5255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_951_LC_7_31_0 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_951_LC_7_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_951_LC_7_31_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i9_4_lut_adj_951_LC_7_31_0  (
            .in0(N__22364),
            .in1(N__29239),
            .in2(N__22282),
            .in3(N__31416),
            .lcout(),
            .ltout(\c0.n25_adj_1957_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_954_LC_7_31_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_954_LC_7_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_954_LC_7_31_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i15_4_lut_adj_954_LC_7_31_1  (
            .in0(N__22342),
            .in1(N__22333),
            .in2(N__22324),
            .in3(N__22645),
            .lcout(\c0.n4465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i18_LC_7_31_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i18_LC_7_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i18_LC_7_31_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i18_LC_7_31_2  (
            .in0(N__30187),
            .in1(N__35652),
            .in2(N__37291),
            .in3(N__22308),
            .lcout(\c0.data_in_field_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i5_LC_7_31_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i5_LC_7_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i5_LC_7_31_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i5_LC_7_31_3  (
            .in0(N__34168),
            .in1(N__22281),
            .in2(_gnd_net_),
            .in3(N__26394),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_854_LC_7_31_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_854_LC_7_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_854_LC_7_31_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_854_LC_7_31_4  (
            .in0(N__27012),
            .in1(N__25452),
            .in2(_gnd_net_),
            .in3(N__31786),
            .lcout(\c0.n1772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i88_LC_7_31_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i88_LC_7_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i88_LC_7_31_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i88_LC_7_31_5  (
            .in0(N__22734),
            .in1(_gnd_net_),
            .in2(N__34379),
            .in3(N__22694),
            .lcout(data_in_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_950_LC_7_31_7 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_950_LC_7_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_950_LC_7_31_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i11_4_lut_adj_950_LC_7_31_7  (
            .in0(N__30153),
            .in1(N__26393),
            .in2(N__29656),
            .in3(N__22663),
            .lcout(\c0.n27_adj_1956 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i19_LC_7_32_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i19_LC_7_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i19_LC_7_32_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i19_LC_7_32_0  (
            .in0(N__34012),
            .in1(N__29412),
            .in2(_gnd_net_),
            .in3(N__29246),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35385),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_952_LC_7_32_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_952_LC_7_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_952_LC_7_32_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_952_LC_7_32_1  (
            .in0(N__24047),
            .in1(N__23892),
            .in2(N__25912),
            .in3(N__23773),
            .lcout(\c0.n26_adj_1958 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_856_LC_7_32_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_856_LC_7_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_856_LC_7_32_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_856_LC_7_32_3  (
            .in0(N__27650),
            .in1(N__22597),
            .in2(N__22572),
            .in3(N__22533),
            .lcout(\c0.n5144 ),
            .ltout(\c0.n5144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_LC_7_32_4 .C_ON=1'b0;
    defparam \c0.i13_4_lut_LC_7_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_LC_7_32_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_LC_7_32_4  (
            .in0(N__23215),
            .in1(N__25201),
            .in2(N__22507),
            .in3(N__22954),
            .lcout(\c0.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i70_LC_7_32_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i70_LC_7_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i70_LC_7_32_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i70_LC_7_32_5  (
            .in0(N__34015),
            .in1(N__27517),
            .in2(_gnd_net_),
            .in3(N__22484),
            .lcout(data_in_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35385),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i64_LC_7_32_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i64_LC_7_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i64_LC_7_32_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i64_LC_7_32_6  (
            .in0(N__34013),
            .in1(N__22464),
            .in2(_gnd_net_),
            .in3(N__24101),
            .lcout(data_in_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35385),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i26_LC_7_32_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i26_LC_7_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i26_LC_7_32_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i26_LC_7_32_7  (
            .in0(N__34014),
            .in1(N__29335),
            .in2(_gnd_net_),
            .in3(N__23774),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35385),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5761_bdd_4_lut_LC_9_23_1 .C_ON=1'b0;
    defparam \c0.n5761_bdd_4_lut_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5761_bdd_4_lut_LC_9_23_1 .LUT_INIT=16'b1100101111001000;
    LogicCell40 \c0.n5761_bdd_4_lut_LC_9_23_1  (
            .in0(N__25770),
            .in1(N__22741),
            .in2(N__32698),
            .in3(N__24840),
            .lcout(),
            .ltout(\c0.n5447_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5420_LC_9_23_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5420_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5420_LC_9_23_2 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5420_LC_9_23_2  (
            .in0(N__34828),
            .in1(N__32124),
            .in2(N__22888),
            .in3(N__22747),
            .lcout(),
            .ltout(\c0.n5755_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5755_bdd_4_lut_LC_9_23_3 .C_ON=1'b0;
    defparam \c0.n5755_bdd_4_lut_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5755_bdd_4_lut_LC_9_23_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5755_bdd_4_lut_LC_9_23_3  (
            .in0(N__34829),
            .in1(N__28219),
            .in2(N__22885),
            .in3(N__22795),
            .lcout(\c0.n5758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5525_LC_9_24_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5525_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5525_LC_9_24_0 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5525_LC_9_24_0  (
            .in0(N__33184),
            .in1(N__22869),
            .in2(N__26671),
            .in3(N__32667),
            .lcout(\c0.n5905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5779_bdd_4_lut_LC_9_24_2 .C_ON=1'b0;
    defparam \c0.n5779_bdd_4_lut_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.n5779_bdd_4_lut_LC_9_24_2 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n5779_bdd_4_lut_LC_9_24_2  (
            .in0(N__27226),
            .in1(N__32674),
            .in2(N__24394),
            .in3(N__22834),
            .lcout(\c0.n5438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5410_LC_9_24_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5410_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5410_LC_9_24_3 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5410_LC_9_24_3  (
            .in0(N__33182),
            .in1(N__22789),
            .in2(N__32697),
            .in3(N__27319),
            .lcout(),
            .ltout(\c0.n5767_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5767_bdd_4_lut_LC_9_24_4 .C_ON=1'b0;
    defparam \c0.n5767_bdd_4_lut_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.n5767_bdd_4_lut_LC_9_24_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5767_bdd_4_lut_LC_9_24_4  (
            .in0(N__32505),
            .in1(N__31204),
            .in2(N__22750),
            .in3(N__30580),
            .lcout(\c0.n5444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5405_LC_9_24_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5405_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5405_LC_9_24_5 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5405_LC_9_24_5  (
            .in0(N__33183),
            .in1(N__30668),
            .in2(N__32696),
            .in3(N__31953),
            .lcout(\c0.n5761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i55_LC_9_25_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i55_LC_9_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i55_LC_9_25_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i55_LC_9_25_0  (
            .in0(N__34466),
            .in1(N__26523),
            .in2(_gnd_net_),
            .in3(N__26195),
            .lcout(data_in_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i97_LC_9_25_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i97_LC_9_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i97_LC_9_25_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i97_LC_9_25_1  (
            .in0(N__36953),
            .in1(N__35862),
            .in2(N__23098),
            .in3(N__22925),
            .lcout(\c0.data_in_field_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_9_25_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_9_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_LC_9_25_2  (
            .in0(N__28456),
            .in1(N__23138),
            .in2(N__22936),
            .in3(N__30572),
            .lcout(\c0.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i85_LC_9_25_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i85_LC_9_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i85_LC_9_25_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i85_LC_9_25_3  (
            .in0(N__27054),
            .in1(N__34467),
            .in2(_gnd_net_),
            .in3(N__26489),
            .lcout(data_in_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_957_LC_9_25_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_957_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_957_LC_9_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_957_LC_9_25_4  (
            .in0(N__23539),
            .in1(N__29294),
            .in2(N__27318),
            .in3(N__28257),
            .lcout(\c0.n2074 ),
            .ltout(\c0.n2074_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_996_LC_9_25_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_996_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_996_LC_9_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_996_LC_9_25_5  (
            .in0(N__23067),
            .in1(N__25533),
            .in2(N__23026),
            .in3(N__25292),
            .lcout(\c0.n5213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_970_LC_9_26_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_970_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_970_LC_9_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_970_LC_9_26_0  (
            .in0(N__25251),
            .in1(N__29799),
            .in2(N__22971),
            .in3(N__32964),
            .lcout(\c0.n10_adj_1888 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_848_LC_9_26_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_848_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_848_LC_9_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_848_LC_9_26_1  (
            .in0(N__25560),
            .in1(N__22926),
            .in2(_gnd_net_),
            .in3(N__23008),
            .lcout(\c0.n1851 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_966_LC_9_26_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_966_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_966_LC_9_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_966_LC_9_26_2  (
            .in0(N__22927),
            .in1(N__28457),
            .in2(N__24740),
            .in3(N__24970),
            .lcout(\c0.n5099 ),
            .ltout(\c0.n5099_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_877_LC_9_26_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_877_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_877_LC_9_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_877_LC_9_26_3  (
            .in0(N__23191),
            .in1(N__23175),
            .in2(N__23164),
            .in3(N__30260),
            .lcout(\c0.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i105_LC_9_26_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i105_LC_9_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i105_LC_9_26_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i105_LC_9_26_4  (
            .in0(N__36194),
            .in1(N__37222),
            .in2(N__23148),
            .in3(N__24382),
            .lcout(\c0.data_in_field_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i7_LC_9_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i7_LC_9_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i7_LC_9_26_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i7_LC_9_26_5  (
            .in0(N__28458),
            .in1(N__23122),
            .in2(N__37272),
            .in3(N__36195),
            .lcout(\c0.data_in_field_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i97_LC_9_26_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i97_LC_9_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i97_LC_9_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i97_LC_9_26_6  (
            .in0(N__34464),
            .in1(N__24381),
            .in2(_gnd_net_),
            .in3(N__23093),
            .lcout(data_in_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i89_LC_9_26_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i89_LC_9_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i89_LC_9_26_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i89_LC_9_26_7  (
            .in0(N__23094),
            .in1(N__34465),
            .in2(_gnd_net_),
            .in3(N__28523),
            .lcout(data_in_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35357),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i65_LC_9_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i65_LC_9_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i65_LC_9_27_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i65_LC_9_27_0  (
            .in0(N__36814),
            .in1(N__36226),
            .in2(N__27772),
            .in3(N__29015),
            .lcout(\c0.data_in_field_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35365),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i41_LC_9_27_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i41_LC_9_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i41_LC_9_27_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i41_LC_9_27_1  (
            .in0(N__28046),
            .in1(N__34474),
            .in2(_gnd_net_),
            .in3(N__26861),
            .lcout(data_in_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35365),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i57_LC_9_27_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i57_LC_9_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i57_LC_9_27_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i57_LC_9_27_2  (
            .in0(N__27768),
            .in1(_gnd_net_),
            .in2(N__34546),
            .in3(N__30929),
            .lcout(data_in_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35365),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i49_LC_9_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i49_LC_9_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i49_LC_9_27_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_0___i49_LC_9_27_3  (
            .in0(N__30930),
            .in1(_gnd_net_),
            .in2(N__28050),
            .in3(N__34478),
            .lcout(data_in_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35365),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i107_LC_9_27_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i107_LC_9_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i107_LC_9_27_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i107_LC_9_27_4  (
            .in0(N__34473),
            .in1(N__29078),
            .in2(_gnd_net_),
            .in3(N__30699),
            .lcout(data_in_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35365),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i90_LC_9_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i90_LC_9_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i90_LC_9_27_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i90_LC_9_27_5  (
            .in0(N__36225),
            .in1(N__36815),
            .in2(N__28609),
            .in3(N__23535),
            .lcout(\c0.data_in_field_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35365),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_912_LC_9_27_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_912_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_912_LC_9_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_912_LC_9_27_6  (
            .in0(N__25763),
            .in1(N__27130),
            .in2(N__30672),
            .in3(N__23499),
            .lcout(\c0.n23_adj_1925 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5435_LC_9_27_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5435_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5435_LC_9_27_7 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5435_LC_9_27_7  (
            .in0(N__33263),
            .in1(N__23436),
            .in2(N__32678),
            .in3(N__31785),
            .lcout(\c0.n5797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_890_LC_9_28_0 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_890_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_890_LC_9_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_890_LC_9_28_0  (
            .in0(N__23379),
            .in1(N__31710),
            .in2(N__25080),
            .in3(N__24894),
            .lcout(\c0.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_955_LC_9_28_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_955_LC_9_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_955_LC_9_28_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_955_LC_9_28_1  (
            .in0(N__26150),
            .in1(N__23319),
            .in2(N__29399),
            .in3(N__27353),
            .lcout(\c0.n25_adj_1960 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i27_LC_9_28_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i27_LC_9_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i27_LC_9_28_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i27_LC_9_28_2  (
            .in0(N__29398),
            .in1(N__34532),
            .in2(_gnd_net_),
            .in3(N__30615),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i1_LC_9_28_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i1_LC_9_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i1_LC_9_28_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i1_LC_9_28_3  (
            .in0(N__34531),
            .in1(N__31417),
            .in2(_gnd_net_),
            .in3(N__27354),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_852_LC_9_28_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_852_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_852_LC_9_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_852_LC_9_28_4  (
            .in0(N__25367),
            .in1(N__29790),
            .in2(N__24836),
            .in3(N__23255),
            .lcout(\c0.n5093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i59_LC_9_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i59_LC_9_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i59_LC_9_28_5 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i59_LC_9_28_5  (
            .in0(N__36197),
            .in1(N__30001),
            .in2(N__37079),
            .in3(N__28294),
            .lcout(\c0.data_in_field_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i58_LC_9_28_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i58_LC_9_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i58_LC_9_28_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i58_LC_9_28_6  (
            .in0(N__34533),
            .in1(N__30297),
            .in2(_gnd_net_),
            .in3(N__23972),
            .lcout(data_in_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5510_LC_9_29_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5510_LC_9_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5510_LC_9_29_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5510_LC_9_29_0  (
            .in0(N__33298),
            .in1(N__23652),
            .in2(N__32666),
            .in3(N__23758),
            .lcout(\c0.n5881 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i30_LC_9_29_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i30_LC_9_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i30_LC_9_29_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i30_LC_9_29_2  (
            .in0(N__36034),
            .in1(N__36955),
            .in2(N__23656),
            .in3(N__27966),
            .lcout(\c0.data_in_field_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i143_LC_9_29_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i143_LC_9_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i143_LC_9_29_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i143_LC_9_29_3  (
            .in0(N__36954),
            .in1(N__36036),
            .in2(N__24184),
            .in3(N__27113),
            .lcout(\c0.data_in_field_142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i6_LC_9_29_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i6_LC_9_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i6_LC_9_29_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i6_LC_9_29_4  (
            .in0(N__36035),
            .in1(N__36956),
            .in2(N__27493),
            .in3(N__25526),
            .lcout(\c0.data_in_field_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i119_LC_9_29_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i119_LC_9_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i119_LC_9_29_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i119_LC_9_29_5  (
            .in0(N__34319),
            .in1(N__23691),
            .in2(_gnd_net_),
            .in3(N__28725),
            .lcout(data_in_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_988_LC_9_29_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_988_LC_9_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_988_LC_9_29_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_988_LC_9_29_6  (
            .in0(N__25652),
            .in1(N__23651),
            .in2(N__27126),
            .in3(N__23911),
            .lcout(\c0.n2046 ),
            .ltout(\c0.n2046_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_824_LC_9_29_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_824_LC_9_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_824_LC_9_29_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_824_LC_9_29_7  (
            .in0(N__23619),
            .in1(N__27370),
            .in2(N__23578),
            .in3(N__25392),
            .lcout(\c0.n5108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i50_LC_9_30_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i50_LC_9_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i50_LC_9_30_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i50_LC_9_30_0  (
            .in0(N__37148),
            .in1(N__35990),
            .in2(N__25997),
            .in3(N__23949),
            .lcout(\c0.data_in_field_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i50_LC_9_30_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i50_LC_9_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i50_LC_9_30_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i50_LC_9_30_1  (
            .in0(N__23948),
            .in1(N__34497),
            .in2(_gnd_net_),
            .in3(N__23979),
            .lcout(data_in_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i142_LC_9_30_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i142_LC_9_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i142_LC_9_30_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i142_LC_9_30_2  (
            .in0(N__37147),
            .in1(N__35989),
            .in2(N__24019),
            .in3(N__23920),
            .lcout(\c0.data_in_field_141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i15_LC_9_30_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i15_LC_9_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i15_LC_9_30_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i15_LC_9_30_3  (
            .in0(N__35986),
            .in1(N__23893),
            .in2(N__28509),
            .in3(N__37151),
            .lcout(\c0.data_in_field_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i48_LC_9_30_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i48_LC_9_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i48_LC_9_30_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i48_LC_9_30_4  (
            .in0(N__34495),
            .in1(N__27737),
            .in2(_gnd_net_),
            .in3(N__23802),
            .lcout(data_in_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i80_LC_9_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i80_LC_9_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i80_LC_9_30_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i80_LC_9_30_5  (
            .in0(N__35988),
            .in1(N__37150),
            .in2(N__25497),
            .in3(N__23844),
            .lcout(\c0.data_in_field_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i56_LC_9_30_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i56_LC_9_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i56_LC_9_30_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i56_LC_9_30_6  (
            .in0(N__34496),
            .in1(N__24114),
            .in2(_gnd_net_),
            .in3(N__23801),
            .lcout(data_in_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i38_LC_9_30_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i38_LC_9_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i38_LC_9_30_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i38_LC_9_30_7  (
            .in0(N__35987),
            .in1(N__37149),
            .in2(N__27802),
            .in3(N__25249),
            .lcout(\c0.data_in_field_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i18_LC_9_31_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i18_LC_9_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i18_LC_9_31_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i18_LC_9_31_0  (
            .in0(N__34493),
            .in1(N__30181),
            .in2(_gnd_net_),
            .in3(N__23787),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35392),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i122_LC_9_31_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i122_LC_9_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i122_LC_9_31_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i122_LC_9_31_1  (
            .in0(N__37143),
            .in1(N__36025),
            .in2(N__31168),
            .in3(N__24068),
            .lcout(\c0.data_in_field_121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35392),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i62_LC_9_31_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i62_LC_9_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i62_LC_9_31_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i62_LC_9_31_2  (
            .in0(N__36024),
            .in1(N__37146),
            .in2(N__25294),
            .in3(N__24250),
            .lcout(\c0.data_in_field_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35392),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i143_LC_9_31_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i143_LC_9_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i143_LC_9_31_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i143_LC_9_31_3  (
            .in0(N__34320),
            .in1(N__24170),
            .in2(_gnd_net_),
            .in3(N__24222),
            .lcout(data_in_17_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35392),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i6_LC_9_31_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i6_LC_9_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i6_LC_9_31_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i6_LC_9_31_4  (
            .in0(N__34494),
            .in1(N__24150),
            .in2(_gnd_net_),
            .in3(N__27488),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35392),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i64_LC_9_31_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i64_LC_9_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i64_LC_9_31_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i64_LC_9_31_5  (
            .in0(N__37144),
            .in1(N__36026),
            .in2(N__24118),
            .in3(N__26715),
            .lcout(\c0.data_in_field_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35392),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i2_LC_9_31_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i2_LC_9_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i2_LC_9_31_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0___i2_LC_9_31_6  (
            .in0(N__25836),
            .in1(N__37145),
            .in2(N__36204),
            .in3(N__29655),
            .lcout(\c0.data_in_field_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35392),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_822_LC_9_31_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_822_LC_9_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_822_LC_9_31_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_822_LC_9_31_7  (
            .in0(N__25282),
            .in1(N__24067),
            .in2(_gnd_net_),
            .in3(N__25835),
            .lcout(\c0.n1830 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i40_LC_9_32_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i40_LC_9_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i40_LC_9_32_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i40_LC_9_32_2  (
            .in0(N__34140),
            .in1(N__27744),
            .in2(_gnd_net_),
            .in3(N__25577),
            .lcout(data_in_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35398),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i32_LC_9_32_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i32_LC_9_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i32_LC_9_32_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i32_LC_9_32_3  (
            .in0(N__25578),
            .in1(N__34141),
            .in2(_gnd_net_),
            .in3(N__24043),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35398),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i33_LC_9_32_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i33_LC_9_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i33_LC_9_32_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i33_LC_9_32_4  (
            .in0(N__34139),
            .in1(N__26874),
            .in2(_gnd_net_),
            .in3(N__29151),
            .lcout(data_in_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35398),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i134_LC_9_32_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i134_LC_9_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i134_LC_9_32_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i134_LC_9_32_7  (
            .in0(N__34138),
            .in1(N__24015),
            .in2(_gnd_net_),
            .in3(N__24461),
            .lcout(data_in_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35398),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i147_LC_10_24_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i147_LC_10_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i147_LC_10_24_1 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \c0.data_in_0___i147_LC_10_24_1  (
            .in0(N__34545),
            .in1(N__24435),
            .in2(N__31237),
            .in3(_gnd_net_),
            .lcout(data_in_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i133_LC_10_24_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i133_LC_10_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i133_LC_10_24_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i133_LC_10_24_2  (
            .in0(N__34523),
            .in1(N__26764),
            .in2(_gnd_net_),
            .in3(N__28178),
            .lcout(data_in_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5425_LC_10_24_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5425_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5425_LC_10_24_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5425_LC_10_24_4  (
            .in0(N__33270),
            .in1(N__29374),
            .in2(N__32712),
            .in3(N__29217),
            .lcout(\c0.n5779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i105_LC_10_24_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i105_LC_10_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i105_LC_10_24_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i105_LC_10_24_5  (
            .in0(N__34544),
            .in1(N__24375),
            .in2(_gnd_net_),
            .in3(N__24363),
            .lcout(data_in_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i113_LC_10_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i113_LC_10_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i113_LC_10_24_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i113_LC_10_24_7  (
            .in0(N__36989),
            .in1(N__36205),
            .in2(N__24323),
            .in3(N__24364),
            .lcout(\c0.data_in_field_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i29_LC_10_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i29_LC_10_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i29_LC_10_25_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i29_LC_10_25_0  (
            .in0(N__24699),
            .in1(N__27928),
            .in2(N__37271),
            .in3(N__36207),
            .lcout(\c0.data_in_field_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35349),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_808_LC_10_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_808_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_808_LC_10_25_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_808_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(N__30529),
            .in2(_gnd_net_),
            .in3(N__24829),
            .lcout(\c0.n1929 ),
            .ltout(\c0.n1929_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_809_LC_10_25_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_809_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_809_LC_10_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_809_LC_10_25_2  (
            .in0(N__24316),
            .in1(N__32889),
            .in2(N__24286),
            .in3(N__28844),
            .lcout(),
            .ltout(\c0.n10_adj_1870_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_10_25_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_10_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_LC_10_25_3  (
            .in0(_gnd_net_),
            .in1(N__30916),
            .in2(N__24283),
            .in3(N__24697),
            .lcout(\c0.n5204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5485_LC_10_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5485_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5485_LC_10_25_4 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5485_LC_10_25_4  (
            .in0(N__24698),
            .in1(N__33315),
            .in2(N__32570),
            .in3(N__24682),
            .lcout(),
            .ltout(\c0.n5851_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5851_bdd_4_lut_LC_10_25_5 .C_ON=1'b0;
    defparam \c0.n5851_bdd_4_lut_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.n5851_bdd_4_lut_LC_10_25_5 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n5851_bdd_4_lut_LC_10_25_5  (
            .in0(N__28916),
            .in1(N__24639),
            .in2(N__24598),
            .in3(N__32475),
            .lcout(\c0.n5408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_984_LC_10_25_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_984_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_984_LC_10_25_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_984_LC_10_25_6  (
            .in0(N__26656),
            .in1(N__24887),
            .in2(_gnd_net_),
            .in3(N__27720),
            .lcout(\c0.n5267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i85_LC_10_25_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i85_LC_10_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i85_LC_10_25_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i85_LC_10_25_7  (
            .in0(N__36206),
            .in1(N__37218),
            .in2(N__26497),
            .in3(N__30530),
            .lcout(\c0.data_in_field_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35349),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5905_bdd_4_lut_LC_10_26_0 .C_ON=1'b0;
    defparam \c0.n5905_bdd_4_lut_LC_10_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.n5905_bdd_4_lut_LC_10_26_0 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n5905_bdd_4_lut_LC_10_26_0  (
            .in0(N__28959),
            .in1(N__32580),
            .in2(N__24550),
            .in3(N__25377),
            .lcout(\c0.n5381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_899_LC_10_26_1 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_899_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_899_LC_10_26_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_899_LC_10_26_1  (
            .in0(N__24535),
            .in1(N__31093),
            .in2(N__24524),
            .in3(N__26729),
            .lcout(\c0.n22_adj_1914 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i52_LC_10_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i52_LC_10_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i52_LC_10_26_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i52_LC_10_26_2  (
            .in0(N__37152),
            .in1(N__36208),
            .in2(N__26620),
            .in3(N__24932),
            .lcout(\c0.data_in_field_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i67_LC_10_26_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i67_LC_10_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i67_LC_10_26_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i67_LC_10_26_3  (
            .in0(N__30571),
            .in1(N__30721),
            .in2(N__36290),
            .in3(N__37153),
            .lcout(\c0.data_in_field_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_831_LC_10_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_831_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_831_LC_10_26_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_831_LC_10_26_4  (
            .in0(_gnd_net_),
            .in1(N__26655),
            .in2(_gnd_net_),
            .in3(N__24885),
            .lcout(),
            .ltout(\c0.n1947_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_10_26_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_10_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_LC_10_26_5  (
            .in0(N__25003),
            .in1(N__24909),
            .in2(N__24973),
            .in3(N__25311),
            .lcout(\c0.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_10_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_10_26_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_LC_10_26_6  (
            .in0(_gnd_net_),
            .in1(N__24931),
            .in2(_gnd_net_),
            .in3(N__30570),
            .lcout(\c0.n1922 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i76_LC_10_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i76_LC_10_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i76_LC_10_26_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i76_LC_10_26_7  (
            .in0(N__24886),
            .in1(N__26442),
            .in2(N__36291),
            .in3(N__37154),
            .lcout(\c0.data_in_field_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5707_bdd_4_lut_LC_10_27_1 .C_ON=1'b0;
    defparam \c0.n5707_bdd_4_lut_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5707_bdd_4_lut_LC_10_27_1 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n5707_bdd_4_lut_LC_10_27_1  (
            .in0(N__27340),
            .in1(N__32657),
            .in2(N__26914),
            .in3(N__30753),
            .lcout(\c0.n5474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_826_LC_10_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_826_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_826_LC_10_27_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_826_LC_10_27_2  (
            .in0(_gnd_net_),
            .in1(N__25185),
            .in2(_gnd_net_),
            .in3(N__25106),
            .lcout(\c0.n5105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_974_LC_10_27_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_974_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_974_LC_10_27_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_974_LC_10_27_3  (
            .in0(N__25107),
            .in1(N__26355),
            .in2(N__25196),
            .in3(N__28914),
            .lcout(\c0.n26_adj_1884 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i99_LC_10_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i99_LC_10_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i99_LC_10_27_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i99_LC_10_27_4  (
            .in0(N__36310),
            .in1(N__36806),
            .in2(N__29065),
            .in3(N__24828),
            .lcout(\c0.data_in_field_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35366),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i104_LC_10_27_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i104_LC_10_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i104_LC_10_27_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i104_LC_10_27_5  (
            .in0(N__36804),
            .in1(N__36311),
            .in2(N__24793),
            .in3(N__24739),
            .lcout(\c0.data_in_field_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35366),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i109_LC_10_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i109_LC_10_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i109_LC_10_27_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i109_LC_10_27_6  (
            .in0(N__36309),
            .in1(N__36805),
            .in2(N__26182),
            .in3(N__27179),
            .lcout(\c0.data_in_field_108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35366),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5500_LC_10_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5500_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5500_LC_10_28_0 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5500_LC_10_28_0  (
            .in0(N__33310),
            .in1(N__25192),
            .in2(N__32628),
            .in3(N__25293),
            .lcout(),
            .ltout(\c0.n5875_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5875_bdd_4_lut_LC_10_28_1 .C_ON=1'b0;
    defparam \c0.n5875_bdd_4_lut_LC_10_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5875_bdd_4_lut_LC_10_28_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5875_bdd_4_lut_LC_10_28_1  (
            .in0(N__32581),
            .in1(N__29607),
            .in2(N__25261),
            .in3(N__25258),
            .lcout(\c0.n5396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i54_LC_10_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i54_LC_10_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i54_LC_10_28_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i54_LC_10_28_2  (
            .in0(N__28108),
            .in1(N__36062),
            .in2(N__25200),
            .in3(N__37199),
            .lcout(\c0.data_in_field_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i44_LC_10_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i44_LC_10_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i44_LC_10_28_3 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i44_LC_10_28_3  (
            .in0(N__26574),
            .in1(N__36251),
            .in2(N__37267),
            .in3(N__25039),
            .lcout(\c0.data_in_field_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i125_LC_10_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i125_LC_10_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i125_LC_10_28_4 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i125_LC_10_28_4  (
            .in0(N__25105),
            .in1(N__37195),
            .in2(N__28162),
            .in3(N__36063),
            .lcout(\c0.data_in_field_124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_839_LC_10_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_839_LC_10_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_839_LC_10_28_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_839_LC_10_28_5  (
            .in0(_gnd_net_),
            .in1(N__25160),
            .in2(_gnd_net_),
            .in3(N__25104),
            .lcout(\c0.n1944 ),
            .ltout(\c0.n1944_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_864_LC_10_28_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_864_LC_10_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_864_LC_10_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_864_LC_10_28_6  (
            .in0(N__33394),
            .in1(N__31542),
            .in2(N__25063),
            .in3(N__28854),
            .lcout(),
            .ltout(\c0.n20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_865_LC_10_28_7 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_865_LC_10_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_865_LC_10_28_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_865_LC_10_28_7  (
            .in0(N__27381),
            .in1(N__28284),
            .in2(N__25060),
            .in3(N__25038),
            .lcout(\c0.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i78_LC_10_29_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i78_LC_10_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i78_LC_10_29_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i78_LC_10_29_0  (
            .in0(N__36085),
            .in1(N__37208),
            .in2(N__25451),
            .in3(N__27513),
            .lcout(\c0.data_in_field_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i40_LC_10_29_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i40_LC_10_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i40_LC_10_29_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i40_LC_10_29_1  (
            .in0(N__37207),
            .in1(N__36087),
            .in2(N__25588),
            .in3(N__25553),
            .lcout(\c0.data_in_field_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_814_LC_10_29_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_814_LC_10_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_814_LC_10_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_814_LC_10_29_2  (
            .in0(N__25552),
            .in1(N__25519),
            .in2(N__25491),
            .in3(N__28631),
            .lcout(),
            .ltout(\c0.n10_adj_1871_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_879_LC_10_29_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_879_LC_10_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_879_LC_10_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_879_LC_10_29_3  (
            .in0(N__25435),
            .in1(N__25870),
            .in2(N__25417),
            .in3(N__25365),
            .lcout(\c0.n5234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_10_29_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_10_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_10_29_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_LC_10_29_4  (
            .in0(N__28955),
            .in1(N__30451),
            .in2(N__28505),
            .in3(N__25780),
            .lcout(\c0.n1975 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i10_LC_10_29_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i10_LC_10_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i10_LC_10_29_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i10_LC_10_29_5  (
            .in0(N__30157),
            .in1(N__36086),
            .in2(N__37269),
            .in3(N__25871),
            .lcout(\c0.data_in_field_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i39_LC_10_29_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i39_LC_10_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i39_LC_10_29_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i39_LC_10_29_6  (
            .in0(N__25366),
            .in1(N__28078),
            .in2(N__36224),
            .in3(N__37212),
            .lcout(\c0.data_in_field_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i128_LC_10_29_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i128_LC_10_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i128_LC_10_29_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i128_LC_10_29_7  (
            .in0(N__25608),
            .in1(_gnd_net_),
            .in2(N__34547),
            .in3(N__27677),
            .lcout(data_in_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i98_LC_10_30_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i98_LC_10_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i98_LC_10_30_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i98_LC_10_30_0  (
            .in0(N__36230),
            .in1(N__37276),
            .in2(N__29795),
            .in3(N__25342),
            .lcout(\c0.data_in_field_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_807_LC_10_30_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_807_LC_10_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_807_LC_10_30_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_807_LC_10_30_1  (
            .in0(_gnd_net_),
            .in1(N__25691),
            .in2(_gnd_net_),
            .in3(N__27706),
            .lcout(\c0.n2062 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_823_LC_10_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_823_LC_10_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_823_LC_10_30_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_823_LC_10_30_2  (
            .in0(_gnd_net_),
            .in1(N__25749),
            .in2(_gnd_net_),
            .in3(N__25791),
            .lcout(\c0.n5141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i107_LC_10_30_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i107_LC_10_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i107_LC_10_30_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i107_LC_10_30_3  (
            .in0(N__37274),
            .in1(N__25759),
            .in2(N__29095),
            .in3(N__36235),
            .lcout(\c0.data_in_field_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i112_LC_10_30_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i112_LC_10_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i112_LC_10_30_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i112_LC_10_30_4  (
            .in0(N__25692),
            .in1(N__25726),
            .in2(N__36293),
            .in3(N__37277),
            .lcout(\c0.data_in_field_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i144_LC_10_30_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i144_LC_10_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i144_LC_10_30_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i144_LC_10_30_5  (
            .in0(N__37273),
            .in1(N__36231),
            .in2(N__25672),
            .in3(N__26020),
            .lcout(\c0.data_in_field_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i129_LC_10_30_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i129_LC_10_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i129_LC_10_30_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i129_LC_10_30_6  (
            .in0(N__36229),
            .in1(N__37275),
            .in2(N__27612),
            .in3(N__29515),
            .lcout(\c0.data_in_field_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i136_LC_10_30_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i136_LC_10_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i136_LC_10_30_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i136_LC_10_30_7  (
            .in0(N__34492),
            .in1(N__26019),
            .in2(_gnd_net_),
            .in3(N__25601),
            .lcout(data_in_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i3_LC_10_31_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i3_LC_10_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i3_LC_10_31_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i3_LC_10_31_0  (
            .in0(N__25911),
            .in1(N__35964),
            .in2(N__37289),
            .in3(N__27217),
            .lcout(\c0.data_in_field_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i101_LC_10_31_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i101_LC_10_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i101_LC_10_31_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i101_LC_10_31_1  (
            .in0(N__26178),
            .in1(N__34491),
            .in2(_gnd_net_),
            .in3(N__28685),
            .lcout(data_in_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i61_LC_10_31_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i61_LC_10_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i61_LC_10_31_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i61_LC_10_31_2  (
            .in0(N__37261),
            .in1(N__35965),
            .in2(N__34591),
            .in3(N__28003),
            .lcout(\c0.data_in_field_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i144_LC_10_31_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i144_LC_10_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i144_LC_10_31_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i144_LC_10_31_3  (
            .in0(N__34498),
            .in1(N__26018),
            .in2(_gnd_net_),
            .in3(N__26050),
            .lcout(data_in_17_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_828_LC_10_31_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_828_LC_10_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_828_LC_10_31_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_828_LC_10_31_4  (
            .in0(_gnd_net_),
            .in1(N__30100),
            .in2(_gnd_net_),
            .in3(N__26702),
            .lcout(),
            .ltout(\c0.n2092_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_836_LC_10_31_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_836_LC_10_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_836_LC_10_31_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_836_LC_10_31_5  (
            .in0(N__25981),
            .in1(N__27973),
            .in2(N__25960),
            .in3(N__25956),
            .lcout(\c0.n5246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i68_LC_10_31_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i68_LC_10_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i68_LC_10_31_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i68_LC_10_31_6  (
            .in0(N__34490),
            .in1(N__26443),
            .in2(_gnd_net_),
            .in3(N__33518),
            .lcout(data_in_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i52_LC_10_31_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i52_LC_10_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i52_LC_10_31_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i52_LC_10_31_7  (
            .in0(N__34499),
            .in1(N__26600),
            .in2(_gnd_net_),
            .in3(N__33501),
            .lcout(data_in_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35393),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i11_LC_10_32_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i11_LC_10_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i11_LC_10_32_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i11_LC_10_32_0  (
            .in0(N__33918),
            .in1(N__27455),
            .in2(_gnd_net_),
            .in3(N__29250),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35399),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i3_LC_10_32_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i3_LC_10_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i3_LC_10_32_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i3_LC_10_32_1  (
            .in0(N__27456),
            .in1(N__33921),
            .in2(_gnd_net_),
            .in3(N__25907),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35399),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i39_LC_10_32_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i39_LC_10_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i39_LC_10_32_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i39_LC_10_32_2  (
            .in0(N__33919),
            .in1(N__27240),
            .in2(_gnd_net_),
            .in3(N__28073),
            .lcout(data_in_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35399),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5749_bdd_4_lut_LC_10_32_4 .C_ON=1'b0;
    defparam \c0.n5749_bdd_4_lut_LC_10_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.n5749_bdd_4_lut_LC_10_32_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5749_bdd_4_lut_LC_10_32_4  (
            .in0(N__32733),
            .in1(N__25881),
            .in2(N__25852),
            .in3(N__25837),
            .lcout(\c0.n5453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i60_LC_10_32_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i60_LC_10_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i60_LC_10_32_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i60_LC_10_32_5  (
            .in0(N__37053),
            .in1(N__36312),
            .in2(N__26247),
            .in3(N__33505),
            .lcout(\c0.data_in_field_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35399),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i47_LC_10_32_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i47_LC_10_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i47_LC_10_32_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i47_LC_10_32_6  (
            .in0(N__33920),
            .in1(N__27239),
            .in2(_gnd_net_),
            .in3(N__26214),
            .lcout(data_in_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35399),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i63_LC_11_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i63_LC_11_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i63_LC_11_22_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i63_LC_11_22_4  (
            .in0(N__28131),
            .in1(_gnd_net_),
            .in2(N__34561),
            .in3(N__26510),
            .lcout(data_in_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i109_LC_11_22_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i109_LC_11_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i109_LC_11_22_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i109_LC_11_22_5  (
            .in0(N__31137),
            .in1(N__34553),
            .in2(_gnd_net_),
            .in3(N__26166),
            .lcout(data_in_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i91_LC_11_23_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i91_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i91_LC_11_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i91_LC_11_23_4  (
            .in0(N__34552),
            .in1(N__29055),
            .in2(_gnd_net_),
            .in3(N__31652),
            .lcout(data_in_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i21_LC_11_24_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i21_LC_11_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i21_LC_11_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i21_LC_11_24_0  (
            .in0(N__27926),
            .in1(N__26143),
            .in2(_gnd_net_),
            .in3(N__34560),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i116_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i116_LC_11_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i116_LC_11_24_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i116_LC_11_24_1  (
            .in0(N__34557),
            .in1(N__31371),
            .in2(_gnd_net_),
            .in3(N__31883),
            .lcout(data_in_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i71_LC_11_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i71_LC_11_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i71_LC_11_24_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i71_LC_11_24_2  (
            .in0(N__36222),
            .in1(N__36705),
            .in2(N__28132),
            .in3(N__32893),
            .lcout(\c0.data_in_field_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i116_LC_11_24_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i116_LC_11_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i116_LC_11_24_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i116_LC_11_24_3  (
            .in0(N__36704),
            .in1(N__36223),
            .in2(N__26091),
            .in3(N__31884),
            .lcout(\c0.data_in_field_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i66_LC_11_24_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i66_LC_11_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i66_LC_11_24_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i66_LC_11_24_6  (
            .in0(N__26538),
            .in1(N__34559),
            .in2(_gnd_net_),
            .in3(N__30284),
            .lcout(data_in_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i74_LC_11_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i74_LC_11_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i74_LC_11_24_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i74_LC_11_24_7  (
            .in0(N__34558),
            .in1(N__26537),
            .in2(_gnd_net_),
            .in3(N__28563),
            .lcout(data_in_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i63_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i63_LC_11_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i63_LC_11_25_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i63_LC_11_25_2  (
            .in0(N__36952),
            .in1(N__35863),
            .in2(N__26524),
            .in3(N__26663),
            .lcout(\c0.data_in_field_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35359),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i77_LC_11_25_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i77_LC_11_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i77_LC_11_25_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i77_LC_11_25_4  (
            .in0(N__34528),
            .in1(N__29702),
            .in2(_gnd_net_),
            .in3(N__26496),
            .lcout(data_in_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35359),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i84_LC_11_25_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i84_LC_11_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i84_LC_11_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i84_LC_11_25_6  (
            .in0(N__34529),
            .in1(N__31810),
            .in2(_gnd_net_),
            .in3(N__26456),
            .lcout(data_in_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35359),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i76_LC_11_25_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i76_LC_11_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i76_LC_11_25_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i76_LC_11_25_7  (
            .in0(N__26457),
            .in1(N__34530),
            .in2(_gnd_net_),
            .in3(N__26432),
            .lcout(data_in_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35359),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_11_26_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_11_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_LC_11_26_0  (
            .in0(N__28882),
            .in1(N__31946),
            .in2(N__26809),
            .in3(N__27178),
            .lcout(\c0.n26_adj_1878 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i5_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i5_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i5_LC_11_26_1 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i5_LC_11_26_1  (
            .in0(N__26404),
            .in1(N__36323),
            .in2(N__37086),
            .in3(N__28917),
            .lcout(\c0.data_in_field_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35367),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i69_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i69_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i69_LC_11_26_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i69_LC_11_26_2  (
            .in0(N__36322),
            .in1(N__36889),
            .in2(N__34617),
            .in3(N__26364),
            .lcout(\c0.data_in_field_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35367),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_926_LC_11_26_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_926_LC_11_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_926_LC_11_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_926_LC_11_26_3  (
            .in0(N__28867),
            .in1(N__27154),
            .in2(N__26329),
            .in3(N__26302),
            .lcout(\c0.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i87_LC_11_26_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i87_LC_11_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i87_LC_11_26_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i87_LC_11_26_4  (
            .in0(N__34526),
            .in1(N__31284),
            .in2(_gnd_net_),
            .in3(N__29957),
            .lcout(data_in_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35367),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i124_LC_11_26_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i124_LC_11_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i124_LC_11_26_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i124_LC_11_26_5  (
            .in0(N__31364),
            .in1(N__34527),
            .in2(_gnd_net_),
            .in3(N__26845),
            .lcout(data_in_15_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35367),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i141_LC_11_26_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i141_LC_11_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i141_LC_11_26_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_0___i141_LC_11_26_6  (
            .in0(N__26807),
            .in1(_gnd_net_),
            .in2(N__26763),
            .in3(N__34525),
            .lcout(data_in_17_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35367),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i141_LC_11_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i141_LC_11_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i141_LC_11_26_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i141_LC_11_26_7  (
            .in0(N__36888),
            .in1(N__26759),
            .in2(N__36331),
            .in3(N__28853),
            .lcout(\c0.data_in_field_140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35367),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_958_LC_11_27_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_958_LC_11_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_958_LC_11_27_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_958_LC_11_27_0  (
            .in0(N__26728),
            .in1(N__28975),
            .in2(N__30119),
            .in3(N__26664),
            .lcout(\c0.n1795 ),
            .ltout(\c0.n1795_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_114_2_lut_LC_11_27_1 .C_ON=1'b0;
    defparam \c0.i1_rep_114_2_lut_LC_11_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_114_2_lut_LC_11_27_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_rep_114_2_lut_LC_11_27_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26632),
            .in3(N__26894),
            .lcout(\c0.n6097 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i79_LC_11_27_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i79_LC_11_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i79_LC_11_27_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i79_LC_11_27_2  (
            .in0(N__32853),
            .in1(N__36807),
            .in2(N__29941),
            .in3(N__36327),
            .lcout(\c0.data_in_field_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35375),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_11_27_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_11_27_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_LC_11_27_3  (
            .in0(N__26930),
            .in1(N__26998),
            .in2(_gnd_net_),
            .in3(N__32852),
            .lcout(\c0.n5179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i44_LC_11_27_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i44_LC_11_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i44_LC_11_27_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i44_LC_11_27_4  (
            .in0(N__34524),
            .in1(N__26619),
            .in2(_gnd_net_),
            .in3(N__26570),
            .lcout(data_in_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35375),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_898_LC_11_27_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_898_LC_11_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_898_LC_11_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_898_LC_11_27_5  (
            .in0(N__27138),
            .in1(N__33393),
            .in2(N__27081),
            .in3(N__28849),
            .lcout(\c0.n11_adj_1913 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i93_LC_11_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i93_LC_11_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i93_LC_11_27_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i93_LC_11_27_6  (
            .in0(N__26999),
            .in1(N__27055),
            .in2(N__37005),
            .in3(N__36328),
            .lcout(\c0.data_in_field_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35375),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i94_LC_11_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i94_LC_11_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i94_LC_11_27_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i94_LC_11_27_7  (
            .in0(N__36329),
            .in1(N__26982),
            .in2(N__37004),
            .in3(N__26936),
            .lcout(\c0.data_in_field_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35375),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5375_LC_11_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5375_LC_11_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5375_LC_11_28_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5375_LC_11_28_0  (
            .in0(N__33256),
            .in1(N__31488),
            .in2(N__32679),
            .in3(N__29483),
            .lcout(\c0.n5707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i119_LC_11_28_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i119_LC_11_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i119_LC_11_28_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i119_LC_11_28_1  (
            .in0(N__36845),
            .in1(N__36083),
            .in2(N__28741),
            .in3(N__33398),
            .lcout(\c0.data_in_field_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35382),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i17_LC_11_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i17_LC_11_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i17_LC_11_28_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i17_LC_11_28_2  (
            .in0(N__36081),
            .in1(N__29484),
            .in2(N__31459),
            .in3(N__36848),
            .lcout(\c0.data_in_field_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35382),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_963_LC_11_28_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_963_LC_11_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_963_LC_11_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_963_LC_11_28_3  (
            .in0(N__28424),
            .in1(N__28714),
            .in2(N__28382),
            .in3(N__27150),
            .lcout(\c0.n1838 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i73_LC_11_28_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i73_LC_11_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i73_LC_11_28_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i73_LC_11_28_4  (
            .in0(N__36082),
            .in1(N__36847),
            .in2(N__29569),
            .in3(N__29457),
            .lcout(\c0.data_in_field_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35382),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i41_LC_11_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i41_LC_11_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i41_LC_11_28_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i41_LC_11_28_5  (
            .in0(N__36846),
            .in1(N__36084),
            .in2(N__26878),
            .in3(N__28635),
            .lcout(\c0.data_in_field_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35382),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_837_LC_11_28_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_837_LC_11_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_837_LC_11_28_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_837_LC_11_28_6  (
            .in0(_gnd_net_),
            .in1(N__29456),
            .in2(_gnd_net_),
            .in3(N__29794),
            .lcout(),
            .ltout(\c0.n6_adj_1876_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_838_LC_11_28_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_838_LC_11_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_838_LC_11_28_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_838_LC_11_28_7  (
            .in0(N__30450),
            .in1(N__30497),
            .in2(N__27436),
            .in3(N__27425),
            .lcout(\c0.n5129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_987_LC_11_29_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_987_LC_11_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_987_LC_11_29_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_987_LC_11_29_0  (
            .in0(N__27334),
            .in1(N__34667),
            .in2(_gnd_net_),
            .in3(N__34647),
            .lcout(\c0.n6_adj_1874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i1_LC_11_29_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i1_LC_11_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i1_LC_11_29_1 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i1_LC_11_29_1  (
            .in0(N__27361),
            .in1(N__36256),
            .in2(N__37270),
            .in3(N__27336),
            .lcout(\c0.data_in_field_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_999_LC_11_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_999_LC_11_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_999_LC_11_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_999_LC_11_29_2  (
            .in0(N__27335),
            .in1(N__27640),
            .in2(_gnd_net_),
            .in3(N__27311),
            .lcout(\c0.n22_adj_1935 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i35_LC_11_29_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i35_LC_11_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i35_LC_11_29_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i35_LC_11_29_4  (
            .in0(N__36255),
            .in1(N__37214),
            .in2(N__30616),
            .in3(N__28249),
            .lcout(\c0.data_in_field_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i47_LC_11_29_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i47_LC_11_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i47_LC_11_29_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i47_LC_11_29_5  (
            .in0(N__37213),
            .in1(N__36257),
            .in2(N__27250),
            .in3(N__28954),
            .lcout(\c0.data_in_field_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i25_LC_11_29_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i25_LC_11_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i25_LC_11_29_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i25_LC_11_29_6  (
            .in0(N__34406),
            .in1(N__29169),
            .in2(_gnd_net_),
            .in3(N__31513),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_815_LC_11_29_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_815_LC_11_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_815_LC_11_29_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_815_LC_11_29_7  (
            .in0(N__27218),
            .in1(N__27180),
            .in2(N__29284),
            .in3(N__29176),
            .lcout(\c0.n5102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i48_LC_11_30_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i48_LC_11_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i48_LC_11_30_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i48_LC_11_30_0  (
            .in0(N__37278),
            .in1(N__36254),
            .in2(N__27748),
            .in3(N__27713),
            .lcout(\c0.data_in_field_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i128_LC_11_30_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i128_LC_11_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i128_LC_11_30_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i128_LC_11_30_1  (
            .in0(N__36252),
            .in1(N__37279),
            .in2(N__27687),
            .in3(N__27641),
            .lcout(\c0.data_in_field_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i129_LC_11_30_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i129_LC_11_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i129_LC_11_30_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i129_LC_11_30_2  (
            .in0(N__34415),
            .in1(N__33432),
            .in2(_gnd_net_),
            .in3(N__27608),
            .lcout(data_in_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i16_LC_11_30_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i16_LC_11_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i16_LC_11_30_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i16_LC_11_30_3  (
            .in0(N__36253),
            .in1(N__27586),
            .in2(N__30353),
            .in3(N__37280),
            .lcout(\c0.data_in_field_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i29_LC_11_30_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i29_LC_11_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i29_LC_11_30_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i29_LC_11_30_4  (
            .in0(N__34416),
            .in1(N__30072),
            .in2(_gnd_net_),
            .in3(N__27919),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i78_LC_11_30_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i78_LC_11_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i78_LC_11_30_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i78_LC_11_30_5  (
            .in0(N__27546),
            .in1(N__34417),
            .in2(_gnd_net_),
            .in3(N__27509),
            .lcout(data_in_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i30_LC_11_30_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i30_LC_11_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i30_LC_11_30_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i30_LC_11_30_6  (
            .in0(N__27795),
            .in1(_gnd_net_),
            .in2(N__34535),
            .in3(N__27956),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i53_LC_11_30_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i53_LC_11_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i53_LC_11_30_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i53_LC_11_30_7  (
            .in0(N__34421),
            .in1(N__34587),
            .in2(_gnd_net_),
            .in3(N__30012),
            .lcout(data_in_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_LC_11_31_0 .C_ON=1'b0;
    defparam \c0.i6_2_lut_LC_11_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_LC_11_31_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i6_2_lut_LC_11_31_0  (
            .in0(N__27489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27454),
            .lcout(\c0.n22_adj_1952 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i46_LC_11_31_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i46_LC_11_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i46_LC_11_31_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i46_LC_11_31_1  (
            .in0(N__28107),
            .in1(_gnd_net_),
            .in2(N__34534),
            .in3(N__29624),
            .lcout(data_in_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35400),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i23_LC_11_31_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i23_LC_11_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i23_LC_11_31_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i23_LC_11_31_2  (
            .in0(N__27836),
            .in1(N__34408),
            .in2(_gnd_net_),
            .in3(N__27869),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35400),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i31_LC_11_31_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i31_LC_11_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i31_LC_11_31_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i31_LC_11_31_3  (
            .in0(N__34407),
            .in1(N__28074),
            .in2(_gnd_net_),
            .in3(N__27837),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35400),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i49_LC_11_31_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i49_LC_11_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i49_LC_11_31_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i49_LC_11_31_4  (
            .in0(N__37265),
            .in1(N__36101),
            .in2(N__30123),
            .in3(N__28057),
            .lcout(\c0.data_in_field_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35400),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_982_LC_11_31_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_982_LC_11_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_982_LC_11_31_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_982_LC_11_31_5  (
            .in0(N__29590),
            .in1(N__27994),
            .in2(_gnd_net_),
            .in3(N__30337),
            .lcout(\c0.n6_adj_1875 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_947_LC_11_31_6 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_947_LC_11_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_947_LC_11_31_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i12_4_lut_adj_947_LC_11_31_6  (
            .in0(N__31517),
            .in1(N__27949),
            .in2(N__27927),
            .in3(N__27868),
            .lcout(),
            .ltout(\c0.n28_adj_1953_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_953_LC_11_31_7 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_953_LC_11_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_953_LC_11_31_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_953_LC_11_31_7  (
            .in0(N__30185),
            .in1(N__27835),
            .in2(N__27820),
            .in3(N__27817),
            .lcout(\c0.n30_adj_1959 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i38_LC_11_32_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i38_LC_11_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i38_LC_11_32_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i38_LC_11_32_0  (
            .in0(N__33922),
            .in1(N__29625),
            .in2(_gnd_net_),
            .in3(N__27788),
            .lcout(data_in_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35405),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i65_LC_12_24_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i65_LC_12_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i65_LC_12_24_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i65_LC_12_24_4  (
            .in0(N__34538),
            .in1(N__29562),
            .in2(_gnd_net_),
            .in3(N__27759),
            .lcout(data_in_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35360),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5415_LC_12_24_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5415_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5415_LC_12_24_5 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5415_LC_12_24_5  (
            .in0(N__33271),
            .in1(N__28306),
            .in2(N__32627),
            .in3(N__30793),
            .lcout(),
            .ltout(\c0.n5773_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5773_bdd_4_lut_LC_12_24_6 .C_ON=1'b0;
    defparam \c0.n5773_bdd_4_lut_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.n5773_bdd_4_lut_LC_12_24_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5773_bdd_4_lut_LC_12_24_6  (
            .in0(N__32576),
            .in1(N__30448),
            .in2(N__28261),
            .in3(N__28258),
            .lcout(\c0.n5441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i117_LC_12_25_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i117_LC_12_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i117_LC_12_25_0 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_0___i117_LC_12_25_0  (
            .in0(_gnd_net_),
            .in1(N__28148),
            .in2(N__34536),
            .in3(N__31130),
            .lcout(data_in_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5701_bdd_4_lut_LC_12_25_1 .C_ON=1'b0;
    defparam \c0.n5701_bdd_4_lut_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5701_bdd_4_lut_LC_12_25_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5701_bdd_4_lut_LC_12_25_1  (
            .in0(N__32464),
            .in1(N__29129),
            .in2(N__30082),
            .in3(N__28636),
            .lcout(\c0.n5477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i123_LC_12_25_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i123_LC_12_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i123_LC_12_25_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i123_LC_12_25_2  (
            .in0(N__34428),
            .in1(N__33630),
            .in2(_gnd_net_),
            .in3(N__31967),
            .lcout(data_in_15_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i125_LC_12_25_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i125_LC_12_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i125_LC_12_25_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_0___i125_LC_12_25_3  (
            .in0(N__28188),
            .in1(_gnd_net_),
            .in2(N__28155),
            .in3(N__34429),
            .lcout(data_in_15_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i69_LC_12_25_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i69_LC_12_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i69_LC_12_25_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i69_LC_12_25_4  (
            .in0(N__29703),
            .in1(_gnd_net_),
            .in2(N__34537),
            .in3(N__34613),
            .lcout(data_in_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i71_LC_12_25_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i71_LC_12_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i71_LC_12_25_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i71_LC_12_25_5  (
            .in0(N__28130),
            .in1(N__29928),
            .in2(_gnd_net_),
            .in3(N__34430),
            .lcout(data_in_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i115_LC_12_25_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i115_LC_12_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i115_LC_12_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i115_LC_12_25_6  (
            .in0(N__34427),
            .in1(N__31968),
            .in2(_gnd_net_),
            .in3(N__30686),
            .lcout(data_in_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i82_LC_12_25_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i82_LC_12_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i82_LC_12_25_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i82_LC_12_25_7  (
            .in0(N__28562),
            .in1(N__28608),
            .in2(_gnd_net_),
            .in3(N__34431),
            .lcout(data_in_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i81_LC_12_26_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i81_LC_12_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i81_LC_12_26_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i81_LC_12_26_0  (
            .in0(N__34449),
            .in1(N__28536),
            .in2(_gnd_net_),
            .in3(N__29906),
            .lcout(data_in_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35376),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5911_bdd_4_lut_LC_12_26_1 .C_ON=1'b0;
    defparam \c0.n5911_bdd_4_lut_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5911_bdd_4_lut_LC_12_26_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n5911_bdd_4_lut_LC_12_26_1  (
            .in0(N__32659),
            .in1(N__28510),
            .in2(N__28480),
            .in3(N__28462),
            .lcout(\c0.n5378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_964_LC_12_26_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_964_LC_12_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_964_LC_12_26_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_964_LC_12_26_5  (
            .in0(N__29857),
            .in1(N__28366),
            .in2(_gnd_net_),
            .in3(N__28409),
            .lcout(\c0.n1899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i139_LC_12_26_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i139_LC_12_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i139_LC_12_26_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i139_LC_12_26_6  (
            .in0(N__28410),
            .in1(N__33658),
            .in2(N__36313),
            .in3(N__36894),
            .lcout(\c0.data_in_field_138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35376),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i131_LC_12_26_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i131_LC_12_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i131_LC_12_26_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i131_LC_12_26_7  (
            .in0(N__36893),
            .in1(N__36266),
            .in2(N__33634),
            .in3(N__28367),
            .lcout(\c0.data_in_field_130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35376),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_812_LC_12_27_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_812_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_812_LC_12_27_0 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_812_LC_12_27_0  (
            .in0(N__30259),
            .in1(_gnd_net_),
            .in2(N__30787),
            .in3(_gnd_net_),
            .lcout(\c0.n5123 ),
            .ltout(\c0.n5123_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_991_LC_12_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_991_LC_12_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_991_LC_12_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_991_LC_12_27_1  (
            .in0(N__28974),
            .in1(N__29029),
            .in2(N__28336),
            .in3(N__29437),
            .lcout(\c0.n5231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_813_LC_12_27_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_813_LC_12_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_813_LC_12_27_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_813_LC_12_27_2  (
            .in0(_gnd_net_),
            .in1(N__31480),
            .in2(_gnd_net_),
            .in3(N__30742),
            .lcout(\c0.n5188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i99_LC_12_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i99_LC_12_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i99_LC_12_27_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i99_LC_12_27_3  (
            .in0(N__34541),
            .in1(N__29091),
            .in2(_gnd_net_),
            .in3(N__29043),
            .lcout(data_in_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35383),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_12_27_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_12_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_12_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_12_27_4  (
            .in0(N__30258),
            .in1(N__29019),
            .in2(N__30788),
            .in3(N__28973),
            .lcout(),
            .ltout(\c0.n1767_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_994_LC_12_27_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_994_LC_12_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_994_LC_12_27_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_994_LC_12_27_5  (
            .in0(N__28960),
            .in1(N__28915),
            .in2(N__28885),
            .in3(N__28878),
            .lcout(\c0.n5126 ),
            .ltout(\c0.n5126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_884_LC_12_27_6 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_884_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_884_LC_12_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_884_LC_12_27_6  (
            .in0(N__28848),
            .in1(N__31083),
            .in2(N__28813),
            .in3(N__28808),
            .lcout(\c0.n20_adj_1899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i111_LC_12_28_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i111_LC_12_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i111_LC_12_28_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i111_LC_12_28_0  (
            .in0(N__34549),
            .in1(N__28737),
            .in2(_gnd_net_),
            .in3(N__29837),
            .lcout(data_in_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_816_LC_12_28_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_816_LC_12_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_816_LC_12_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_816_LC_12_28_1  (
            .in0(N__31575),
            .in1(N__31330),
            .in2(N__31932),
            .in3(N__28654),
            .lcout(\c0.n10_adj_1872 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i101_LC_12_28_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i101_LC_12_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i101_LC_12_28_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i101_LC_12_28_2  (
            .in0(N__36171),
            .in1(N__37167),
            .in2(N__28707),
            .in3(N__28665),
            .lcout(\c0.data_in_field_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_841_LC_12_28_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_841_LC_12_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_841_LC_12_28_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_841_LC_12_28_3  (
            .in0(_gnd_net_),
            .in1(N__28655),
            .in2(_gnd_net_),
            .in3(N__28630),
            .lcout(\c0.n1969 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i103_LC_12_28_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i103_LC_12_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i103_LC_12_28_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i103_LC_12_28_4  (
            .in0(N__34548),
            .in1(N__31299),
            .in2(_gnd_net_),
            .in3(N__29838),
            .lcout(data_in_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_LC_12_28_5 .C_ON=1'b0;
    defparam \c0.i2_4_lut_LC_12_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_LC_12_28_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_LC_12_28_5  (
            .in0(N__29527),
            .in1(N__31999),
            .in2(N__29488),
            .in3(N__29455),
            .lcout(\c0.n5138 ),
            .ltout(\c0.n5138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_992_LC_12_28_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_992_LC_12_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_992_LC_12_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_992_LC_12_28_6  (
            .in0(N__29361),
            .in1(N__29436),
            .in2(N__29425),
            .in3(N__32162),
            .lcout(\c0.n15_adj_1968 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i27_LC_12_28_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i27_LC_12_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i27_LC_12_28_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i27_LC_12_28_7  (
            .in0(N__29365),
            .in1(N__29413),
            .in2(N__37250),
            .in3(N__36170),
            .lcout(\c0.data_in_field_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i34_LC_12_29_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i34_LC_12_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i34_LC_12_29_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i34_LC_12_29_0  (
            .in0(N__37054),
            .in1(N__36163),
            .in2(N__29298),
            .in3(N__29334),
            .lcout(\c0.data_in_field_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35395),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i19_LC_12_29_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i19_LC_12_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i19_LC_12_29_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i19_LC_12_29_2  (
            .in0(N__29195),
            .in1(N__37060),
            .in2(N__29257),
            .in3(N__36202),
            .lcout(\c0.data_in_field_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35395),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_868_LC_12_29_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_868_LC_12_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_868_LC_12_29_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_868_LC_12_29_3  (
            .in0(N__31693),
            .in1(N__29194),
            .in2(_gnd_net_),
            .in3(N__29113),
            .lcout(\c0.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i33_LC_12_29_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i33_LC_12_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i33_LC_12_29_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i33_LC_12_29_4  (
            .in0(N__29114),
            .in1(N__29170),
            .in2(N__37194),
            .in3(N__36203),
            .lcout(\c0.data_in_field_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35395),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_844_LC_12_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_844_LC_12_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_844_LC_12_29_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_844_LC_12_29_5  (
            .in0(N__29674),
            .in1(N__31184),
            .in2(_gnd_net_),
            .in3(N__31767),
            .lcout(\c0.n5219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i111_LC_12_29_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i111_LC_12_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i111_LC_12_29_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i111_LC_12_29_7  (
            .in0(N__37059),
            .in1(N__29839),
            .in2(N__36270),
            .in3(N__32166),
            .lcout(\c0.data_in_field_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35395),
            .ce(),
            .sr(_gnd_net_));
    defparam i4988_4_lut_LC_12_30_0.C_ON=1'b0;
    defparam i4988_4_lut_LC_12_30_0.SEQ_MODE=4'b0000;
    defparam i4988_4_lut_LC_12_30_0.LUT_INIT=16'b1111111011000100;
    LogicCell40 i4988_4_lut_LC_12_30_0 (
            .in0(N__37438),
            .in1(N__37413),
            .in2(N__37387),
            .in3(N__37462),
            .lcout(n5332),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4987_4_lut_LC_12_30_1.C_ON=1'b0;
    defparam i4987_4_lut_LC_12_30_1.SEQ_MODE=4'b0000;
    defparam i4987_4_lut_LC_12_30_1.LUT_INIT=16'b1011101000100010;
    LogicCell40 i4987_4_lut_LC_12_30_1 (
            .in0(N__37461),
            .in1(N__37383),
            .in2(N__37414),
            .in3(N__37437),
            .lcout(),
            .ltout(n5331_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4989_3_lut_LC_12_30_2.C_ON=1'b0;
    defparam i4989_3_lut_LC_12_30_2.SEQ_MODE=4'b0000;
    defparam i4989_3_lut_LC_12_30_2.LUT_INIT=16'b0011001100001111;
    LogicCell40 i4989_3_lut_LC_12_30_2 (
            .in0(_gnd_net_),
            .in1(N__29824),
            .in2(N__29818),
            .in3(N__37357),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_12_30_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_12_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_12_30_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_12_30_3  (
            .in0(N__29675),
            .in1(N__31768),
            .in2(_gnd_net_),
            .in3(N__29786),
            .lcout(\c0.n1972 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i77_LC_12_30_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i77_LC_12_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i77_LC_12_30_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i77_LC_12_30_4  (
            .in0(N__37058),
            .in1(N__36174),
            .in2(N__29713),
            .in3(N__29676),
            .lcout(\c0.data_in_field_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35401),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i2_LC_12_31_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i2_LC_12_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i2_LC_12_31_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i2_LC_12_31_0  (
            .in0(N__34413),
            .in1(N__30149),
            .in2(_gnd_net_),
            .in3(N__29645),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35406),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i46_LC_12_31_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i46_LC_12_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i46_LC_12_31_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i46_LC_12_31_1  (
            .in0(N__37188),
            .in1(N__35966),
            .in2(N__29629),
            .in3(N__29597),
            .lcout(\c0.data_in_field_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35406),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i73_LC_12_31_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i73_LC_12_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i73_LC_12_31_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i73_LC_12_31_2  (
            .in0(N__34414),
            .in1(N__29550),
            .in2(_gnd_net_),
            .in3(N__29911),
            .lcout(data_in_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35406),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i10_LC_12_31_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i10_LC_12_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i10_LC_12_31_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i10_LC_12_31_6  (
            .in0(N__34412),
            .in1(N__30186),
            .in2(_gnd_net_),
            .in3(N__30148),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35406),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i51_LC_13_24_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i51_LC_13_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i51_LC_13_24_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i51_LC_13_24_1  (
            .in0(N__34540),
            .in1(N__30806),
            .in2(_gnd_net_),
            .in3(N__29994),
            .lcout(data_in_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35369),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i43_LC_13_24_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i43_LC_13_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i43_LC_13_24_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i43_LC_13_24_5  (
            .in0(N__34539),
            .in1(N__30807),
            .in2(_gnd_net_),
            .in3(N__30462),
            .lcout(data_in_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35369),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5356_LC_13_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5356_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5356_LC_13_25_0 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5356_LC_13_25_0  (
            .in0(N__33299),
            .in1(N__30915),
            .in2(N__30127),
            .in3(N__32465),
            .lcout(\c0.n5701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i37_LC_13_25_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i37_LC_13_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i37_LC_13_25_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i37_LC_13_25_1  (
            .in0(N__31599),
            .in1(N__34425),
            .in2(_gnd_net_),
            .in3(N__30053),
            .lcout(data_in_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i45_LC_13_25_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i45_LC_13_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i45_LC_13_25_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i45_LC_13_25_2  (
            .in0(N__34422),
            .in1(N__31598),
            .in2(_gnd_net_),
            .in3(N__30030),
            .lcout(data_in_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i59_LC_13_25_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i59_LC_13_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i59_LC_13_25_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i59_LC_13_25_3  (
            .in0(N__30714),
            .in1(N__34426),
            .in2(_gnd_net_),
            .in3(N__29993),
            .lcout(data_in_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i79_LC_13_25_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i79_LC_13_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i79_LC_13_25_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i79_LC_13_25_4  (
            .in0(N__34424),
            .in1(N__29927),
            .in2(_gnd_net_),
            .in3(N__29970),
            .lcout(data_in_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i81_LC_13_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i81_LC_13_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i81_LC_13_25_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i81_LC_13_25_5  (
            .in0(N__37009),
            .in1(N__35864),
            .in2(N__29875),
            .in3(N__29910),
            .lcout(\c0.data_in_field_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i67_LC_13_25_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i67_LC_13_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i67_LC_13_25_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i67_LC_13_25_6  (
            .in0(N__34423),
            .in1(N__33558),
            .in2(_gnd_net_),
            .in3(N__30713),
            .lcout(data_in_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i115_LC_13_26_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i115_LC_13_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i115_LC_13_26_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i115_LC_13_26_0  (
            .in0(N__37006),
            .in1(N__36265),
            .in2(N__30700),
            .in3(N__30648),
            .lcout(\c0.data_in_field_114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i35_LC_13_26_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i35_LC_13_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i35_LC_13_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i35_LC_13_26_1  (
            .in0(N__34448),
            .in1(N__30468),
            .in2(_gnd_net_),
            .in3(N__30596),
            .lcout(data_in_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_13_26_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_13_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_LC_13_26_2  (
            .in0(N__32010),
            .in1(N__30579),
            .in2(N__30547),
            .in3(N__30504),
            .lcout(\c0.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i43_LC_13_26_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i43_LC_13_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i43_LC_13_26_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i43_LC_13_26_3  (
            .in0(N__36263),
            .in1(N__37007),
            .in2(N__30449),
            .in3(N__30469),
            .lcout(\c0.data_in_field_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_976_LC_13_26_4 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_976_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_976_LC_13_26_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_976_LC_13_26_4  (
            .in0(N__30886),
            .in1(N__31936),
            .in2(N__30409),
            .in3(N__30354),
            .lcout(\c0.n20_adj_1916 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i66_LC_13_26_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i66_LC_13_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i66_LC_13_26_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i66_LC_13_26_5  (
            .in0(N__36264),
            .in1(N__37008),
            .in2(N__30301),
            .in3(N__30257),
            .lcout(\c0.data_in_field_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i122_LC_13_26_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i122_LC_13_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i122_LC_13_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i122_LC_13_26_6  (
            .in0(N__34446),
            .in1(N__30216),
            .in2(_gnd_net_),
            .in3(N__31154),
            .lcout(data_in_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i114_LC_13_26_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i114_LC_13_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i114_LC_13_26_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i114_LC_13_26_7  (
            .in0(N__31155),
            .in1(N__34447),
            .in2(_gnd_net_),
            .in3(N__30992),
            .lcout(data_in_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i117_LC_13_27_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i117_LC_13_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i117_LC_13_27_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i117_LC_13_27_0  (
            .in0(N__31107),
            .in1(N__37189),
            .in2(N__31141),
            .in3(N__36217),
            .lcout(\c0.data_in_field_116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35390),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_842_LC_13_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_842_LC_13_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_842_LC_13_27_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_842_LC_13_27_1  (
            .in0(_gnd_net_),
            .in1(N__31106),
            .in2(_gnd_net_),
            .in3(N__32960),
            .lcout(\c0.n1815 ),
            .ltout(\c0.n1815_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_13_27_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_13_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_LC_13_27_2  (
            .in0(N__30907),
            .in1(N__31481),
            .in2(N__31072),
            .in3(N__31068),
            .lcout(\c0.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i106_LC_13_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i106_LC_13_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i106_LC_13_27_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i106_LC_13_27_3  (
            .in0(N__34542),
            .in1(N__30956),
            .in2(_gnd_net_),
            .in3(N__30999),
            .lcout(data_in_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35390),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i57_LC_13_27_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i57_LC_13_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i57_LC_13_27_4 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i57_LC_13_27_4  (
            .in0(N__30908),
            .in1(N__37190),
            .in2(N__30940),
            .in3(N__36218),
            .lcout(\c0.data_in_field_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35390),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_910_LC_13_27_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_910_LC_13_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_910_LC_13_27_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_910_LC_13_27_5  (
            .in0(_gnd_net_),
            .in1(N__31247),
            .in2(_gnd_net_),
            .in3(N__30885),
            .lcout(\c0.n15_adj_1923 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i51_LC_13_27_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i51_LC_13_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i51_LC_13_27_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i51_LC_13_27_6  (
            .in0(N__30814),
            .in1(N__36216),
            .in2(N__30792),
            .in3(N__36803),
            .lcout(\c0.data_in_field_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35390),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i9_LC_13_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i9_LC_13_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i9_LC_13_27_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i9_LC_13_27_7  (
            .in0(N__36215),
            .in1(N__36802),
            .in2(N__31409),
            .in3(N__30749),
            .lcout(\c0.data_in_field_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35390),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i103_LC_13_28_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i103_LC_13_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i103_LC_13_28_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i103_LC_13_28_0  (
            .in0(N__37184),
            .in1(N__36162),
            .in2(N__32829),
            .in3(N__31306),
            .lcout(\c0.data_in_field_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35396),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i45_LC_13_28_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i45_LC_13_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i45_LC_13_28_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i45_LC_13_28_1  (
            .in0(N__36161),
            .in1(N__37186),
            .in2(N__31609),
            .in3(N__31574),
            .lcout(\c0.data_in_field_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35396),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_840_LC_13_28_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_840_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_840_LC_13_28_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_840_LC_13_28_2  (
            .in0(_gnd_net_),
            .in1(N__32809),
            .in2(_gnd_net_),
            .in3(N__32161),
            .lcout(\c0.n1962 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i25_LC_13_28_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i25_LC_13_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i25_LC_13_28_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i25_LC_13_28_3  (
            .in0(N__36160),
            .in1(N__31524),
            .in2(N__31489),
            .in3(N__37187),
            .lcout(\c0.data_in_field_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35396),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i9_LC_13_28_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i9_LC_13_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i9_LC_13_28_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i9_LC_13_28_4  (
            .in0(N__31402),
            .in1(N__31458),
            .in2(_gnd_net_),
            .in3(N__34451),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35396),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i124_LC_13_28_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i124_LC_13_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i124_LC_13_28_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i124_LC_13_28_5  (
            .in0(N__36159),
            .in1(N__37185),
            .in2(N__31378),
            .in3(N__31331),
            .lcout(\c0.data_in_field_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35396),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i95_LC_13_28_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i95_LC_13_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i95_LC_13_28_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i95_LC_13_28_6  (
            .in0(N__34550),
            .in1(N__31305),
            .in2(_gnd_net_),
            .in3(N__31274),
            .lcout(data_in_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35396),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i139_LC_13_28_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i139_LC_13_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i139_LC_13_28_7 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \c0.data_in_0___i139_LC_13_28_7  (
            .in0(N__34450),
            .in1(N__33650),
            .in2(N__31252),
            .in3(_gnd_net_),
            .lcout(data_in_17_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35396),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i75_LC_13_29_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i75_LC_13_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i75_LC_13_29_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i75_LC_13_29_0  (
            .in0(N__31190),
            .in1(N__36168),
            .in2(N__33559),
            .in3(N__37163),
            .lcout(\c0.data_in_field_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i137_LC_13_29_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i137_LC_13_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i137_LC_13_29_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i137_LC_13_29_1  (
            .in0(N__37165),
            .in1(N__36172),
            .in2(N__33433),
            .in3(N__32006),
            .lcout(\c0.data_in_field_136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i123_LC_13_29_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i123_LC_13_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i123_LC_13_29_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i123_LC_13_29_2  (
            .in0(N__31931),
            .in1(N__36167),
            .in2(N__31978),
            .in3(N__37162),
            .lcout(\c0.data_in_field_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i108_LC_13_29_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i108_LC_13_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i108_LC_13_29_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i108_LC_13_29_3  (
            .in0(N__34500),
            .in1(N__31853),
            .in2(_gnd_net_),
            .in3(N__31894),
            .lcout(data_in_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i100_LC_13_29_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i100_LC_13_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i100_LC_13_29_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i100_LC_13_29_4  (
            .in0(N__31854),
            .in1(N__34501),
            .in2(_gnd_net_),
            .in3(N__31823),
            .lcout(data_in_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i92_LC_13_29_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i92_LC_13_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i92_LC_13_29_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i92_LC_13_29_5  (
            .in0(N__31824),
            .in1(_gnd_net_),
            .in2(N__34551),
            .in3(N__31799),
            .lcout(data_in_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i92_LC_13_29_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i92_LC_13_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i92_LC_13_29_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i92_LC_13_29_6  (
            .in0(N__31775),
            .in1(N__36169),
            .in2(N__31806),
            .in3(N__37164),
            .lcout(\c0.data_in_field_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i4_LC_13_29_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i4_LC_13_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i4_LC_13_29_7 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i4_LC_13_29_7  (
            .in0(N__37166),
            .in1(N__31744),
            .in2(N__31709),
            .in3(N__36173),
            .lcout(\c0.data_in_field_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35402),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i83_LC_13_30_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i83_LC_13_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i83_LC_13_30_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i83_LC_13_30_0  (
            .in0(N__34281),
            .in1(N__31671),
            .in2(_gnd_net_),
            .in3(N__31622),
            .lcout(data_in_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35407),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i75_LC_13_30_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i75_LC_13_30_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i75_LC_13_30_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i75_LC_13_30_2  (
            .in0(N__34280),
            .in1(N__33551),
            .in2(_gnd_net_),
            .in3(N__31623),
            .lcout(data_in_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35407),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i60_LC_13_30_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i60_LC_13_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i60_LC_13_30_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i60_LC_13_30_6  (
            .in0(N__34279),
            .in1(N__33531),
            .in2(_gnd_net_),
            .in3(N__33489),
            .lcout(data_in_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35407),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i137_LC_13_31_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i137_LC_13_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i137_LC_13_31_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i137_LC_13_31_1  (
            .in0(N__34278),
            .in1(N__33419),
            .in2(_gnd_net_),
            .in3(N__33478),
            .lcout(data_in_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35410),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5515_LC_14_25_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5515_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5515_LC_14_25_1 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5515_LC_14_25_1  (
            .in0(N__33316),
            .in1(N__33402),
            .in2(N__32564),
            .in3(N__33361),
            .lcout(\c0.n5893 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5520_LC_14_26_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5520_LC_14_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5520_LC_14_26_0 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5520_LC_14_26_0  (
            .in0(N__33311),
            .in1(N__33001),
            .in2(N__32658),
            .in3(N__32965),
            .lcout(),
            .ltout(\c0.n5899_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5899_bdd_4_lut_LC_14_26_1 .C_ON=1'b0;
    defparam \c0.n5899_bdd_4_lut_LC_14_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5899_bdd_4_lut_LC_14_26_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5899_bdd_4_lut_LC_14_26_1  (
            .in0(N__32713),
            .in1(N__32909),
            .in2(N__32863),
            .in3(N__32860),
            .lcout(\c0.n5384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5893_bdd_4_lut_LC_14_26_3 .C_ON=1'b0;
    defparam \c0.n5893_bdd_4_lut_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5893_bdd_4_lut_LC_14_26_3 .LUT_INIT=16'b1010111010100100;
    LogicCell40 \c0.n5893_bdd_4_lut_LC_14_26_3  (
            .in0(N__32839),
            .in1(N__32825),
            .in2(N__32734),
            .in3(N__32170),
            .lcout(),
            .ltout(\c0.n5387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_14_26_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_14_26_4 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_LC_14_26_4  (
            .in0(N__34830),
            .in1(N__32140),
            .in2(N__32134),
            .in3(N__32131),
            .lcout(),
            .ltout(\c0.n5887_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5887_bdd_4_lut_LC_14_26_5 .C_ON=1'b0;
    defparam \c0.n5887_bdd_4_lut_LC_14_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.n5887_bdd_4_lut_LC_14_26_5 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n5887_bdd_4_lut_LC_14_26_5  (
            .in0(N__32047),
            .in1(N__32038),
            .in2(N__34834),
            .in3(N__34831),
            .lcout(\c0.n5890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_817_LC_14_28_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_817_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_817_LC_14_28_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_817_LC_14_28_2  (
            .in0(_gnd_net_),
            .in1(N__34680),
            .in2(_gnd_net_),
            .in3(N__34651),
            .lcout(\c0.n1896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i61_LC_14_28_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i61_LC_14_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i61_LC_14_28_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i61_LC_14_28_3  (
            .in0(N__34459),
            .in1(N__34618),
            .in2(_gnd_net_),
            .in3(N__34572),
            .lcout(data_in_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i131_LC_14_28_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i131_LC_14_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i131_LC_14_28_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i131_LC_14_28_5  (
            .in0(N__34458),
            .in1(N__33651),
            .in2(_gnd_net_),
            .in3(N__33615),
            .lcout(data_in_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35403),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i0_LC_15_25_0.C_ON=1'b1;
    defparam blink_counter_523__i0_LC_15_25_0.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i0_LC_15_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i0_LC_15_25_0 (
            .in0(_gnd_net_),
            .in1(N__33604),
            .in2(_gnd_net_),
            .in3(N__33598),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(n4437),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i1_LC_15_25_1.C_ON=1'b1;
    defparam blink_counter_523__i1_LC_15_25_1.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i1_LC_15_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i1_LC_15_25_1 (
            .in0(_gnd_net_),
            .in1(N__33595),
            .in2(_gnd_net_),
            .in3(N__33589),
            .lcout(n25),
            .ltout(),
            .carryin(n4437),
            .carryout(n4438),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i2_LC_15_25_2.C_ON=1'b1;
    defparam blink_counter_523__i2_LC_15_25_2.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i2_LC_15_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i2_LC_15_25_2 (
            .in0(_gnd_net_),
            .in1(N__33586),
            .in2(_gnd_net_),
            .in3(N__33580),
            .lcout(n24),
            .ltout(),
            .carryin(n4438),
            .carryout(n4439),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i3_LC_15_25_3.C_ON=1'b1;
    defparam blink_counter_523__i3_LC_15_25_3.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i3_LC_15_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i3_LC_15_25_3 (
            .in0(_gnd_net_),
            .in1(N__33577),
            .in2(_gnd_net_),
            .in3(N__33571),
            .lcout(n23),
            .ltout(),
            .carryin(n4439),
            .carryout(n4440),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i4_LC_15_25_4.C_ON=1'b1;
    defparam blink_counter_523__i4_LC_15_25_4.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i4_LC_15_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i4_LC_15_25_4 (
            .in0(_gnd_net_),
            .in1(N__33568),
            .in2(_gnd_net_),
            .in3(N__33562),
            .lcout(n22),
            .ltout(),
            .carryin(n4440),
            .carryout(n4441),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i5_LC_15_25_5.C_ON=1'b1;
    defparam blink_counter_523__i5_LC_15_25_5.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i5_LC_15_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i5_LC_15_25_5 (
            .in0(_gnd_net_),
            .in1(N__34906),
            .in2(_gnd_net_),
            .in3(N__34900),
            .lcout(n21),
            .ltout(),
            .carryin(n4441),
            .carryout(n4442),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i6_LC_15_25_6.C_ON=1'b1;
    defparam blink_counter_523__i6_LC_15_25_6.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i6_LC_15_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i6_LC_15_25_6 (
            .in0(_gnd_net_),
            .in1(N__34897),
            .in2(_gnd_net_),
            .in3(N__34891),
            .lcout(n20),
            .ltout(),
            .carryin(n4442),
            .carryout(n4443),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i7_LC_15_25_7.C_ON=1'b1;
    defparam blink_counter_523__i7_LC_15_25_7.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i7_LC_15_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i7_LC_15_25_7 (
            .in0(_gnd_net_),
            .in1(N__34888),
            .in2(_gnd_net_),
            .in3(N__34882),
            .lcout(n19),
            .ltout(),
            .carryin(n4443),
            .carryout(n4444),
            .clk(N__35391),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i8_LC_15_26_0.C_ON=1'b1;
    defparam blink_counter_523__i8_LC_15_26_0.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i8_LC_15_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i8_LC_15_26_0 (
            .in0(_gnd_net_),
            .in1(N__34879),
            .in2(_gnd_net_),
            .in3(N__34873),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(n4445),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i9_LC_15_26_1.C_ON=1'b1;
    defparam blink_counter_523__i9_LC_15_26_1.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i9_LC_15_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i9_LC_15_26_1 (
            .in0(_gnd_net_),
            .in1(N__34870),
            .in2(_gnd_net_),
            .in3(N__34864),
            .lcout(n17),
            .ltout(),
            .carryin(n4445),
            .carryout(n4446),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i10_LC_15_26_2.C_ON=1'b1;
    defparam blink_counter_523__i10_LC_15_26_2.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i10_LC_15_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i10_LC_15_26_2 (
            .in0(_gnd_net_),
            .in1(N__34861),
            .in2(_gnd_net_),
            .in3(N__34855),
            .lcout(n16),
            .ltout(),
            .carryin(n4446),
            .carryout(n4447),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i11_LC_15_26_3.C_ON=1'b1;
    defparam blink_counter_523__i11_LC_15_26_3.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i11_LC_15_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i11_LC_15_26_3 (
            .in0(_gnd_net_),
            .in1(N__34852),
            .in2(_gnd_net_),
            .in3(N__34846),
            .lcout(n15),
            .ltout(),
            .carryin(n4447),
            .carryout(n4448),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i12_LC_15_26_4.C_ON=1'b1;
    defparam blink_counter_523__i12_LC_15_26_4.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i12_LC_15_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i12_LC_15_26_4 (
            .in0(_gnd_net_),
            .in1(N__34843),
            .in2(_gnd_net_),
            .in3(N__34837),
            .lcout(n14),
            .ltout(),
            .carryin(n4448),
            .carryout(n4449),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i13_LC_15_26_5.C_ON=1'b1;
    defparam blink_counter_523__i13_LC_15_26_5.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i13_LC_15_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i13_LC_15_26_5 (
            .in0(_gnd_net_),
            .in1(N__34978),
            .in2(_gnd_net_),
            .in3(N__34972),
            .lcout(n13),
            .ltout(),
            .carryin(n4449),
            .carryout(n4450),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i14_LC_15_26_6.C_ON=1'b1;
    defparam blink_counter_523__i14_LC_15_26_6.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i14_LC_15_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i14_LC_15_26_6 (
            .in0(_gnd_net_),
            .in1(N__34969),
            .in2(_gnd_net_),
            .in3(N__34963),
            .lcout(n12),
            .ltout(),
            .carryin(n4450),
            .carryout(n4451),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i15_LC_15_26_7.C_ON=1'b1;
    defparam blink_counter_523__i15_LC_15_26_7.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i15_LC_15_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i15_LC_15_26_7 (
            .in0(_gnd_net_),
            .in1(N__34960),
            .in2(_gnd_net_),
            .in3(N__34954),
            .lcout(n11),
            .ltout(),
            .carryin(n4451),
            .carryout(n4452),
            .clk(N__35397),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i16_LC_15_27_0.C_ON=1'b1;
    defparam blink_counter_523__i16_LC_15_27_0.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i16_LC_15_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i16_LC_15_27_0 (
            .in0(_gnd_net_),
            .in1(N__34951),
            .in2(_gnd_net_),
            .in3(N__34945),
            .lcout(n10),
            .ltout(),
            .carryin(bfn_15_27_0_),
            .carryout(n4453),
            .clk(N__35404),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i17_LC_15_27_1.C_ON=1'b1;
    defparam blink_counter_523__i17_LC_15_27_1.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i17_LC_15_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i17_LC_15_27_1 (
            .in0(_gnd_net_),
            .in1(N__34942),
            .in2(_gnd_net_),
            .in3(N__34936),
            .lcout(n9),
            .ltout(),
            .carryin(n4453),
            .carryout(n4454),
            .clk(N__35404),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i18_LC_15_27_2.C_ON=1'b1;
    defparam blink_counter_523__i18_LC_15_27_2.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i18_LC_15_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i18_LC_15_27_2 (
            .in0(_gnd_net_),
            .in1(N__34933),
            .in2(_gnd_net_),
            .in3(N__34927),
            .lcout(n8_adj_1989),
            .ltout(),
            .carryin(n4454),
            .carryout(n4455),
            .clk(N__35404),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i19_LC_15_27_3.C_ON=1'b1;
    defparam blink_counter_523__i19_LC_15_27_3.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i19_LC_15_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i19_LC_15_27_3 (
            .in0(_gnd_net_),
            .in1(N__34924),
            .in2(_gnd_net_),
            .in3(N__34918),
            .lcout(n7),
            .ltout(),
            .carryin(n4455),
            .carryout(n4456),
            .clk(N__35404),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i20_LC_15_27_4.C_ON=1'b1;
    defparam blink_counter_523__i20_LC_15_27_4.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i20_LC_15_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i20_LC_15_27_4 (
            .in0(_gnd_net_),
            .in1(N__34915),
            .in2(_gnd_net_),
            .in3(N__34909),
            .lcout(n6),
            .ltout(),
            .carryin(n4456),
            .carryout(n4457),
            .clk(N__35404),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i21_LC_15_27_5.C_ON=1'b1;
    defparam blink_counter_523__i21_LC_15_27_5.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i21_LC_15_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i21_LC_15_27_5 (
            .in0(_gnd_net_),
            .in1(N__37452),
            .in2(_gnd_net_),
            .in3(N__37441),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n4457),
            .carryout(n4458),
            .clk(N__35404),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i22_LC_15_27_6.C_ON=1'b1;
    defparam blink_counter_523__i22_LC_15_27_6.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i22_LC_15_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i22_LC_15_27_6 (
            .in0(_gnd_net_),
            .in1(N__37428),
            .in2(_gnd_net_),
            .in3(N__37417),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n4458),
            .carryout(n4459),
            .clk(N__35404),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i23_LC_15_27_7.C_ON=1'b1;
    defparam blink_counter_523__i23_LC_15_27_7.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i23_LC_15_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i23_LC_15_27_7 (
            .in0(_gnd_net_),
            .in1(N__37401),
            .in2(_gnd_net_),
            .in3(N__37390),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n4459),
            .carryout(n4460),
            .clk(N__35404),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i24_LC_15_28_0.C_ON=1'b1;
    defparam blink_counter_523__i24_LC_15_28_0.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i24_LC_15_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i24_LC_15_28_0 (
            .in0(_gnd_net_),
            .in1(N__37374),
            .in2(_gnd_net_),
            .in3(N__37363),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_15_28_0_),
            .carryout(n4461),
            .clk(N__35408),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i25_LC_15_28_1.C_ON=1'b0;
    defparam blink_counter_523__i25_LC_15_28_1.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i25_LC_15_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i25_LC_15_28_1 (
            .in0(_gnd_net_),
            .in1(N__37350),
            .in2(_gnd_net_),
            .in3(N__37360),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35408),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i157_LC_16_27_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i157_LC_16_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i157_LC_16_27_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i157_LC_16_27_7  (
            .in0(N__35424),
            .in1(N__37339),
            .in2(N__37266),
            .in3(N__36292),
            .lcout(\c0.data_in_frame_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35409),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
