-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Sep 18 2019 23:28:45

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    PIN_9 : out std_logic;
    PIN_8 : in std_logic;
    PIN_7 : in std_logic;
    PIN_6 : inout std_logic;
    PIN_5 : inout std_logic;
    PIN_4 : inout std_logic;
    PIN_3 : out std_logic;
    PIN_24 : out std_logic;
    PIN_23 : out std_logic;
    PIN_22 : out std_logic;
    PIN_21 : in std_logic;
    PIN_20 : in std_logic;
    PIN_2 : out std_logic;
    PIN_19 : in std_logic;
    PIN_18 : in std_logic;
    PIN_17 : in std_logic;
    PIN_16 : in std_logic;
    PIN_15 : in std_logic;
    PIN_14 : in std_logic;
    PIN_13 : in std_logic;
    PIN_12 : in std_logic;
    PIN_11 : inout std_logic;
    PIN_10 : inout std_logic;
    PIN_1 : out std_logic;
    LED : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__70064\ : std_logic;
signal \N__70063\ : std_logic;
signal \N__70062\ : std_logic;
signal \N__70055\ : std_logic;
signal \N__70054\ : std_logic;
signal \N__70053\ : std_logic;
signal \N__70046\ : std_logic;
signal \N__70045\ : std_logic;
signal \N__70044\ : std_logic;
signal \N__70037\ : std_logic;
signal \N__70036\ : std_logic;
signal \N__70035\ : std_logic;
signal \N__70028\ : std_logic;
signal \N__70027\ : std_logic;
signal \N__70026\ : std_logic;
signal \N__70019\ : std_logic;
signal \N__70018\ : std_logic;
signal \N__70017\ : std_logic;
signal \N__70010\ : std_logic;
signal \N__70009\ : std_logic;
signal \N__70008\ : std_logic;
signal \N__70001\ : std_logic;
signal \N__70000\ : std_logic;
signal \N__69999\ : std_logic;
signal \N__69992\ : std_logic;
signal \N__69991\ : std_logic;
signal \N__69990\ : std_logic;
signal \N__69983\ : std_logic;
signal \N__69982\ : std_logic;
signal \N__69981\ : std_logic;
signal \N__69974\ : std_logic;
signal \N__69973\ : std_logic;
signal \N__69972\ : std_logic;
signal \N__69965\ : std_logic;
signal \N__69964\ : std_logic;
signal \N__69963\ : std_logic;
signal \N__69956\ : std_logic;
signal \N__69955\ : std_logic;
signal \N__69954\ : std_logic;
signal \N__69947\ : std_logic;
signal \N__69946\ : std_logic;
signal \N__69945\ : std_logic;
signal \N__69938\ : std_logic;
signal \N__69937\ : std_logic;
signal \N__69936\ : std_logic;
signal \N__69929\ : std_logic;
signal \N__69928\ : std_logic;
signal \N__69927\ : std_logic;
signal \N__69920\ : std_logic;
signal \N__69919\ : std_logic;
signal \N__69918\ : std_logic;
signal \N__69911\ : std_logic;
signal \N__69910\ : std_logic;
signal \N__69909\ : std_logic;
signal \N__69902\ : std_logic;
signal \N__69901\ : std_logic;
signal \N__69900\ : std_logic;
signal \N__69883\ : std_logic;
signal \N__69882\ : std_logic;
signal \N__69881\ : std_logic;
signal \N__69880\ : std_logic;
signal \N__69879\ : std_logic;
signal \N__69878\ : std_logic;
signal \N__69877\ : std_logic;
signal \N__69876\ : std_logic;
signal \N__69873\ : std_logic;
signal \N__69872\ : std_logic;
signal \N__69871\ : std_logic;
signal \N__69868\ : std_logic;
signal \N__69867\ : std_logic;
signal \N__69866\ : std_logic;
signal \N__69865\ : std_logic;
signal \N__69864\ : std_logic;
signal \N__69861\ : std_logic;
signal \N__69860\ : std_logic;
signal \N__69857\ : std_logic;
signal \N__69854\ : std_logic;
signal \N__69851\ : std_logic;
signal \N__69848\ : std_logic;
signal \N__69847\ : std_logic;
signal \N__69846\ : std_logic;
signal \N__69845\ : std_logic;
signal \N__69844\ : std_logic;
signal \N__69841\ : std_logic;
signal \N__69840\ : std_logic;
signal \N__69839\ : std_logic;
signal \N__69836\ : std_logic;
signal \N__69833\ : std_logic;
signal \N__69830\ : std_logic;
signal \N__69827\ : std_logic;
signal \N__69824\ : std_logic;
signal \N__69821\ : std_logic;
signal \N__69818\ : std_logic;
signal \N__69815\ : std_logic;
signal \N__69810\ : std_logic;
signal \N__69807\ : std_logic;
signal \N__69806\ : std_logic;
signal \N__69803\ : std_logic;
signal \N__69802\ : std_logic;
signal \N__69801\ : std_logic;
signal \N__69798\ : std_logic;
signal \N__69795\ : std_logic;
signal \N__69794\ : std_logic;
signal \N__69791\ : std_logic;
signal \N__69784\ : std_logic;
signal \N__69781\ : std_logic;
signal \N__69778\ : std_logic;
signal \N__69777\ : std_logic;
signal \N__69774\ : std_logic;
signal \N__69771\ : std_logic;
signal \N__69766\ : std_logic;
signal \N__69761\ : std_logic;
signal \N__69758\ : std_logic;
signal \N__69751\ : std_logic;
signal \N__69750\ : std_logic;
signal \N__69747\ : std_logic;
signal \N__69744\ : std_logic;
signal \N__69741\ : std_logic;
signal \N__69736\ : std_logic;
signal \N__69731\ : std_logic;
signal \N__69730\ : std_logic;
signal \N__69727\ : std_logic;
signal \N__69720\ : std_logic;
signal \N__69717\ : std_logic;
signal \N__69716\ : std_logic;
signal \N__69713\ : std_logic;
signal \N__69710\ : std_logic;
signal \N__69703\ : std_logic;
signal \N__69698\ : std_logic;
signal \N__69697\ : std_logic;
signal \N__69696\ : std_logic;
signal \N__69695\ : std_logic;
signal \N__69692\ : std_logic;
signal \N__69687\ : std_logic;
signal \N__69680\ : std_logic;
signal \N__69677\ : std_logic;
signal \N__69674\ : std_logic;
signal \N__69669\ : std_logic;
signal \N__69666\ : std_logic;
signal \N__69663\ : std_logic;
signal \N__69656\ : std_logic;
signal \N__69649\ : std_logic;
signal \N__69646\ : std_logic;
signal \N__69641\ : std_logic;
signal \N__69638\ : std_logic;
signal \N__69633\ : std_logic;
signal \N__69630\ : std_logic;
signal \N__69625\ : std_logic;
signal \N__69616\ : std_logic;
signal \N__69613\ : std_logic;
signal \N__69608\ : std_logic;
signal \N__69605\ : std_logic;
signal \N__69602\ : std_logic;
signal \N__69595\ : std_logic;
signal \N__69594\ : std_logic;
signal \N__69591\ : std_logic;
signal \N__69588\ : std_logic;
signal \N__69585\ : std_logic;
signal \N__69584\ : std_logic;
signal \N__69581\ : std_logic;
signal \N__69578\ : std_logic;
signal \N__69575\ : std_logic;
signal \N__69568\ : std_logic;
signal \N__69567\ : std_logic;
signal \N__69566\ : std_logic;
signal \N__69565\ : std_logic;
signal \N__69564\ : std_logic;
signal \N__69563\ : std_logic;
signal \N__69562\ : std_logic;
signal \N__69561\ : std_logic;
signal \N__69560\ : std_logic;
signal \N__69559\ : std_logic;
signal \N__69558\ : std_logic;
signal \N__69557\ : std_logic;
signal \N__69556\ : std_logic;
signal \N__69555\ : std_logic;
signal \N__69552\ : std_logic;
signal \N__69549\ : std_logic;
signal \N__69548\ : std_logic;
signal \N__69545\ : std_logic;
signal \N__69542\ : std_logic;
signal \N__69539\ : std_logic;
signal \N__69538\ : std_logic;
signal \N__69537\ : std_logic;
signal \N__69534\ : std_logic;
signal \N__69529\ : std_logic;
signal \N__69526\ : std_logic;
signal \N__69521\ : std_logic;
signal \N__69518\ : std_logic;
signal \N__69513\ : std_logic;
signal \N__69510\ : std_logic;
signal \N__69507\ : std_logic;
signal \N__69504\ : std_logic;
signal \N__69503\ : std_logic;
signal \N__69502\ : std_logic;
signal \N__69497\ : std_logic;
signal \N__69494\ : std_logic;
signal \N__69493\ : std_logic;
signal \N__69492\ : std_logic;
signal \N__69491\ : std_logic;
signal \N__69488\ : std_logic;
signal \N__69487\ : std_logic;
signal \N__69486\ : std_logic;
signal \N__69483\ : std_logic;
signal \N__69482\ : std_logic;
signal \N__69481\ : std_logic;
signal \N__69480\ : std_logic;
signal \N__69477\ : std_logic;
signal \N__69474\ : std_logic;
signal \N__69471\ : std_logic;
signal \N__69468\ : std_logic;
signal \N__69465\ : std_logic;
signal \N__69456\ : std_logic;
signal \N__69453\ : std_logic;
signal \N__69452\ : std_logic;
signal \N__69451\ : std_logic;
signal \N__69450\ : std_logic;
signal \N__69447\ : std_logic;
signal \N__69442\ : std_logic;
signal \N__69439\ : std_logic;
signal \N__69436\ : std_logic;
signal \N__69433\ : std_logic;
signal \N__69430\ : std_logic;
signal \N__69427\ : std_logic;
signal \N__69424\ : std_logic;
signal \N__69421\ : std_logic;
signal \N__69418\ : std_logic;
signal \N__69413\ : std_logic;
signal \N__69410\ : std_logic;
signal \N__69405\ : std_logic;
signal \N__69400\ : std_logic;
signal \N__69397\ : std_logic;
signal \N__69394\ : std_logic;
signal \N__69391\ : std_logic;
signal \N__69388\ : std_logic;
signal \N__69385\ : std_logic;
signal \N__69376\ : std_logic;
signal \N__69375\ : std_logic;
signal \N__69374\ : std_logic;
signal \N__69371\ : std_logic;
signal \N__69368\ : std_logic;
signal \N__69365\ : std_logic;
signal \N__69360\ : std_logic;
signal \N__69355\ : std_logic;
signal \N__69352\ : std_logic;
signal \N__69349\ : std_logic;
signal \N__69344\ : std_logic;
signal \N__69341\ : std_logic;
signal \N__69338\ : std_logic;
signal \N__69335\ : std_logic;
signal \N__69330\ : std_logic;
signal \N__69327\ : std_logic;
signal \N__69324\ : std_logic;
signal \N__69319\ : std_logic;
signal \N__69314\ : std_logic;
signal \N__69309\ : std_logic;
signal \N__69304\ : std_logic;
signal \N__69295\ : std_logic;
signal \N__69280\ : std_logic;
signal \N__69279\ : std_logic;
signal \N__69276\ : std_logic;
signal \N__69273\ : std_logic;
signal \N__69270\ : std_logic;
signal \N__69269\ : std_logic;
signal \N__69266\ : std_logic;
signal \N__69263\ : std_logic;
signal \N__69260\ : std_logic;
signal \N__69253\ : std_logic;
signal \N__69250\ : std_logic;
signal \N__69249\ : std_logic;
signal \N__69246\ : std_logic;
signal \N__69245\ : std_logic;
signal \N__69244\ : std_logic;
signal \N__69241\ : std_logic;
signal \N__69238\ : std_logic;
signal \N__69235\ : std_logic;
signal \N__69234\ : std_logic;
signal \N__69233\ : std_logic;
signal \N__69232\ : std_logic;
signal \N__69231\ : std_logic;
signal \N__69228\ : std_logic;
signal \N__69227\ : std_logic;
signal \N__69226\ : std_logic;
signal \N__69223\ : std_logic;
signal \N__69220\ : std_logic;
signal \N__69217\ : std_logic;
signal \N__69214\ : std_logic;
signal \N__69213\ : std_logic;
signal \N__69212\ : std_logic;
signal \N__69211\ : std_logic;
signal \N__69210\ : std_logic;
signal \N__69207\ : std_logic;
signal \N__69206\ : std_logic;
signal \N__69205\ : std_logic;
signal \N__69204\ : std_logic;
signal \N__69203\ : std_logic;
signal \N__69200\ : std_logic;
signal \N__69199\ : std_logic;
signal \N__69198\ : std_logic;
signal \N__69197\ : std_logic;
signal \N__69194\ : std_logic;
signal \N__69193\ : std_logic;
signal \N__69192\ : std_logic;
signal \N__69191\ : std_logic;
signal \N__69184\ : std_logic;
signal \N__69177\ : std_logic;
signal \N__69174\ : std_logic;
signal \N__69169\ : std_logic;
signal \N__69168\ : std_logic;
signal \N__69165\ : std_logic;
signal \N__69162\ : std_logic;
signal \N__69155\ : std_logic;
signal \N__69152\ : std_logic;
signal \N__69151\ : std_logic;
signal \N__69148\ : std_logic;
signal \N__69143\ : std_logic;
signal \N__69138\ : std_logic;
signal \N__69135\ : std_logic;
signal \N__69132\ : std_logic;
signal \N__69129\ : std_logic;
signal \N__69126\ : std_logic;
signal \N__69125\ : std_logic;
signal \N__69124\ : std_logic;
signal \N__69119\ : std_logic;
signal \N__69116\ : std_logic;
signal \N__69113\ : std_logic;
signal \N__69110\ : std_logic;
signal \N__69107\ : std_logic;
signal \N__69100\ : std_logic;
signal \N__69097\ : std_logic;
signal \N__69094\ : std_logic;
signal \N__69089\ : std_logic;
signal \N__69086\ : std_logic;
signal \N__69081\ : std_logic;
signal \N__69078\ : std_logic;
signal \N__69075\ : std_logic;
signal \N__69072\ : std_logic;
signal \N__69069\ : std_logic;
signal \N__69066\ : std_logic;
signal \N__69065\ : std_logic;
signal \N__69064\ : std_logic;
signal \N__69063\ : std_logic;
signal \N__69062\ : std_logic;
signal \N__69059\ : std_logic;
signal \N__69056\ : std_logic;
signal \N__69053\ : std_logic;
signal \N__69050\ : std_logic;
signal \N__69043\ : std_logic;
signal \N__69034\ : std_logic;
signal \N__69027\ : std_logic;
signal \N__69018\ : std_logic;
signal \N__69015\ : std_logic;
signal \N__69008\ : std_logic;
signal \N__69005\ : std_logic;
signal \N__69000\ : std_logic;
signal \N__68989\ : std_logic;
signal \N__68988\ : std_logic;
signal \N__68987\ : std_logic;
signal \N__68984\ : std_logic;
signal \N__68981\ : std_logic;
signal \N__68980\ : std_logic;
signal \N__68979\ : std_logic;
signal \N__68976\ : std_logic;
signal \N__68975\ : std_logic;
signal \N__68974\ : std_logic;
signal \N__68973\ : std_logic;
signal \N__68972\ : std_logic;
signal \N__68971\ : std_logic;
signal \N__68970\ : std_logic;
signal \N__68965\ : std_logic;
signal \N__68962\ : std_logic;
signal \N__68959\ : std_logic;
signal \N__68958\ : std_logic;
signal \N__68957\ : std_logic;
signal \N__68956\ : std_logic;
signal \N__68955\ : std_logic;
signal \N__68954\ : std_logic;
signal \N__68951\ : std_logic;
signal \N__68948\ : std_logic;
signal \N__68945\ : std_logic;
signal \N__68944\ : std_logic;
signal \N__68941\ : std_logic;
signal \N__68940\ : std_logic;
signal \N__68939\ : std_logic;
signal \N__68938\ : std_logic;
signal \N__68935\ : std_logic;
signal \N__68932\ : std_logic;
signal \N__68929\ : std_logic;
signal \N__68926\ : std_logic;
signal \N__68921\ : std_logic;
signal \N__68916\ : std_logic;
signal \N__68913\ : std_logic;
signal \N__68910\ : std_logic;
signal \N__68909\ : std_logic;
signal \N__68908\ : std_logic;
signal \N__68905\ : std_logic;
signal \N__68900\ : std_logic;
signal \N__68897\ : std_logic;
signal \N__68894\ : std_logic;
signal \N__68889\ : std_logic;
signal \N__68884\ : std_logic;
signal \N__68883\ : std_logic;
signal \N__68882\ : std_logic;
signal \N__68881\ : std_logic;
signal \N__68880\ : std_logic;
signal \N__68877\ : std_logic;
signal \N__68876\ : std_logic;
signal \N__68873\ : std_logic;
signal \N__68868\ : std_logic;
signal \N__68867\ : std_logic;
signal \N__68866\ : std_logic;
signal \N__68865\ : std_logic;
signal \N__68862\ : std_logic;
signal \N__68855\ : std_logic;
signal \N__68852\ : std_logic;
signal \N__68849\ : std_logic;
signal \N__68846\ : std_logic;
signal \N__68837\ : std_logic;
signal \N__68834\ : std_logic;
signal \N__68831\ : std_logic;
signal \N__68826\ : std_logic;
signal \N__68823\ : std_logic;
signal \N__68820\ : std_logic;
signal \N__68817\ : std_logic;
signal \N__68812\ : std_logic;
signal \N__68809\ : std_logic;
signal \N__68806\ : std_logic;
signal \N__68803\ : std_logic;
signal \N__68800\ : std_logic;
signal \N__68797\ : std_logic;
signal \N__68792\ : std_logic;
signal \N__68789\ : std_logic;
signal \N__68786\ : std_logic;
signal \N__68785\ : std_logic;
signal \N__68784\ : std_logic;
signal \N__68781\ : std_logic;
signal \N__68776\ : std_logic;
signal \N__68771\ : std_logic;
signal \N__68766\ : std_logic;
signal \N__68763\ : std_logic;
signal \N__68756\ : std_logic;
signal \N__68753\ : std_logic;
signal \N__68746\ : std_logic;
signal \N__68743\ : std_logic;
signal \N__68740\ : std_logic;
signal \N__68731\ : std_logic;
signal \N__68722\ : std_logic;
signal \N__68713\ : std_logic;
signal \N__68712\ : std_logic;
signal \N__68709\ : std_logic;
signal \N__68706\ : std_logic;
signal \N__68705\ : std_logic;
signal \N__68702\ : std_logic;
signal \N__68699\ : std_logic;
signal \N__68696\ : std_logic;
signal \N__68695\ : std_logic;
signal \N__68690\ : std_logic;
signal \N__68685\ : std_logic;
signal \N__68680\ : std_logic;
signal \N__68679\ : std_logic;
signal \N__68678\ : std_logic;
signal \N__68675\ : std_logic;
signal \N__68674\ : std_logic;
signal \N__68673\ : std_logic;
signal \N__68672\ : std_logic;
signal \N__68671\ : std_logic;
signal \N__68670\ : std_logic;
signal \N__68669\ : std_logic;
signal \N__68666\ : std_logic;
signal \N__68663\ : std_logic;
signal \N__68660\ : std_logic;
signal \N__68659\ : std_logic;
signal \N__68658\ : std_logic;
signal \N__68655\ : std_logic;
signal \N__68650\ : std_logic;
signal \N__68647\ : std_logic;
signal \N__68644\ : std_logic;
signal \N__68639\ : std_logic;
signal \N__68638\ : std_logic;
signal \N__68633\ : std_logic;
signal \N__68632\ : std_logic;
signal \N__68629\ : std_logic;
signal \N__68628\ : std_logic;
signal \N__68625\ : std_logic;
signal \N__68620\ : std_logic;
signal \N__68617\ : std_logic;
signal \N__68614\ : std_logic;
signal \N__68611\ : std_logic;
signal \N__68608\ : std_logic;
signal \N__68605\ : std_logic;
signal \N__68602\ : std_logic;
signal \N__68601\ : std_logic;
signal \N__68600\ : std_logic;
signal \N__68595\ : std_logic;
signal \N__68592\ : std_logic;
signal \N__68591\ : std_logic;
signal \N__68590\ : std_logic;
signal \N__68589\ : std_logic;
signal \N__68584\ : std_logic;
signal \N__68579\ : std_logic;
signal \N__68576\ : std_logic;
signal \N__68571\ : std_logic;
signal \N__68570\ : std_logic;
signal \N__68569\ : std_logic;
signal \N__68568\ : std_logic;
signal \N__68565\ : std_logic;
signal \N__68562\ : std_logic;
signal \N__68557\ : std_logic;
signal \N__68554\ : std_logic;
signal \N__68553\ : std_logic;
signal \N__68552\ : std_logic;
signal \N__68549\ : std_logic;
signal \N__68546\ : std_logic;
signal \N__68545\ : std_logic;
signal \N__68542\ : std_logic;
signal \N__68539\ : std_logic;
signal \N__68536\ : std_logic;
signal \N__68533\ : std_logic;
signal \N__68530\ : std_logic;
signal \N__68527\ : std_logic;
signal \N__68524\ : std_logic;
signal \N__68517\ : std_logic;
signal \N__68516\ : std_logic;
signal \N__68513\ : std_logic;
signal \N__68506\ : std_logic;
signal \N__68503\ : std_logic;
signal \N__68500\ : std_logic;
signal \N__68493\ : std_logic;
signal \N__68488\ : std_logic;
signal \N__68485\ : std_logic;
signal \N__68480\ : std_logic;
signal \N__68477\ : std_logic;
signal \N__68468\ : std_logic;
signal \N__68463\ : std_logic;
signal \N__68460\ : std_logic;
signal \N__68457\ : std_logic;
signal \N__68450\ : std_logic;
signal \N__68443\ : std_logic;
signal \N__68442\ : std_logic;
signal \N__68441\ : std_logic;
signal \N__68438\ : std_logic;
signal \N__68437\ : std_logic;
signal \N__68436\ : std_logic;
signal \N__68435\ : std_logic;
signal \N__68434\ : std_logic;
signal \N__68433\ : std_logic;
signal \N__68430\ : std_logic;
signal \N__68427\ : std_logic;
signal \N__68426\ : std_logic;
signal \N__68423\ : std_logic;
signal \N__68420\ : std_logic;
signal \N__68419\ : std_logic;
signal \N__68418\ : std_logic;
signal \N__68417\ : std_logic;
signal \N__68416\ : std_logic;
signal \N__68413\ : std_logic;
signal \N__68412\ : std_logic;
signal \N__68411\ : std_logic;
signal \N__68410\ : std_logic;
signal \N__68407\ : std_logic;
signal \N__68404\ : std_logic;
signal \N__68399\ : std_logic;
signal \N__68396\ : std_logic;
signal \N__68395\ : std_logic;
signal \N__68394\ : std_logic;
signal \N__68393\ : std_logic;
signal \N__68390\ : std_logic;
signal \N__68385\ : std_logic;
signal \N__68378\ : std_logic;
signal \N__68377\ : std_logic;
signal \N__68374\ : std_logic;
signal \N__68373\ : std_logic;
signal \N__68370\ : std_logic;
signal \N__68369\ : std_logic;
signal \N__68366\ : std_logic;
signal \N__68363\ : std_logic;
signal \N__68360\ : std_logic;
signal \N__68359\ : std_logic;
signal \N__68358\ : std_logic;
signal \N__68357\ : std_logic;
signal \N__68356\ : std_logic;
signal \N__68355\ : std_logic;
signal \N__68354\ : std_logic;
signal \N__68353\ : std_logic;
signal \N__68352\ : std_logic;
signal \N__68349\ : std_logic;
signal \N__68346\ : std_logic;
signal \N__68341\ : std_logic;
signal \N__68338\ : std_logic;
signal \N__68333\ : std_logic;
signal \N__68330\ : std_logic;
signal \N__68325\ : std_logic;
signal \N__68322\ : std_logic;
signal \N__68319\ : std_logic;
signal \N__68316\ : std_logic;
signal \N__68313\ : std_logic;
signal \N__68310\ : std_logic;
signal \N__68307\ : std_logic;
signal \N__68304\ : std_logic;
signal \N__68301\ : std_logic;
signal \N__68296\ : std_logic;
signal \N__68293\ : std_logic;
signal \N__68290\ : std_logic;
signal \N__68289\ : std_logic;
signal \N__68288\ : std_logic;
signal \N__68285\ : std_logic;
signal \N__68280\ : std_logic;
signal \N__68277\ : std_logic;
signal \N__68274\ : std_logic;
signal \N__68269\ : std_logic;
signal \N__68262\ : std_logic;
signal \N__68259\ : std_logic;
signal \N__68256\ : std_logic;
signal \N__68251\ : std_logic;
signal \N__68248\ : std_logic;
signal \N__68243\ : std_logic;
signal \N__68238\ : std_logic;
signal \N__68235\ : std_logic;
signal \N__68230\ : std_logic;
signal \N__68227\ : std_logic;
signal \N__68224\ : std_logic;
signal \N__68219\ : std_logic;
signal \N__68216\ : std_logic;
signal \N__68211\ : std_logic;
signal \N__68208\ : std_logic;
signal \N__68205\ : std_logic;
signal \N__68196\ : std_logic;
signal \N__68189\ : std_logic;
signal \N__68178\ : std_logic;
signal \N__68167\ : std_logic;
signal \N__68166\ : std_logic;
signal \N__68165\ : std_logic;
signal \N__68164\ : std_logic;
signal \N__68163\ : std_logic;
signal \N__68162\ : std_logic;
signal \N__68161\ : std_logic;
signal \N__68160\ : std_logic;
signal \N__68159\ : std_logic;
signal \N__68158\ : std_logic;
signal \N__68157\ : std_logic;
signal \N__68156\ : std_logic;
signal \N__68155\ : std_logic;
signal \N__68152\ : std_logic;
signal \N__68149\ : std_logic;
signal \N__68148\ : std_logic;
signal \N__68147\ : std_logic;
signal \N__68146\ : std_logic;
signal \N__68145\ : std_logic;
signal \N__68144\ : std_logic;
signal \N__68143\ : std_logic;
signal \N__68142\ : std_logic;
signal \N__68141\ : std_logic;
signal \N__68140\ : std_logic;
signal \N__68139\ : std_logic;
signal \N__68138\ : std_logic;
signal \N__68137\ : std_logic;
signal \N__68136\ : std_logic;
signal \N__68135\ : std_logic;
signal \N__68132\ : std_logic;
signal \N__68129\ : std_logic;
signal \N__68122\ : std_logic;
signal \N__68117\ : std_logic;
signal \N__68112\ : std_logic;
signal \N__68111\ : std_logic;
signal \N__68110\ : std_logic;
signal \N__68109\ : std_logic;
signal \N__68104\ : std_logic;
signal \N__68101\ : std_logic;
signal \N__68098\ : std_logic;
signal \N__68097\ : std_logic;
signal \N__68096\ : std_logic;
signal \N__68095\ : std_logic;
signal \N__68094\ : std_logic;
signal \N__68093\ : std_logic;
signal \N__68092\ : std_logic;
signal \N__68091\ : std_logic;
signal \N__68088\ : std_logic;
signal \N__68087\ : std_logic;
signal \N__68086\ : std_logic;
signal \N__68083\ : std_logic;
signal \N__68078\ : std_logic;
signal \N__68071\ : std_logic;
signal \N__68070\ : std_logic;
signal \N__68069\ : std_logic;
signal \N__68068\ : std_logic;
signal \N__68067\ : std_logic;
signal \N__68066\ : std_logic;
signal \N__68065\ : std_logic;
signal \N__68062\ : std_logic;
signal \N__68057\ : std_logic;
signal \N__68048\ : std_logic;
signal \N__68045\ : std_logic;
signal \N__68044\ : std_logic;
signal \N__68043\ : std_logic;
signal \N__68042\ : std_logic;
signal \N__68039\ : std_logic;
signal \N__68036\ : std_logic;
signal \N__68033\ : std_logic;
signal \N__68030\ : std_logic;
signal \N__68023\ : std_logic;
signal \N__68020\ : std_logic;
signal \N__68019\ : std_logic;
signal \N__68018\ : std_logic;
signal \N__68017\ : std_logic;
signal \N__68012\ : std_logic;
signal \N__68009\ : std_logic;
signal \N__68008\ : std_logic;
signal \N__68007\ : std_logic;
signal \N__68006\ : std_logic;
signal \N__68003\ : std_logic;
signal \N__68000\ : std_logic;
signal \N__67995\ : std_logic;
signal \N__67990\ : std_logic;
signal \N__67987\ : std_logic;
signal \N__67984\ : std_logic;
signal \N__67979\ : std_logic;
signal \N__67974\ : std_logic;
signal \N__67971\ : std_logic;
signal \N__67966\ : std_logic;
signal \N__67959\ : std_logic;
signal \N__67954\ : std_logic;
signal \N__67949\ : std_logic;
signal \N__67946\ : std_logic;
signal \N__67941\ : std_logic;
signal \N__67938\ : std_logic;
signal \N__67933\ : std_logic;
signal \N__67926\ : std_logic;
signal \N__67919\ : std_logic;
signal \N__67916\ : std_logic;
signal \N__67913\ : std_logic;
signal \N__67912\ : std_logic;
signal \N__67911\ : std_logic;
signal \N__67904\ : std_logic;
signal \N__67901\ : std_logic;
signal \N__67892\ : std_logic;
signal \N__67885\ : std_logic;
signal \N__67874\ : std_logic;
signal \N__67871\ : std_logic;
signal \N__67866\ : std_logic;
signal \N__67861\ : std_logic;
signal \N__67854\ : std_logic;
signal \N__67849\ : std_logic;
signal \N__67838\ : std_logic;
signal \N__67831\ : std_logic;
signal \N__67828\ : std_logic;
signal \N__67819\ : std_logic;
signal \N__67818\ : std_logic;
signal \N__67815\ : std_logic;
signal \N__67812\ : std_logic;
signal \N__67811\ : std_logic;
signal \N__67808\ : std_logic;
signal \N__67805\ : std_logic;
signal \N__67802\ : std_logic;
signal \N__67795\ : std_logic;
signal \N__67794\ : std_logic;
signal \N__67793\ : std_logic;
signal \N__67792\ : std_logic;
signal \N__67791\ : std_logic;
signal \N__67784\ : std_logic;
signal \N__67779\ : std_logic;
signal \N__67778\ : std_logic;
signal \N__67777\ : std_logic;
signal \N__67776\ : std_logic;
signal \N__67775\ : std_logic;
signal \N__67770\ : std_logic;
signal \N__67765\ : std_logic;
signal \N__67764\ : std_logic;
signal \N__67763\ : std_logic;
signal \N__67762\ : std_logic;
signal \N__67761\ : std_logic;
signal \N__67760\ : std_logic;
signal \N__67759\ : std_logic;
signal \N__67758\ : std_logic;
signal \N__67757\ : std_logic;
signal \N__67756\ : std_logic;
signal \N__67753\ : std_logic;
signal \N__67752\ : std_logic;
signal \N__67751\ : std_logic;
signal \N__67750\ : std_logic;
signal \N__67749\ : std_logic;
signal \N__67748\ : std_logic;
signal \N__67745\ : std_logic;
signal \N__67744\ : std_logic;
signal \N__67739\ : std_logic;
signal \N__67734\ : std_logic;
signal \N__67733\ : std_logic;
signal \N__67732\ : std_logic;
signal \N__67731\ : std_logic;
signal \N__67724\ : std_logic;
signal \N__67721\ : std_logic;
signal \N__67718\ : std_logic;
signal \N__67715\ : std_logic;
signal \N__67712\ : std_logic;
signal \N__67709\ : std_logic;
signal \N__67708\ : std_logic;
signal \N__67707\ : std_logic;
signal \N__67706\ : std_logic;
signal \N__67705\ : std_logic;
signal \N__67702\ : std_logic;
signal \N__67699\ : std_logic;
signal \N__67692\ : std_logic;
signal \N__67689\ : std_logic;
signal \N__67686\ : std_logic;
signal \N__67685\ : std_logic;
signal \N__67682\ : std_logic;
signal \N__67679\ : std_logic;
signal \N__67678\ : std_logic;
signal \N__67677\ : std_logic;
signal \N__67676\ : std_logic;
signal \N__67675\ : std_logic;
signal \N__67674\ : std_logic;
signal \N__67673\ : std_logic;
signal \N__67672\ : std_logic;
signal \N__67665\ : std_logic;
signal \N__67662\ : std_logic;
signal \N__67659\ : std_logic;
signal \N__67656\ : std_logic;
signal \N__67649\ : std_logic;
signal \N__67646\ : std_logic;
signal \N__67643\ : std_logic;
signal \N__67638\ : std_logic;
signal \N__67633\ : std_logic;
signal \N__67630\ : std_logic;
signal \N__67625\ : std_logic;
signal \N__67624\ : std_logic;
signal \N__67623\ : std_logic;
signal \N__67622\ : std_logic;
signal \N__67621\ : std_logic;
signal \N__67620\ : std_logic;
signal \N__67617\ : std_logic;
signal \N__67612\ : std_logic;
signal \N__67611\ : std_logic;
signal \N__67610\ : std_logic;
signal \N__67609\ : std_logic;
signal \N__67606\ : std_logic;
signal \N__67603\ : std_logic;
signal \N__67600\ : std_logic;
signal \N__67597\ : std_logic;
signal \N__67592\ : std_logic;
signal \N__67589\ : std_logic;
signal \N__67586\ : std_logic;
signal \N__67583\ : std_logic;
signal \N__67576\ : std_logic;
signal \N__67573\ : std_logic;
signal \N__67564\ : std_logic;
signal \N__67561\ : std_logic;
signal \N__67556\ : std_logic;
signal \N__67553\ : std_logic;
signal \N__67548\ : std_logic;
signal \N__67545\ : std_logic;
signal \N__67542\ : std_logic;
signal \N__67539\ : std_logic;
signal \N__67536\ : std_logic;
signal \N__67533\ : std_logic;
signal \N__67522\ : std_logic;
signal \N__67513\ : std_logic;
signal \N__67506\ : std_logic;
signal \N__67495\ : std_logic;
signal \N__67480\ : std_logic;
signal \N__67479\ : std_logic;
signal \N__67478\ : std_logic;
signal \N__67477\ : std_logic;
signal \N__67476\ : std_logic;
signal \N__67475\ : std_logic;
signal \N__67472\ : std_logic;
signal \N__67471\ : std_logic;
signal \N__67470\ : std_logic;
signal \N__67469\ : std_logic;
signal \N__67466\ : std_logic;
signal \N__67463\ : std_logic;
signal \N__67462\ : std_logic;
signal \N__67461\ : std_logic;
signal \N__67460\ : std_logic;
signal \N__67459\ : std_logic;
signal \N__67458\ : std_logic;
signal \N__67457\ : std_logic;
signal \N__67454\ : std_logic;
signal \N__67453\ : std_logic;
signal \N__67452\ : std_logic;
signal \N__67451\ : std_logic;
signal \N__67446\ : std_logic;
signal \N__67445\ : std_logic;
signal \N__67440\ : std_logic;
signal \N__67437\ : std_logic;
signal \N__67434\ : std_logic;
signal \N__67425\ : std_logic;
signal \N__67418\ : std_logic;
signal \N__67415\ : std_logic;
signal \N__67412\ : std_logic;
signal \N__67409\ : std_logic;
signal \N__67408\ : std_logic;
signal \N__67407\ : std_logic;
signal \N__67404\ : std_logic;
signal \N__67403\ : std_logic;
signal \N__67402\ : std_logic;
signal \N__67399\ : std_logic;
signal \N__67396\ : std_logic;
signal \N__67393\ : std_logic;
signal \N__67392\ : std_logic;
signal \N__67391\ : std_logic;
signal \N__67386\ : std_logic;
signal \N__67383\ : std_logic;
signal \N__67380\ : std_logic;
signal \N__67379\ : std_logic;
signal \N__67376\ : std_logic;
signal \N__67373\ : std_logic;
signal \N__67368\ : std_logic;
signal \N__67365\ : std_logic;
signal \N__67364\ : std_logic;
signal \N__67363\ : std_logic;
signal \N__67362\ : std_logic;
signal \N__67361\ : std_logic;
signal \N__67358\ : std_logic;
signal \N__67355\ : std_logic;
signal \N__67352\ : std_logic;
signal \N__67349\ : std_logic;
signal \N__67348\ : std_logic;
signal \N__67345\ : std_logic;
signal \N__67340\ : std_logic;
signal \N__67339\ : std_logic;
signal \N__67334\ : std_logic;
signal \N__67331\ : std_logic;
signal \N__67326\ : std_logic;
signal \N__67323\ : std_logic;
signal \N__67320\ : std_logic;
signal \N__67317\ : std_logic;
signal \N__67312\ : std_logic;
signal \N__67307\ : std_logic;
signal \N__67304\ : std_logic;
signal \N__67301\ : std_logic;
signal \N__67296\ : std_logic;
signal \N__67293\ : std_logic;
signal \N__67290\ : std_logic;
signal \N__67287\ : std_logic;
signal \N__67282\ : std_logic;
signal \N__67279\ : std_logic;
signal \N__67272\ : std_logic;
signal \N__67269\ : std_logic;
signal \N__67262\ : std_logic;
signal \N__67251\ : std_logic;
signal \N__67240\ : std_logic;
signal \N__67237\ : std_logic;
signal \N__67234\ : std_logic;
signal \N__67231\ : std_logic;
signal \N__67228\ : std_logic;
signal \N__67219\ : std_logic;
signal \N__67218\ : std_logic;
signal \N__67217\ : std_logic;
signal \N__67216\ : std_logic;
signal \N__67215\ : std_logic;
signal \N__67214\ : std_logic;
signal \N__67211\ : std_logic;
signal \N__67210\ : std_logic;
signal \N__67209\ : std_logic;
signal \N__67208\ : std_logic;
signal \N__67207\ : std_logic;
signal \N__67206\ : std_logic;
signal \N__67203\ : std_logic;
signal \N__67202\ : std_logic;
signal \N__67201\ : std_logic;
signal \N__67196\ : std_logic;
signal \N__67193\ : std_logic;
signal \N__67190\ : std_logic;
signal \N__67187\ : std_logic;
signal \N__67186\ : std_logic;
signal \N__67183\ : std_logic;
signal \N__67180\ : std_logic;
signal \N__67177\ : std_logic;
signal \N__67172\ : std_logic;
signal \N__67171\ : std_logic;
signal \N__67170\ : std_logic;
signal \N__67167\ : std_logic;
signal \N__67164\ : std_logic;
signal \N__67163\ : std_logic;
signal \N__67162\ : std_logic;
signal \N__67161\ : std_logic;
signal \N__67158\ : std_logic;
signal \N__67157\ : std_logic;
signal \N__67154\ : std_logic;
signal \N__67149\ : std_logic;
signal \N__67146\ : std_logic;
signal \N__67143\ : std_logic;
signal \N__67142\ : std_logic;
signal \N__67139\ : std_logic;
signal \N__67134\ : std_logic;
signal \N__67131\ : std_logic;
signal \N__67128\ : std_logic;
signal \N__67125\ : std_logic;
signal \N__67124\ : std_logic;
signal \N__67123\ : std_logic;
signal \N__67122\ : std_logic;
signal \N__67117\ : std_logic;
signal \N__67114\ : std_logic;
signal \N__67111\ : std_logic;
signal \N__67108\ : std_logic;
signal \N__67105\ : std_logic;
signal \N__67104\ : std_logic;
signal \N__67103\ : std_logic;
signal \N__67100\ : std_logic;
signal \N__67097\ : std_logic;
signal \N__67094\ : std_logic;
signal \N__67089\ : std_logic;
signal \N__67086\ : std_logic;
signal \N__67083\ : std_logic;
signal \N__67080\ : std_logic;
signal \N__67079\ : std_logic;
signal \N__67076\ : std_logic;
signal \N__67071\ : std_logic;
signal \N__67070\ : std_logic;
signal \N__67067\ : std_logic;
signal \N__67064\ : std_logic;
signal \N__67063\ : std_logic;
signal \N__67060\ : std_logic;
signal \N__67057\ : std_logic;
signal \N__67054\ : std_logic;
signal \N__67051\ : std_logic;
signal \N__67046\ : std_logic;
signal \N__67043\ : std_logic;
signal \N__67040\ : std_logic;
signal \N__67033\ : std_logic;
signal \N__67030\ : std_logic;
signal \N__67027\ : std_logic;
signal \N__67022\ : std_logic;
signal \N__67019\ : std_logic;
signal \N__67014\ : std_logic;
signal \N__67011\ : std_logic;
signal \N__67006\ : std_logic;
signal \N__67005\ : std_logic;
signal \N__67002\ : std_logic;
signal \N__66991\ : std_logic;
signal \N__66982\ : std_logic;
signal \N__66979\ : std_logic;
signal \N__66976\ : std_logic;
signal \N__66975\ : std_logic;
signal \N__66974\ : std_logic;
signal \N__66971\ : std_logic;
signal \N__66968\ : std_logic;
signal \N__66963\ : std_logic;
signal \N__66960\ : std_logic;
signal \N__66953\ : std_logic;
signal \N__66948\ : std_logic;
signal \N__66945\ : std_logic;
signal \N__66942\ : std_logic;
signal \N__66939\ : std_logic;
signal \N__66934\ : std_logic;
signal \N__66929\ : std_logic;
signal \N__66926\ : std_logic;
signal \N__66913\ : std_logic;
signal \N__66912\ : std_logic;
signal \N__66909\ : std_logic;
signal \N__66908\ : std_logic;
signal \N__66905\ : std_logic;
signal \N__66902\ : std_logic;
signal \N__66899\ : std_logic;
signal \N__66896\ : std_logic;
signal \N__66893\ : std_logic;
signal \N__66890\ : std_logic;
signal \N__66883\ : std_logic;
signal \N__66880\ : std_logic;
signal \N__66877\ : std_logic;
signal \N__66876\ : std_logic;
signal \N__66875\ : std_logic;
signal \N__66872\ : std_logic;
signal \N__66871\ : std_logic;
signal \N__66870\ : std_logic;
signal \N__66869\ : std_logic;
signal \N__66868\ : std_logic;
signal \N__66867\ : std_logic;
signal \N__66866\ : std_logic;
signal \N__66865\ : std_logic;
signal \N__66864\ : std_logic;
signal \N__66863\ : std_logic;
signal \N__66862\ : std_logic;
signal \N__66861\ : std_logic;
signal \N__66860\ : std_logic;
signal \N__66859\ : std_logic;
signal \N__66858\ : std_logic;
signal \N__66857\ : std_logic;
signal \N__66856\ : std_logic;
signal \N__66855\ : std_logic;
signal \N__66854\ : std_logic;
signal \N__66853\ : std_logic;
signal \N__66852\ : std_logic;
signal \N__66851\ : std_logic;
signal \N__66850\ : std_logic;
signal \N__66849\ : std_logic;
signal \N__66848\ : std_logic;
signal \N__66847\ : std_logic;
signal \N__66846\ : std_logic;
signal \N__66845\ : std_logic;
signal \N__66844\ : std_logic;
signal \N__66843\ : std_logic;
signal \N__66842\ : std_logic;
signal \N__66841\ : std_logic;
signal \N__66840\ : std_logic;
signal \N__66839\ : std_logic;
signal \N__66838\ : std_logic;
signal \N__66837\ : std_logic;
signal \N__66836\ : std_logic;
signal \N__66835\ : std_logic;
signal \N__66834\ : std_logic;
signal \N__66833\ : std_logic;
signal \N__66832\ : std_logic;
signal \N__66831\ : std_logic;
signal \N__66830\ : std_logic;
signal \N__66829\ : std_logic;
signal \N__66828\ : std_logic;
signal \N__66827\ : std_logic;
signal \N__66826\ : std_logic;
signal \N__66825\ : std_logic;
signal \N__66824\ : std_logic;
signal \N__66823\ : std_logic;
signal \N__66822\ : std_logic;
signal \N__66821\ : std_logic;
signal \N__66820\ : std_logic;
signal \N__66819\ : std_logic;
signal \N__66818\ : std_logic;
signal \N__66817\ : std_logic;
signal \N__66816\ : std_logic;
signal \N__66815\ : std_logic;
signal \N__66814\ : std_logic;
signal \N__66813\ : std_logic;
signal \N__66812\ : std_logic;
signal \N__66811\ : std_logic;
signal \N__66810\ : std_logic;
signal \N__66809\ : std_logic;
signal \N__66808\ : std_logic;
signal \N__66807\ : std_logic;
signal \N__66806\ : std_logic;
signal \N__66805\ : std_logic;
signal \N__66804\ : std_logic;
signal \N__66803\ : std_logic;
signal \N__66802\ : std_logic;
signal \N__66801\ : std_logic;
signal \N__66800\ : std_logic;
signal \N__66799\ : std_logic;
signal \N__66798\ : std_logic;
signal \N__66797\ : std_logic;
signal \N__66796\ : std_logic;
signal \N__66795\ : std_logic;
signal \N__66794\ : std_logic;
signal \N__66793\ : std_logic;
signal \N__66792\ : std_logic;
signal \N__66791\ : std_logic;
signal \N__66790\ : std_logic;
signal \N__66789\ : std_logic;
signal \N__66788\ : std_logic;
signal \N__66787\ : std_logic;
signal \N__66786\ : std_logic;
signal \N__66785\ : std_logic;
signal \N__66784\ : std_logic;
signal \N__66783\ : std_logic;
signal \N__66782\ : std_logic;
signal \N__66781\ : std_logic;
signal \N__66780\ : std_logic;
signal \N__66779\ : std_logic;
signal \N__66778\ : std_logic;
signal \N__66777\ : std_logic;
signal \N__66776\ : std_logic;
signal \N__66775\ : std_logic;
signal \N__66774\ : std_logic;
signal \N__66773\ : std_logic;
signal \N__66772\ : std_logic;
signal \N__66771\ : std_logic;
signal \N__66770\ : std_logic;
signal \N__66769\ : std_logic;
signal \N__66768\ : std_logic;
signal \N__66767\ : std_logic;
signal \N__66766\ : std_logic;
signal \N__66765\ : std_logic;
signal \N__66764\ : std_logic;
signal \N__66763\ : std_logic;
signal \N__66762\ : std_logic;
signal \N__66761\ : std_logic;
signal \N__66760\ : std_logic;
signal \N__66759\ : std_logic;
signal \N__66758\ : std_logic;
signal \N__66757\ : std_logic;
signal \N__66756\ : std_logic;
signal \N__66755\ : std_logic;
signal \N__66754\ : std_logic;
signal \N__66753\ : std_logic;
signal \N__66752\ : std_logic;
signal \N__66751\ : std_logic;
signal \N__66750\ : std_logic;
signal \N__66749\ : std_logic;
signal \N__66748\ : std_logic;
signal \N__66747\ : std_logic;
signal \N__66746\ : std_logic;
signal \N__66745\ : std_logic;
signal \N__66744\ : std_logic;
signal \N__66743\ : std_logic;
signal \N__66742\ : std_logic;
signal \N__66741\ : std_logic;
signal \N__66740\ : std_logic;
signal \N__66739\ : std_logic;
signal \N__66738\ : std_logic;
signal \N__66737\ : std_logic;
signal \N__66736\ : std_logic;
signal \N__66735\ : std_logic;
signal \N__66734\ : std_logic;
signal \N__66733\ : std_logic;
signal \N__66732\ : std_logic;
signal \N__66731\ : std_logic;
signal \N__66730\ : std_logic;
signal \N__66729\ : std_logic;
signal \N__66728\ : std_logic;
signal \N__66727\ : std_logic;
signal \N__66726\ : std_logic;
signal \N__66725\ : std_logic;
signal \N__66724\ : std_logic;
signal \N__66723\ : std_logic;
signal \N__66722\ : std_logic;
signal \N__66721\ : std_logic;
signal \N__66720\ : std_logic;
signal \N__66719\ : std_logic;
signal \N__66718\ : std_logic;
signal \N__66717\ : std_logic;
signal \N__66716\ : std_logic;
signal \N__66715\ : std_logic;
signal \N__66714\ : std_logic;
signal \N__66713\ : std_logic;
signal \N__66712\ : std_logic;
signal \N__66711\ : std_logic;
signal \N__66710\ : std_logic;
signal \N__66709\ : std_logic;
signal \N__66708\ : std_logic;
signal \N__66707\ : std_logic;
signal \N__66706\ : std_logic;
signal \N__66705\ : std_logic;
signal \N__66704\ : std_logic;
signal \N__66703\ : std_logic;
signal \N__66702\ : std_logic;
signal \N__66701\ : std_logic;
signal \N__66700\ : std_logic;
signal \N__66699\ : std_logic;
signal \N__66698\ : std_logic;
signal \N__66697\ : std_logic;
signal \N__66696\ : std_logic;
signal \N__66695\ : std_logic;
signal \N__66694\ : std_logic;
signal \N__66693\ : std_logic;
signal \N__66692\ : std_logic;
signal \N__66691\ : std_logic;
signal \N__66690\ : std_logic;
signal \N__66689\ : std_logic;
signal \N__66688\ : std_logic;
signal \N__66687\ : std_logic;
signal \N__66686\ : std_logic;
signal \N__66685\ : std_logic;
signal \N__66684\ : std_logic;
signal \N__66683\ : std_logic;
signal \N__66682\ : std_logic;
signal \N__66681\ : std_logic;
signal \N__66680\ : std_logic;
signal \N__66679\ : std_logic;
signal \N__66678\ : std_logic;
signal \N__66677\ : std_logic;
signal \N__66676\ : std_logic;
signal \N__66675\ : std_logic;
signal \N__66674\ : std_logic;
signal \N__66673\ : std_logic;
signal \N__66672\ : std_logic;
signal \N__66671\ : std_logic;
signal \N__66670\ : std_logic;
signal \N__66669\ : std_logic;
signal \N__66668\ : std_logic;
signal \N__66667\ : std_logic;
signal \N__66666\ : std_logic;
signal \N__66665\ : std_logic;
signal \N__66664\ : std_logic;
signal \N__66663\ : std_logic;
signal \N__66662\ : std_logic;
signal \N__66661\ : std_logic;
signal \N__66660\ : std_logic;
signal \N__66659\ : std_logic;
signal \N__66658\ : std_logic;
signal \N__66657\ : std_logic;
signal \N__66656\ : std_logic;
signal \N__66655\ : std_logic;
signal \N__66654\ : std_logic;
signal \N__66653\ : std_logic;
signal \N__66652\ : std_logic;
signal \N__66651\ : std_logic;
signal \N__66650\ : std_logic;
signal \N__66649\ : std_logic;
signal \N__66648\ : std_logic;
signal \N__66647\ : std_logic;
signal \N__66646\ : std_logic;
signal \N__66645\ : std_logic;
signal \N__66644\ : std_logic;
signal \N__66643\ : std_logic;
signal \N__66642\ : std_logic;
signal \N__66641\ : std_logic;
signal \N__66640\ : std_logic;
signal \N__66639\ : std_logic;
signal \N__66638\ : std_logic;
signal \N__66637\ : std_logic;
signal \N__66636\ : std_logic;
signal \N__66635\ : std_logic;
signal \N__66634\ : std_logic;
signal \N__66633\ : std_logic;
signal \N__66632\ : std_logic;
signal \N__66631\ : std_logic;
signal \N__66630\ : std_logic;
signal \N__66139\ : std_logic;
signal \N__66136\ : std_logic;
signal \N__66135\ : std_logic;
signal \N__66132\ : std_logic;
signal \N__66129\ : std_logic;
signal \N__66128\ : std_logic;
signal \N__66125\ : std_logic;
signal \N__66124\ : std_logic;
signal \N__66121\ : std_logic;
signal \N__66118\ : std_logic;
signal \N__66115\ : std_logic;
signal \N__66112\ : std_logic;
signal \N__66107\ : std_logic;
signal \N__66104\ : std_logic;
signal \N__66097\ : std_logic;
signal \N__66096\ : std_logic;
signal \N__66095\ : std_logic;
signal \N__66092\ : std_logic;
signal \N__66089\ : std_logic;
signal \N__66086\ : std_logic;
signal \N__66083\ : std_logic;
signal \N__66080\ : std_logic;
signal \N__66077\ : std_logic;
signal \N__66072\ : std_logic;
signal \N__66067\ : std_logic;
signal \N__66066\ : std_logic;
signal \N__66065\ : std_logic;
signal \N__66060\ : std_logic;
signal \N__66057\ : std_logic;
signal \N__66054\ : std_logic;
signal \N__66049\ : std_logic;
signal \N__66048\ : std_logic;
signal \N__66045\ : std_logic;
signal \N__66042\ : std_logic;
signal \N__66039\ : std_logic;
signal \N__66034\ : std_logic;
signal \N__66031\ : std_logic;
signal \N__66030\ : std_logic;
signal \N__66029\ : std_logic;
signal \N__66028\ : std_logic;
signal \N__66025\ : std_logic;
signal \N__66022\ : std_logic;
signal \N__66021\ : std_logic;
signal \N__66020\ : std_logic;
signal \N__66019\ : std_logic;
signal \N__66016\ : std_logic;
signal \N__66015\ : std_logic;
signal \N__66014\ : std_logic;
signal \N__66013\ : std_logic;
signal \N__66012\ : std_logic;
signal \N__66009\ : std_logic;
signal \N__66008\ : std_logic;
signal \N__66007\ : std_logic;
signal \N__66004\ : std_logic;
signal \N__66003\ : std_logic;
signal \N__66002\ : std_logic;
signal \N__66001\ : std_logic;
signal \N__65998\ : std_logic;
signal \N__65993\ : std_logic;
signal \N__65992\ : std_logic;
signal \N__65991\ : std_logic;
signal \N__65988\ : std_logic;
signal \N__65985\ : std_logic;
signal \N__65982\ : std_logic;
signal \N__65977\ : std_logic;
signal \N__65974\ : std_logic;
signal \N__65973\ : std_logic;
signal \N__65972\ : std_logic;
signal \N__65971\ : std_logic;
signal \N__65970\ : std_logic;
signal \N__65969\ : std_logic;
signal \N__65964\ : std_logic;
signal \N__65961\ : std_logic;
signal \N__65958\ : std_logic;
signal \N__65953\ : std_logic;
signal \N__65950\ : std_logic;
signal \N__65949\ : std_logic;
signal \N__65944\ : std_logic;
signal \N__65941\ : std_logic;
signal \N__65940\ : std_logic;
signal \N__65939\ : std_logic;
signal \N__65938\ : std_logic;
signal \N__65937\ : std_logic;
signal \N__65936\ : std_logic;
signal \N__65933\ : std_logic;
signal \N__65932\ : std_logic;
signal \N__65929\ : std_logic;
signal \N__65926\ : std_logic;
signal \N__65923\ : std_logic;
signal \N__65920\ : std_logic;
signal \N__65917\ : std_logic;
signal \N__65908\ : std_logic;
signal \N__65905\ : std_logic;
signal \N__65900\ : std_logic;
signal \N__65899\ : std_logic;
signal \N__65894\ : std_logic;
signal \N__65891\ : std_logic;
signal \N__65888\ : std_logic;
signal \N__65885\ : std_logic;
signal \N__65882\ : std_logic;
signal \N__65879\ : std_logic;
signal \N__65876\ : std_logic;
signal \N__65869\ : std_logic;
signal \N__65866\ : std_logic;
signal \N__65865\ : std_logic;
signal \N__65862\ : std_logic;
signal \N__65859\ : std_logic;
signal \N__65850\ : std_logic;
signal \N__65847\ : std_logic;
signal \N__65842\ : std_logic;
signal \N__65839\ : std_logic;
signal \N__65834\ : std_logic;
signal \N__65825\ : std_logic;
signal \N__65822\ : std_logic;
signal \N__65819\ : std_logic;
signal \N__65816\ : std_logic;
signal \N__65813\ : std_logic;
signal \N__65806\ : std_logic;
signal \N__65801\ : std_logic;
signal \N__65798\ : std_logic;
signal \N__65793\ : std_logic;
signal \N__65788\ : std_logic;
signal \N__65785\ : std_logic;
signal \N__65780\ : std_logic;
signal \N__65777\ : std_logic;
signal \N__65772\ : std_logic;
signal \N__65761\ : std_logic;
signal \N__65760\ : std_logic;
signal \N__65759\ : std_logic;
signal \N__65756\ : std_logic;
signal \N__65751\ : std_logic;
signal \N__65750\ : std_logic;
signal \N__65747\ : std_logic;
signal \N__65744\ : std_logic;
signal \N__65741\ : std_logic;
signal \N__65738\ : std_logic;
signal \N__65735\ : std_logic;
signal \N__65732\ : std_logic;
signal \N__65729\ : std_logic;
signal \N__65726\ : std_logic;
signal \N__65719\ : std_logic;
signal \N__65718\ : std_logic;
signal \N__65715\ : std_logic;
signal \N__65712\ : std_logic;
signal \N__65709\ : std_logic;
signal \N__65706\ : std_logic;
signal \N__65703\ : std_logic;
signal \N__65698\ : std_logic;
signal \N__65697\ : std_logic;
signal \N__65696\ : std_logic;
signal \N__65693\ : std_logic;
signal \N__65690\ : std_logic;
signal \N__65689\ : std_logic;
signal \N__65686\ : std_logic;
signal \N__65681\ : std_logic;
signal \N__65678\ : std_logic;
signal \N__65675\ : std_logic;
signal \N__65674\ : std_logic;
signal \N__65673\ : std_logic;
signal \N__65672\ : std_logic;
signal \N__65671\ : std_logic;
signal \N__65670\ : std_logic;
signal \N__65667\ : std_logic;
signal \N__65662\ : std_logic;
signal \N__65661\ : std_logic;
signal \N__65658\ : std_logic;
signal \N__65655\ : std_logic;
signal \N__65650\ : std_logic;
signal \N__65649\ : std_logic;
signal \N__65648\ : std_logic;
signal \N__65647\ : std_logic;
signal \N__65644\ : std_logic;
signal \N__65639\ : std_logic;
signal \N__65636\ : std_logic;
signal \N__65631\ : std_logic;
signal \N__65628\ : std_logic;
signal \N__65625\ : std_logic;
signal \N__65624\ : std_logic;
signal \N__65623\ : std_logic;
signal \N__65620\ : std_logic;
signal \N__65617\ : std_logic;
signal \N__65604\ : std_logic;
signal \N__65601\ : std_logic;
signal \N__65598\ : std_logic;
signal \N__65595\ : std_logic;
signal \N__65592\ : std_logic;
signal \N__65591\ : std_logic;
signal \N__65588\ : std_logic;
signal \N__65583\ : std_logic;
signal \N__65582\ : std_logic;
signal \N__65577\ : std_logic;
signal \N__65576\ : std_logic;
signal \N__65575\ : std_logic;
signal \N__65574\ : std_logic;
signal \N__65573\ : std_logic;
signal \N__65572\ : std_logic;
signal \N__65571\ : std_logic;
signal \N__65570\ : std_logic;
signal \N__65569\ : std_logic;
signal \N__65568\ : std_logic;
signal \N__65567\ : std_logic;
signal \N__65564\ : std_logic;
signal \N__65563\ : std_logic;
signal \N__65562\ : std_logic;
signal \N__65557\ : std_logic;
signal \N__65554\ : std_logic;
signal \N__65551\ : std_logic;
signal \N__65548\ : std_logic;
signal \N__65545\ : std_logic;
signal \N__65542\ : std_logic;
signal \N__65537\ : std_logic;
signal \N__65532\ : std_logic;
signal \N__65529\ : std_logic;
signal \N__65524\ : std_logic;
signal \N__65521\ : std_logic;
signal \N__65518\ : std_logic;
signal \N__65515\ : std_logic;
signal \N__65512\ : std_logic;
signal \N__65509\ : std_logic;
signal \N__65504\ : std_logic;
signal \N__65503\ : std_logic;
signal \N__65502\ : std_logic;
signal \N__65501\ : std_logic;
signal \N__65498\ : std_logic;
signal \N__65495\ : std_logic;
signal \N__65492\ : std_logic;
signal \N__65489\ : std_logic;
signal \N__65486\ : std_logic;
signal \N__65481\ : std_logic;
signal \N__65470\ : std_logic;
signal \N__65465\ : std_logic;
signal \N__65462\ : std_logic;
signal \N__65459\ : std_logic;
signal \N__65454\ : std_logic;
signal \N__65451\ : std_logic;
signal \N__65446\ : std_logic;
signal \N__65443\ : std_logic;
signal \N__65428\ : std_logic;
signal \N__65425\ : std_logic;
signal \N__65424\ : std_logic;
signal \N__65421\ : std_logic;
signal \N__65418\ : std_logic;
signal \N__65417\ : std_logic;
signal \N__65414\ : std_logic;
signal \N__65409\ : std_logic;
signal \N__65404\ : std_logic;
signal \N__65401\ : std_logic;
signal \N__65400\ : std_logic;
signal \N__65397\ : std_logic;
signal \N__65394\ : std_logic;
signal \N__65391\ : std_logic;
signal \N__65388\ : std_logic;
signal \N__65385\ : std_logic;
signal \N__65380\ : std_logic;
signal \N__65379\ : std_logic;
signal \N__65378\ : std_logic;
signal \N__65375\ : std_logic;
signal \N__65370\ : std_logic;
signal \N__65365\ : std_logic;
signal \N__65364\ : std_logic;
signal \N__65361\ : std_logic;
signal \N__65358\ : std_logic;
signal \N__65357\ : std_logic;
signal \N__65356\ : std_logic;
signal \N__65355\ : std_logic;
signal \N__65352\ : std_logic;
signal \N__65349\ : std_logic;
signal \N__65344\ : std_logic;
signal \N__65341\ : std_logic;
signal \N__65338\ : std_logic;
signal \N__65335\ : std_logic;
signal \N__65326\ : std_logic;
signal \N__65323\ : std_logic;
signal \N__65322\ : std_logic;
signal \N__65319\ : std_logic;
signal \N__65316\ : std_logic;
signal \N__65311\ : std_logic;
signal \N__65308\ : std_logic;
signal \N__65305\ : std_logic;
signal \N__65304\ : std_logic;
signal \N__65301\ : std_logic;
signal \N__65298\ : std_logic;
signal \N__65297\ : std_logic;
signal \N__65292\ : std_logic;
signal \N__65289\ : std_logic;
signal \N__65286\ : std_logic;
signal \N__65283\ : std_logic;
signal \N__65280\ : std_logic;
signal \N__65275\ : std_logic;
signal \N__65272\ : std_logic;
signal \N__65269\ : std_logic;
signal \N__65266\ : std_logic;
signal \N__65265\ : std_logic;
signal \N__65262\ : std_logic;
signal \N__65259\ : std_logic;
signal \N__65256\ : std_logic;
signal \N__65253\ : std_logic;
signal \N__65248\ : std_logic;
signal \N__65247\ : std_logic;
signal \N__65246\ : std_logic;
signal \N__65245\ : std_logic;
signal \N__65242\ : std_logic;
signal \N__65239\ : std_logic;
signal \N__65234\ : std_logic;
signal \N__65231\ : std_logic;
signal \N__65230\ : std_logic;
signal \N__65227\ : std_logic;
signal \N__65224\ : std_logic;
signal \N__65221\ : std_logic;
signal \N__65218\ : std_logic;
signal \N__65213\ : std_logic;
signal \N__65206\ : std_logic;
signal \N__65203\ : std_logic;
signal \N__65200\ : std_logic;
signal \N__65197\ : std_logic;
signal \N__65194\ : std_logic;
signal \N__65193\ : std_logic;
signal \N__65192\ : std_logic;
signal \N__65189\ : std_logic;
signal \N__65186\ : std_logic;
signal \N__65183\ : std_logic;
signal \N__65180\ : std_logic;
signal \N__65179\ : std_logic;
signal \N__65176\ : std_logic;
signal \N__65173\ : std_logic;
signal \N__65170\ : std_logic;
signal \N__65167\ : std_logic;
signal \N__65164\ : std_logic;
signal \N__65155\ : std_logic;
signal \N__65154\ : std_logic;
signal \N__65153\ : std_logic;
signal \N__65150\ : std_logic;
signal \N__65147\ : std_logic;
signal \N__65146\ : std_logic;
signal \N__65143\ : std_logic;
signal \N__65140\ : std_logic;
signal \N__65137\ : std_logic;
signal \N__65134\ : std_logic;
signal \N__65131\ : std_logic;
signal \N__65128\ : std_logic;
signal \N__65123\ : std_logic;
signal \N__65120\ : std_logic;
signal \N__65113\ : std_logic;
signal \N__65110\ : std_logic;
signal \N__65107\ : std_logic;
signal \N__65104\ : std_logic;
signal \N__65103\ : std_logic;
signal \N__65100\ : std_logic;
signal \N__65097\ : std_logic;
signal \N__65094\ : std_logic;
signal \N__65091\ : std_logic;
signal \N__65086\ : std_logic;
signal \N__65083\ : std_logic;
signal \N__65080\ : std_logic;
signal \N__65077\ : std_logic;
signal \N__65074\ : std_logic;
signal \N__65073\ : std_logic;
signal \N__65070\ : std_logic;
signal \N__65067\ : std_logic;
signal \N__65062\ : std_logic;
signal \N__65061\ : std_logic;
signal \N__65060\ : std_logic;
signal \N__65059\ : std_logic;
signal \N__65054\ : std_logic;
signal \N__65053\ : std_logic;
signal \N__65050\ : std_logic;
signal \N__65047\ : std_logic;
signal \N__65044\ : std_logic;
signal \N__65041\ : std_logic;
signal \N__65038\ : std_logic;
signal \N__65035\ : std_logic;
signal \N__65032\ : std_logic;
signal \N__65029\ : std_logic;
signal \N__65020\ : std_logic;
signal \N__65017\ : std_logic;
signal \N__65016\ : std_logic;
signal \N__65013\ : std_logic;
signal \N__65010\ : std_logic;
signal \N__65007\ : std_logic;
signal \N__65004\ : std_logic;
signal \N__65001\ : std_logic;
signal \N__64998\ : std_logic;
signal \N__64995\ : std_logic;
signal \N__64990\ : std_logic;
signal \N__64989\ : std_logic;
signal \N__64986\ : std_logic;
signal \N__64983\ : std_logic;
signal \N__64980\ : std_logic;
signal \N__64975\ : std_logic;
signal \N__64972\ : std_logic;
signal \N__64969\ : std_logic;
signal \N__64966\ : std_logic;
signal \N__64963\ : std_logic;
signal \N__64962\ : std_logic;
signal \N__64957\ : std_logic;
signal \N__64954\ : std_logic;
signal \N__64951\ : std_logic;
signal \N__64948\ : std_logic;
signal \N__64947\ : std_logic;
signal \N__64944\ : std_logic;
signal \N__64941\ : std_logic;
signal \N__64938\ : std_logic;
signal \N__64933\ : std_logic;
signal \N__64932\ : std_logic;
signal \N__64929\ : std_logic;
signal \N__64926\ : std_logic;
signal \N__64923\ : std_logic;
signal \N__64920\ : std_logic;
signal \N__64917\ : std_logic;
signal \N__64912\ : std_logic;
signal \N__64911\ : std_logic;
signal \N__64908\ : std_logic;
signal \N__64905\ : std_logic;
signal \N__64900\ : std_logic;
signal \N__64897\ : std_logic;
signal \N__64894\ : std_logic;
signal \N__64893\ : std_logic;
signal \N__64892\ : std_logic;
signal \N__64889\ : std_logic;
signal \N__64888\ : std_logic;
signal \N__64887\ : std_logic;
signal \N__64886\ : std_logic;
signal \N__64885\ : std_logic;
signal \N__64884\ : std_logic;
signal \N__64883\ : std_logic;
signal \N__64880\ : std_logic;
signal \N__64879\ : std_logic;
signal \N__64876\ : std_logic;
signal \N__64875\ : std_logic;
signal \N__64874\ : std_logic;
signal \N__64873\ : std_logic;
signal \N__64872\ : std_logic;
signal \N__64871\ : std_logic;
signal \N__64868\ : std_logic;
signal \N__64865\ : std_logic;
signal \N__64864\ : std_logic;
signal \N__64863\ : std_logic;
signal \N__64862\ : std_logic;
signal \N__64859\ : std_logic;
signal \N__64854\ : std_logic;
signal \N__64853\ : std_logic;
signal \N__64852\ : std_logic;
signal \N__64851\ : std_logic;
signal \N__64846\ : std_logic;
signal \N__64843\ : std_logic;
signal \N__64840\ : std_logic;
signal \N__64837\ : std_logic;
signal \N__64836\ : std_logic;
signal \N__64833\ : std_logic;
signal \N__64830\ : std_logic;
signal \N__64827\ : std_logic;
signal \N__64826\ : std_logic;
signal \N__64825\ : std_logic;
signal \N__64824\ : std_logic;
signal \N__64823\ : std_logic;
signal \N__64820\ : std_logic;
signal \N__64819\ : std_logic;
signal \N__64818\ : std_logic;
signal \N__64815\ : std_logic;
signal \N__64812\ : std_logic;
signal \N__64809\ : std_logic;
signal \N__64806\ : std_logic;
signal \N__64803\ : std_logic;
signal \N__64800\ : std_logic;
signal \N__64797\ : std_logic;
signal \N__64794\ : std_logic;
signal \N__64789\ : std_logic;
signal \N__64786\ : std_logic;
signal \N__64781\ : std_logic;
signal \N__64778\ : std_logic;
signal \N__64775\ : std_logic;
signal \N__64772\ : std_logic;
signal \N__64767\ : std_logic;
signal \N__64764\ : std_logic;
signal \N__64761\ : std_logic;
signal \N__64758\ : std_logic;
signal \N__64755\ : std_logic;
signal \N__64752\ : std_logic;
signal \N__64749\ : std_logic;
signal \N__64748\ : std_logic;
signal \N__64745\ : std_logic;
signal \N__64742\ : std_logic;
signal \N__64739\ : std_logic;
signal \N__64734\ : std_logic;
signal \N__64731\ : std_logic;
signal \N__64726\ : std_logic;
signal \N__64721\ : std_logic;
signal \N__64718\ : std_logic;
signal \N__64715\ : std_logic;
signal \N__64706\ : std_logic;
signal \N__64701\ : std_logic;
signal \N__64700\ : std_logic;
signal \N__64699\ : std_logic;
signal \N__64698\ : std_logic;
signal \N__64695\ : std_logic;
signal \N__64692\ : std_logic;
signal \N__64689\ : std_logic;
signal \N__64686\ : std_logic;
signal \N__64683\ : std_logic;
signal \N__64678\ : std_logic;
signal \N__64671\ : std_logic;
signal \N__64668\ : std_logic;
signal \N__64665\ : std_logic;
signal \N__64660\ : std_logic;
signal \N__64653\ : std_logic;
signal \N__64650\ : std_logic;
signal \N__64645\ : std_logic;
signal \N__64642\ : std_logic;
signal \N__64633\ : std_logic;
signal \N__64626\ : std_logic;
signal \N__64621\ : std_logic;
signal \N__64618\ : std_logic;
signal \N__64603\ : std_logic;
signal \N__64600\ : std_logic;
signal \N__64599\ : std_logic;
signal \N__64596\ : std_logic;
signal \N__64593\ : std_logic;
signal \N__64588\ : std_logic;
signal \N__64587\ : std_logic;
signal \N__64584\ : std_logic;
signal \N__64581\ : std_logic;
signal \N__64578\ : std_logic;
signal \N__64575\ : std_logic;
signal \N__64572\ : std_logic;
signal \N__64567\ : std_logic;
signal \N__64566\ : std_logic;
signal \N__64565\ : std_logic;
signal \N__64562\ : std_logic;
signal \N__64561\ : std_logic;
signal \N__64560\ : std_logic;
signal \N__64557\ : std_logic;
signal \N__64556\ : std_logic;
signal \N__64553\ : std_logic;
signal \N__64552\ : std_logic;
signal \N__64551\ : std_logic;
signal \N__64550\ : std_logic;
signal \N__64549\ : std_logic;
signal \N__64546\ : std_logic;
signal \N__64543\ : std_logic;
signal \N__64540\ : std_logic;
signal \N__64537\ : std_logic;
signal \N__64536\ : std_logic;
signal \N__64535\ : std_logic;
signal \N__64534\ : std_logic;
signal \N__64533\ : std_logic;
signal \N__64532\ : std_logic;
signal \N__64531\ : std_logic;
signal \N__64528\ : std_logic;
signal \N__64527\ : std_logic;
signal \N__64524\ : std_logic;
signal \N__64523\ : std_logic;
signal \N__64520\ : std_logic;
signal \N__64519\ : std_logic;
signal \N__64518\ : std_logic;
signal \N__64517\ : std_logic;
signal \N__64514\ : std_logic;
signal \N__64513\ : std_logic;
signal \N__64512\ : std_logic;
signal \N__64511\ : std_logic;
signal \N__64508\ : std_logic;
signal \N__64505\ : std_logic;
signal \N__64502\ : std_logic;
signal \N__64499\ : std_logic;
signal \N__64498\ : std_logic;
signal \N__64495\ : std_logic;
signal \N__64492\ : std_logic;
signal \N__64487\ : std_logic;
signal \N__64482\ : std_logic;
signal \N__64481\ : std_logic;
signal \N__64478\ : std_logic;
signal \N__64473\ : std_logic;
signal \N__64470\ : std_logic;
signal \N__64467\ : std_logic;
signal \N__64464\ : std_logic;
signal \N__64459\ : std_logic;
signal \N__64458\ : std_logic;
signal \N__64455\ : std_logic;
signal \N__64452\ : std_logic;
signal \N__64451\ : std_logic;
signal \N__64448\ : std_logic;
signal \N__64441\ : std_logic;
signal \N__64438\ : std_logic;
signal \N__64435\ : std_logic;
signal \N__64430\ : std_logic;
signal \N__64427\ : std_logic;
signal \N__64420\ : std_logic;
signal \N__64417\ : std_logic;
signal \N__64414\ : std_logic;
signal \N__64411\ : std_logic;
signal \N__64404\ : std_logic;
signal \N__64399\ : std_logic;
signal \N__64396\ : std_logic;
signal \N__64391\ : std_logic;
signal \N__64388\ : std_logic;
signal \N__64385\ : std_logic;
signal \N__64382\ : std_logic;
signal \N__64375\ : std_logic;
signal \N__64372\ : std_logic;
signal \N__64365\ : std_logic;
signal \N__64358\ : std_logic;
signal \N__64357\ : std_logic;
signal \N__64356\ : std_logic;
signal \N__64353\ : std_logic;
signal \N__64350\ : std_logic;
signal \N__64347\ : std_logic;
signal \N__64346\ : std_logic;
signal \N__64345\ : std_logic;
signal \N__64342\ : std_logic;
signal \N__64339\ : std_logic;
signal \N__64336\ : std_logic;
signal \N__64333\ : std_logic;
signal \N__64328\ : std_logic;
signal \N__64323\ : std_logic;
signal \N__64316\ : std_logic;
signal \N__64313\ : std_logic;
signal \N__64310\ : std_logic;
signal \N__64305\ : std_logic;
signal \N__64302\ : std_logic;
signal \N__64299\ : std_logic;
signal \N__64296\ : std_logic;
signal \N__64291\ : std_logic;
signal \N__64276\ : std_logic;
signal \N__64275\ : std_logic;
signal \N__64272\ : std_logic;
signal \N__64269\ : std_logic;
signal \N__64266\ : std_logic;
signal \N__64263\ : std_logic;
signal \N__64258\ : std_logic;
signal \N__64257\ : std_logic;
signal \N__64254\ : std_logic;
signal \N__64251\ : std_logic;
signal \N__64248\ : std_logic;
signal \N__64245\ : std_logic;
signal \N__64244\ : std_logic;
signal \N__64239\ : std_logic;
signal \N__64236\ : std_logic;
signal \N__64231\ : std_logic;
signal \N__64228\ : std_logic;
signal \N__64225\ : std_logic;
signal \N__64224\ : std_logic;
signal \N__64221\ : std_logic;
signal \N__64220\ : std_logic;
signal \N__64219\ : std_logic;
signal \N__64216\ : std_logic;
signal \N__64213\ : std_logic;
signal \N__64208\ : std_logic;
signal \N__64207\ : std_logic;
signal \N__64204\ : std_logic;
signal \N__64199\ : std_logic;
signal \N__64196\ : std_logic;
signal \N__64189\ : std_logic;
signal \N__64186\ : std_logic;
signal \N__64183\ : std_logic;
signal \N__64180\ : std_logic;
signal \N__64177\ : std_logic;
signal \N__64174\ : std_logic;
signal \N__64173\ : std_logic;
signal \N__64170\ : std_logic;
signal \N__64167\ : std_logic;
signal \N__64164\ : std_logic;
signal \N__64161\ : std_logic;
signal \N__64156\ : std_logic;
signal \N__64153\ : std_logic;
signal \N__64152\ : std_logic;
signal \N__64149\ : std_logic;
signal \N__64146\ : std_logic;
signal \N__64141\ : std_logic;
signal \N__64138\ : std_logic;
signal \N__64135\ : std_logic;
signal \N__64132\ : std_logic;
signal \N__64129\ : std_logic;
signal \N__64126\ : std_logic;
signal \N__64123\ : std_logic;
signal \N__64122\ : std_logic;
signal \N__64119\ : std_logic;
signal \N__64116\ : std_logic;
signal \N__64111\ : std_logic;
signal \N__64110\ : std_logic;
signal \N__64109\ : std_logic;
signal \N__64106\ : std_logic;
signal \N__64101\ : std_logic;
signal \N__64098\ : std_logic;
signal \N__64095\ : std_logic;
signal \N__64092\ : std_logic;
signal \N__64089\ : std_logic;
signal \N__64084\ : std_logic;
signal \N__64081\ : std_logic;
signal \N__64078\ : std_logic;
signal \N__64075\ : std_logic;
signal \N__64072\ : std_logic;
signal \N__64069\ : std_logic;
signal \N__64066\ : std_logic;
signal \N__64065\ : std_logic;
signal \N__64062\ : std_logic;
signal \N__64059\ : std_logic;
signal \N__64054\ : std_logic;
signal \N__64051\ : std_logic;
signal \N__64048\ : std_logic;
signal \N__64045\ : std_logic;
signal \N__64042\ : std_logic;
signal \N__64039\ : std_logic;
signal \N__64036\ : std_logic;
signal \N__64035\ : std_logic;
signal \N__64034\ : std_logic;
signal \N__64031\ : std_logic;
signal \N__64030\ : std_logic;
signal \N__64027\ : std_logic;
signal \N__64024\ : std_logic;
signal \N__64021\ : std_logic;
signal \N__64018\ : std_logic;
signal \N__64017\ : std_logic;
signal \N__64014\ : std_logic;
signal \N__64011\ : std_logic;
signal \N__64008\ : std_logic;
signal \N__64003\ : std_logic;
signal \N__63994\ : std_logic;
signal \N__63991\ : std_logic;
signal \N__63988\ : std_logic;
signal \N__63985\ : std_logic;
signal \N__63982\ : std_logic;
signal \N__63979\ : std_logic;
signal \N__63976\ : std_logic;
signal \N__63973\ : std_logic;
signal \N__63970\ : std_logic;
signal \N__63969\ : std_logic;
signal \N__63966\ : std_logic;
signal \N__63963\ : std_logic;
signal \N__63958\ : std_logic;
signal \N__63957\ : std_logic;
signal \N__63956\ : std_logic;
signal \N__63953\ : std_logic;
signal \N__63950\ : std_logic;
signal \N__63947\ : std_logic;
signal \N__63944\ : std_logic;
signal \N__63941\ : std_logic;
signal \N__63938\ : std_logic;
signal \N__63935\ : std_logic;
signal \N__63932\ : std_logic;
signal \N__63929\ : std_logic;
signal \N__63922\ : std_logic;
signal \N__63919\ : std_logic;
signal \N__63918\ : std_logic;
signal \N__63917\ : std_logic;
signal \N__63914\ : std_logic;
signal \N__63911\ : std_logic;
signal \N__63908\ : std_logic;
signal \N__63905\ : std_logic;
signal \N__63902\ : std_logic;
signal \N__63901\ : std_logic;
signal \N__63900\ : std_logic;
signal \N__63897\ : std_logic;
signal \N__63894\ : std_logic;
signal \N__63891\ : std_logic;
signal \N__63886\ : std_logic;
signal \N__63877\ : std_logic;
signal \N__63876\ : std_logic;
signal \N__63873\ : std_logic;
signal \N__63870\ : std_logic;
signal \N__63865\ : std_logic;
signal \N__63864\ : std_logic;
signal \N__63863\ : std_logic;
signal \N__63862\ : std_logic;
signal \N__63861\ : std_logic;
signal \N__63860\ : std_logic;
signal \N__63859\ : std_logic;
signal \N__63856\ : std_logic;
signal \N__63855\ : std_logic;
signal \N__63854\ : std_logic;
signal \N__63853\ : std_logic;
signal \N__63852\ : std_logic;
signal \N__63851\ : std_logic;
signal \N__63850\ : std_logic;
signal \N__63849\ : std_logic;
signal \N__63846\ : std_logic;
signal \N__63843\ : std_logic;
signal \N__63840\ : std_logic;
signal \N__63835\ : std_logic;
signal \N__63832\ : std_logic;
signal \N__63831\ : std_logic;
signal \N__63830\ : std_logic;
signal \N__63827\ : std_logic;
signal \N__63826\ : std_logic;
signal \N__63825\ : std_logic;
signal \N__63820\ : std_logic;
signal \N__63817\ : std_logic;
signal \N__63816\ : std_logic;
signal \N__63815\ : std_logic;
signal \N__63814\ : std_logic;
signal \N__63813\ : std_logic;
signal \N__63810\ : std_logic;
signal \N__63807\ : std_logic;
signal \N__63804\ : std_logic;
signal \N__63801\ : std_logic;
signal \N__63800\ : std_logic;
signal \N__63797\ : std_logic;
signal \N__63794\ : std_logic;
signal \N__63793\ : std_logic;
signal \N__63790\ : std_logic;
signal \N__63785\ : std_logic;
signal \N__63782\ : std_logic;
signal \N__63781\ : std_logic;
signal \N__63780\ : std_logic;
signal \N__63779\ : std_logic;
signal \N__63776\ : std_logic;
signal \N__63773\ : std_logic;
signal \N__63770\ : std_logic;
signal \N__63769\ : std_logic;
signal \N__63768\ : std_logic;
signal \N__63765\ : std_logic;
signal \N__63764\ : std_logic;
signal \N__63761\ : std_logic;
signal \N__63758\ : std_logic;
signal \N__63753\ : std_logic;
signal \N__63750\ : std_logic;
signal \N__63747\ : std_logic;
signal \N__63744\ : std_logic;
signal \N__63741\ : std_logic;
signal \N__63738\ : std_logic;
signal \N__63735\ : std_logic;
signal \N__63732\ : std_logic;
signal \N__63727\ : std_logic;
signal \N__63724\ : std_logic;
signal \N__63717\ : std_logic;
signal \N__63716\ : std_logic;
signal \N__63713\ : std_logic;
signal \N__63710\ : std_logic;
signal \N__63707\ : std_logic;
signal \N__63700\ : std_logic;
signal \N__63695\ : std_logic;
signal \N__63692\ : std_logic;
signal \N__63689\ : std_logic;
signal \N__63686\ : std_logic;
signal \N__63679\ : std_logic;
signal \N__63672\ : std_logic;
signal \N__63665\ : std_logic;
signal \N__63660\ : std_logic;
signal \N__63657\ : std_logic;
signal \N__63654\ : std_logic;
signal \N__63651\ : std_logic;
signal \N__63644\ : std_logic;
signal \N__63643\ : std_logic;
signal \N__63638\ : std_logic;
signal \N__63633\ : std_logic;
signal \N__63626\ : std_logic;
signal \N__63623\ : std_logic;
signal \N__63620\ : std_logic;
signal \N__63617\ : std_logic;
signal \N__63612\ : std_logic;
signal \N__63609\ : std_logic;
signal \N__63606\ : std_logic;
signal \N__63603\ : std_logic;
signal \N__63600\ : std_logic;
signal \N__63597\ : std_logic;
signal \N__63592\ : std_logic;
signal \N__63589\ : std_logic;
signal \N__63574\ : std_logic;
signal \N__63573\ : std_logic;
signal \N__63570\ : std_logic;
signal \N__63567\ : std_logic;
signal \N__63564\ : std_logic;
signal \N__63561\ : std_logic;
signal \N__63560\ : std_logic;
signal \N__63555\ : std_logic;
signal \N__63552\ : std_logic;
signal \N__63547\ : std_logic;
signal \N__63546\ : std_logic;
signal \N__63543\ : std_logic;
signal \N__63540\ : std_logic;
signal \N__63539\ : std_logic;
signal \N__63538\ : std_logic;
signal \N__63535\ : std_logic;
signal \N__63532\ : std_logic;
signal \N__63529\ : std_logic;
signal \N__63526\ : std_logic;
signal \N__63523\ : std_logic;
signal \N__63520\ : std_logic;
signal \N__63517\ : std_logic;
signal \N__63510\ : std_logic;
signal \N__63505\ : std_logic;
signal \N__63502\ : std_logic;
signal \N__63501\ : std_logic;
signal \N__63498\ : std_logic;
signal \N__63495\ : std_logic;
signal \N__63490\ : std_logic;
signal \N__63487\ : std_logic;
signal \N__63486\ : std_logic;
signal \N__63485\ : std_logic;
signal \N__63482\ : std_logic;
signal \N__63479\ : std_logic;
signal \N__63476\ : std_logic;
signal \N__63475\ : std_logic;
signal \N__63470\ : std_logic;
signal \N__63467\ : std_logic;
signal \N__63464\ : std_logic;
signal \N__63459\ : std_logic;
signal \N__63456\ : std_logic;
signal \N__63455\ : std_logic;
signal \N__63450\ : std_logic;
signal \N__63447\ : std_logic;
signal \N__63444\ : std_logic;
signal \N__63439\ : std_logic;
signal \N__63436\ : std_logic;
signal \N__63433\ : std_logic;
signal \N__63432\ : std_logic;
signal \N__63429\ : std_logic;
signal \N__63426\ : std_logic;
signal \N__63421\ : std_logic;
signal \N__63418\ : std_logic;
signal \N__63417\ : std_logic;
signal \N__63416\ : std_logic;
signal \N__63413\ : std_logic;
signal \N__63410\ : std_logic;
signal \N__63407\ : std_logic;
signal \N__63404\ : std_logic;
signal \N__63401\ : std_logic;
signal \N__63398\ : std_logic;
signal \N__63395\ : std_logic;
signal \N__63388\ : std_logic;
signal \N__63387\ : std_logic;
signal \N__63384\ : std_logic;
signal \N__63381\ : std_logic;
signal \N__63378\ : std_logic;
signal \N__63375\ : std_logic;
signal \N__63372\ : std_logic;
signal \N__63369\ : std_logic;
signal \N__63364\ : std_logic;
signal \N__63361\ : std_logic;
signal \N__63358\ : std_logic;
signal \N__63357\ : std_logic;
signal \N__63356\ : std_logic;
signal \N__63355\ : std_logic;
signal \N__63352\ : std_logic;
signal \N__63351\ : std_logic;
signal \N__63348\ : std_logic;
signal \N__63345\ : std_logic;
signal \N__63342\ : std_logic;
signal \N__63339\ : std_logic;
signal \N__63336\ : std_logic;
signal \N__63331\ : std_logic;
signal \N__63328\ : std_logic;
signal \N__63321\ : std_logic;
signal \N__63316\ : std_logic;
signal \N__63313\ : std_logic;
signal \N__63310\ : std_logic;
signal \N__63309\ : std_logic;
signal \N__63308\ : std_logic;
signal \N__63305\ : std_logic;
signal \N__63304\ : std_logic;
signal \N__63301\ : std_logic;
signal \N__63296\ : std_logic;
signal \N__63295\ : std_logic;
signal \N__63292\ : std_logic;
signal \N__63289\ : std_logic;
signal \N__63286\ : std_logic;
signal \N__63283\ : std_logic;
signal \N__63280\ : std_logic;
signal \N__63275\ : std_logic;
signal \N__63268\ : std_logic;
signal \N__63267\ : std_logic;
signal \N__63264\ : std_logic;
signal \N__63261\ : std_logic;
signal \N__63258\ : std_logic;
signal \N__63257\ : std_logic;
signal \N__63254\ : std_logic;
signal \N__63251\ : std_logic;
signal \N__63248\ : std_logic;
signal \N__63245\ : std_logic;
signal \N__63238\ : std_logic;
signal \N__63235\ : std_logic;
signal \N__63232\ : std_logic;
signal \N__63229\ : std_logic;
signal \N__63226\ : std_logic;
signal \N__63225\ : std_logic;
signal \N__63222\ : std_logic;
signal \N__63219\ : std_logic;
signal \N__63218\ : std_logic;
signal \N__63217\ : std_logic;
signal \N__63216\ : std_logic;
signal \N__63213\ : std_logic;
signal \N__63210\ : std_logic;
signal \N__63207\ : std_logic;
signal \N__63206\ : std_logic;
signal \N__63205\ : std_logic;
signal \N__63204\ : std_logic;
signal \N__63201\ : std_logic;
signal \N__63198\ : std_logic;
signal \N__63195\ : std_logic;
signal \N__63192\ : std_logic;
signal \N__63189\ : std_logic;
signal \N__63188\ : std_logic;
signal \N__63185\ : std_logic;
signal \N__63182\ : std_logic;
signal \N__63179\ : std_logic;
signal \N__63178\ : std_logic;
signal \N__63177\ : std_logic;
signal \N__63176\ : std_logic;
signal \N__63175\ : std_logic;
signal \N__63174\ : std_logic;
signal \N__63173\ : std_logic;
signal \N__63172\ : std_logic;
signal \N__63171\ : std_logic;
signal \N__63170\ : std_logic;
signal \N__63165\ : std_logic;
signal \N__63162\ : std_logic;
signal \N__63161\ : std_logic;
signal \N__63156\ : std_logic;
signal \N__63153\ : std_logic;
signal \N__63150\ : std_logic;
signal \N__63147\ : std_logic;
signal \N__63146\ : std_logic;
signal \N__63145\ : std_logic;
signal \N__63144\ : std_logic;
signal \N__63143\ : std_logic;
signal \N__63140\ : std_logic;
signal \N__63139\ : std_logic;
signal \N__63136\ : std_logic;
signal \N__63133\ : std_logic;
signal \N__63130\ : std_logic;
signal \N__63125\ : std_logic;
signal \N__63124\ : std_logic;
signal \N__63123\ : std_logic;
signal \N__63120\ : std_logic;
signal \N__63117\ : std_logic;
signal \N__63114\ : std_logic;
signal \N__63111\ : std_logic;
signal \N__63108\ : std_logic;
signal \N__63107\ : std_logic;
signal \N__63106\ : std_logic;
signal \N__63103\ : std_logic;
signal \N__63100\ : std_logic;
signal \N__63093\ : std_logic;
signal \N__63092\ : std_logic;
signal \N__63089\ : std_logic;
signal \N__63086\ : std_logic;
signal \N__63083\ : std_logic;
signal \N__63078\ : std_logic;
signal \N__63075\ : std_logic;
signal \N__63072\ : std_logic;
signal \N__63069\ : std_logic;
signal \N__63062\ : std_logic;
signal \N__63059\ : std_logic;
signal \N__63058\ : std_logic;
signal \N__63055\ : std_logic;
signal \N__63052\ : std_logic;
signal \N__63049\ : std_logic;
signal \N__63046\ : std_logic;
signal \N__63041\ : std_logic;
signal \N__63038\ : std_logic;
signal \N__63035\ : std_logic;
signal \N__63030\ : std_logic;
signal \N__63027\ : std_logic;
signal \N__63024\ : std_logic;
signal \N__63021\ : std_logic;
signal \N__63018\ : std_logic;
signal \N__63015\ : std_logic;
signal \N__63010\ : std_logic;
signal \N__63001\ : std_logic;
signal \N__63000\ : std_logic;
signal \N__62997\ : std_logic;
signal \N__62990\ : std_logic;
signal \N__62985\ : std_logic;
signal \N__62982\ : std_logic;
signal \N__62979\ : std_logic;
signal \N__62976\ : std_logic;
signal \N__62975\ : std_logic;
signal \N__62972\ : std_logic;
signal \N__62967\ : std_logic;
signal \N__62964\ : std_logic;
signal \N__62961\ : std_logic;
signal \N__62956\ : std_logic;
signal \N__62953\ : std_logic;
signal \N__62944\ : std_logic;
signal \N__62941\ : std_logic;
signal \N__62938\ : std_logic;
signal \N__62935\ : std_logic;
signal \N__62932\ : std_logic;
signal \N__62929\ : std_logic;
signal \N__62922\ : std_logic;
signal \N__62913\ : std_logic;
signal \N__62902\ : std_logic;
signal \N__62901\ : std_logic;
signal \N__62900\ : std_logic;
signal \N__62897\ : std_logic;
signal \N__62894\ : std_logic;
signal \N__62893\ : std_logic;
signal \N__62890\ : std_logic;
signal \N__62887\ : std_logic;
signal \N__62884\ : std_logic;
signal \N__62881\ : std_logic;
signal \N__62874\ : std_logic;
signal \N__62869\ : std_logic;
signal \N__62866\ : std_logic;
signal \N__62863\ : std_logic;
signal \N__62860\ : std_logic;
signal \N__62857\ : std_logic;
signal \N__62854\ : std_logic;
signal \N__62851\ : std_logic;
signal \N__62850\ : std_logic;
signal \N__62847\ : std_logic;
signal \N__62844\ : std_logic;
signal \N__62839\ : std_logic;
signal \N__62836\ : std_logic;
signal \N__62833\ : std_logic;
signal \N__62830\ : std_logic;
signal \N__62827\ : std_logic;
signal \N__62826\ : std_logic;
signal \N__62823\ : std_logic;
signal \N__62822\ : std_logic;
signal \N__62819\ : std_logic;
signal \N__62816\ : std_logic;
signal \N__62815\ : std_logic;
signal \N__62812\ : std_logic;
signal \N__62807\ : std_logic;
signal \N__62804\ : std_logic;
signal \N__62801\ : std_logic;
signal \N__62798\ : std_logic;
signal \N__62791\ : std_logic;
signal \N__62788\ : std_logic;
signal \N__62787\ : std_logic;
signal \N__62784\ : std_logic;
signal \N__62781\ : std_logic;
signal \N__62778\ : std_logic;
signal \N__62775\ : std_logic;
signal \N__62770\ : std_logic;
signal \N__62767\ : std_logic;
signal \N__62766\ : std_logic;
signal \N__62765\ : std_logic;
signal \N__62762\ : std_logic;
signal \N__62757\ : std_logic;
signal \N__62752\ : std_logic;
signal \N__62751\ : std_logic;
signal \N__62748\ : std_logic;
signal \N__62745\ : std_logic;
signal \N__62742\ : std_logic;
signal \N__62739\ : std_logic;
signal \N__62736\ : std_logic;
signal \N__62733\ : std_logic;
signal \N__62730\ : std_logic;
signal \N__62729\ : std_logic;
signal \N__62726\ : std_logic;
signal \N__62723\ : std_logic;
signal \N__62720\ : std_logic;
signal \N__62717\ : std_logic;
signal \N__62714\ : std_logic;
signal \N__62707\ : std_logic;
signal \N__62706\ : std_logic;
signal \N__62703\ : std_logic;
signal \N__62702\ : std_logic;
signal \N__62699\ : std_logic;
signal \N__62698\ : std_logic;
signal \N__62695\ : std_logic;
signal \N__62690\ : std_logic;
signal \N__62687\ : std_logic;
signal \N__62682\ : std_logic;
signal \N__62677\ : std_logic;
signal \N__62676\ : std_logic;
signal \N__62673\ : std_logic;
signal \N__62672\ : std_logic;
signal \N__62671\ : std_logic;
signal \N__62668\ : std_logic;
signal \N__62665\ : std_logic;
signal \N__62662\ : std_logic;
signal \N__62661\ : std_logic;
signal \N__62658\ : std_logic;
signal \N__62655\ : std_logic;
signal \N__62650\ : std_logic;
signal \N__62647\ : std_logic;
signal \N__62644\ : std_logic;
signal \N__62635\ : std_logic;
signal \N__62632\ : std_logic;
signal \N__62631\ : std_logic;
signal \N__62630\ : std_logic;
signal \N__62627\ : std_logic;
signal \N__62624\ : std_logic;
signal \N__62621\ : std_logic;
signal \N__62618\ : std_logic;
signal \N__62615\ : std_logic;
signal \N__62612\ : std_logic;
signal \N__62609\ : std_logic;
signal \N__62606\ : std_logic;
signal \N__62599\ : std_logic;
signal \N__62598\ : std_logic;
signal \N__62595\ : std_logic;
signal \N__62592\ : std_logic;
signal \N__62591\ : std_logic;
signal \N__62590\ : std_logic;
signal \N__62587\ : std_logic;
signal \N__62584\ : std_logic;
signal \N__62581\ : std_logic;
signal \N__62578\ : std_logic;
signal \N__62573\ : std_logic;
signal \N__62570\ : std_logic;
signal \N__62567\ : std_logic;
signal \N__62564\ : std_logic;
signal \N__62557\ : std_logic;
signal \N__62556\ : std_logic;
signal \N__62555\ : std_logic;
signal \N__62554\ : std_logic;
signal \N__62551\ : std_logic;
signal \N__62546\ : std_logic;
signal \N__62545\ : std_logic;
signal \N__62544\ : std_logic;
signal \N__62543\ : std_logic;
signal \N__62542\ : std_logic;
signal \N__62541\ : std_logic;
signal \N__62540\ : std_logic;
signal \N__62539\ : std_logic;
signal \N__62538\ : std_logic;
signal \N__62535\ : std_logic;
signal \N__62532\ : std_logic;
signal \N__62531\ : std_logic;
signal \N__62530\ : std_logic;
signal \N__62529\ : std_logic;
signal \N__62528\ : std_logic;
signal \N__62527\ : std_logic;
signal \N__62526\ : std_logic;
signal \N__62525\ : std_logic;
signal \N__62524\ : std_logic;
signal \N__62523\ : std_logic;
signal \N__62522\ : std_logic;
signal \N__62519\ : std_logic;
signal \N__62514\ : std_logic;
signal \N__62511\ : std_logic;
signal \N__62510\ : std_logic;
signal \N__62509\ : std_logic;
signal \N__62508\ : std_logic;
signal \N__62507\ : std_logic;
signal \N__62506\ : std_logic;
signal \N__62505\ : std_logic;
signal \N__62504\ : std_logic;
signal \N__62503\ : std_logic;
signal \N__62502\ : std_logic;
signal \N__62501\ : std_logic;
signal \N__62500\ : std_logic;
signal \N__62499\ : std_logic;
signal \N__62498\ : std_logic;
signal \N__62497\ : std_logic;
signal \N__62496\ : std_logic;
signal \N__62495\ : std_logic;
signal \N__62494\ : std_logic;
signal \N__62493\ : std_logic;
signal \N__62492\ : std_logic;
signal \N__62491\ : std_logic;
signal \N__62490\ : std_logic;
signal \N__62487\ : std_logic;
signal \N__62484\ : std_logic;
signal \N__62477\ : std_logic;
signal \N__62472\ : std_logic;
signal \N__62465\ : std_logic;
signal \N__62458\ : std_logic;
signal \N__62449\ : std_logic;
signal \N__62444\ : std_logic;
signal \N__62441\ : std_logic;
signal \N__62436\ : std_logic;
signal \N__62433\ : std_logic;
signal \N__62432\ : std_logic;
signal \N__62431\ : std_logic;
signal \N__62430\ : std_logic;
signal \N__62429\ : std_logic;
signal \N__62428\ : std_logic;
signal \N__62427\ : std_logic;
signal \N__62422\ : std_logic;
signal \N__62417\ : std_logic;
signal \N__62412\ : std_logic;
signal \N__62409\ : std_logic;
signal \N__62406\ : std_logic;
signal \N__62397\ : std_logic;
signal \N__62396\ : std_logic;
signal \N__62383\ : std_logic;
signal \N__62380\ : std_logic;
signal \N__62379\ : std_logic;
signal \N__62378\ : std_logic;
signal \N__62377\ : std_logic;
signal \N__62376\ : std_logic;
signal \N__62375\ : std_logic;
signal \N__62374\ : std_logic;
signal \N__62365\ : std_logic;
signal \N__62360\ : std_logic;
signal \N__62357\ : std_logic;
signal \N__62352\ : std_logic;
signal \N__62351\ : std_logic;
signal \N__62348\ : std_logic;
signal \N__62343\ : std_logic;
signal \N__62340\ : std_logic;
signal \N__62333\ : std_logic;
signal \N__62330\ : std_logic;
signal \N__62327\ : std_logic;
signal \N__62324\ : std_logic;
signal \N__62317\ : std_logic;
signal \N__62314\ : std_logic;
signal \N__62311\ : std_logic;
signal \N__62308\ : std_logic;
signal \N__62305\ : std_logic;
signal \N__62302\ : std_logic;
signal \N__62299\ : std_logic;
signal \N__62292\ : std_logic;
signal \N__62289\ : std_logic;
signal \N__62282\ : std_logic;
signal \N__62279\ : std_logic;
signal \N__62276\ : std_logic;
signal \N__62273\ : std_logic;
signal \N__62260\ : std_logic;
signal \N__62257\ : std_logic;
signal \N__62252\ : std_logic;
signal \N__62249\ : std_logic;
signal \N__62236\ : std_logic;
signal \N__62233\ : std_logic;
signal \N__62230\ : std_logic;
signal \N__62227\ : std_logic;
signal \N__62222\ : std_logic;
signal \N__62217\ : std_logic;
signal \N__62206\ : std_logic;
signal \N__62205\ : std_logic;
signal \N__62204\ : std_logic;
signal \N__62203\ : std_logic;
signal \N__62202\ : std_logic;
signal \N__62199\ : std_logic;
signal \N__62198\ : std_logic;
signal \N__62197\ : std_logic;
signal \N__62194\ : std_logic;
signal \N__62191\ : std_logic;
signal \N__62190\ : std_logic;
signal \N__62189\ : std_logic;
signal \N__62188\ : std_logic;
signal \N__62187\ : std_logic;
signal \N__62186\ : std_logic;
signal \N__62185\ : std_logic;
signal \N__62184\ : std_logic;
signal \N__62183\ : std_logic;
signal \N__62182\ : std_logic;
signal \N__62181\ : std_logic;
signal \N__62178\ : std_logic;
signal \N__62177\ : std_logic;
signal \N__62174\ : std_logic;
signal \N__62171\ : std_logic;
signal \N__62168\ : std_logic;
signal \N__62167\ : std_logic;
signal \N__62166\ : std_logic;
signal \N__62161\ : std_logic;
signal \N__62160\ : std_logic;
signal \N__62157\ : std_logic;
signal \N__62154\ : std_logic;
signal \N__62151\ : std_logic;
signal \N__62150\ : std_logic;
signal \N__62149\ : std_logic;
signal \N__62148\ : std_logic;
signal \N__62145\ : std_logic;
signal \N__62142\ : std_logic;
signal \N__62137\ : std_logic;
signal \N__62132\ : std_logic;
signal \N__62125\ : std_logic;
signal \N__62122\ : std_logic;
signal \N__62121\ : std_logic;
signal \N__62120\ : std_logic;
signal \N__62117\ : std_logic;
signal \N__62112\ : std_logic;
signal \N__62107\ : std_logic;
signal \N__62104\ : std_logic;
signal \N__62101\ : std_logic;
signal \N__62098\ : std_logic;
signal \N__62095\ : std_logic;
signal \N__62092\ : std_logic;
signal \N__62089\ : std_logic;
signal \N__62088\ : std_logic;
signal \N__62087\ : std_logic;
signal \N__62086\ : std_logic;
signal \N__62083\ : std_logic;
signal \N__62080\ : std_logic;
signal \N__62077\ : std_logic;
signal \N__62074\ : std_logic;
signal \N__62071\ : std_logic;
signal \N__62068\ : std_logic;
signal \N__62065\ : std_logic;
signal \N__62062\ : std_logic;
signal \N__62059\ : std_logic;
signal \N__62058\ : std_logic;
signal \N__62055\ : std_logic;
signal \N__62052\ : std_logic;
signal \N__62049\ : std_logic;
signal \N__62046\ : std_logic;
signal \N__62043\ : std_logic;
signal \N__62038\ : std_logic;
signal \N__62033\ : std_logic;
signal \N__62030\ : std_logic;
signal \N__62027\ : std_logic;
signal \N__62024\ : std_logic;
signal \N__62021\ : std_logic;
signal \N__62018\ : std_logic;
signal \N__62015\ : std_logic;
signal \N__62010\ : std_logic;
signal \N__62007\ : std_logic;
signal \N__62004\ : std_logic;
signal \N__62001\ : std_logic;
signal \N__61998\ : std_logic;
signal \N__61995\ : std_logic;
signal \N__61992\ : std_logic;
signal \N__61989\ : std_logic;
signal \N__61982\ : std_logic;
signal \N__61977\ : std_logic;
signal \N__61974\ : std_logic;
signal \N__61971\ : std_logic;
signal \N__61970\ : std_logic;
signal \N__61969\ : std_logic;
signal \N__61966\ : std_logic;
signal \N__61961\ : std_logic;
signal \N__61950\ : std_logic;
signal \N__61945\ : std_logic;
signal \N__61934\ : std_logic;
signal \N__61929\ : std_logic;
signal \N__61924\ : std_logic;
signal \N__61921\ : std_logic;
signal \N__61918\ : std_logic;
signal \N__61915\ : std_logic;
signal \N__61910\ : std_logic;
signal \N__61907\ : std_logic;
signal \N__61894\ : std_logic;
signal \N__61891\ : std_logic;
signal \N__61888\ : std_logic;
signal \N__61887\ : std_logic;
signal \N__61886\ : std_logic;
signal \N__61885\ : std_logic;
signal \N__61884\ : std_logic;
signal \N__61881\ : std_logic;
signal \N__61878\ : std_logic;
signal \N__61875\ : std_logic;
signal \N__61872\ : std_logic;
signal \N__61869\ : std_logic;
signal \N__61866\ : std_logic;
signal \N__61861\ : std_logic;
signal \N__61852\ : std_logic;
signal \N__61849\ : std_logic;
signal \N__61848\ : std_logic;
signal \N__61845\ : std_logic;
signal \N__61842\ : std_logic;
signal \N__61839\ : std_logic;
signal \N__61836\ : std_logic;
signal \N__61833\ : std_logic;
signal \N__61828\ : std_logic;
signal \N__61825\ : std_logic;
signal \N__61824\ : std_logic;
signal \N__61823\ : std_logic;
signal \N__61820\ : std_logic;
signal \N__61817\ : std_logic;
signal \N__61814\ : std_logic;
signal \N__61813\ : std_logic;
signal \N__61808\ : std_logic;
signal \N__61807\ : std_logic;
signal \N__61804\ : std_logic;
signal \N__61801\ : std_logic;
signal \N__61798\ : std_logic;
signal \N__61795\ : std_logic;
signal \N__61786\ : std_logic;
signal \N__61783\ : std_logic;
signal \N__61780\ : std_logic;
signal \N__61777\ : std_logic;
signal \N__61774\ : std_logic;
signal \N__61773\ : std_logic;
signal \N__61770\ : std_logic;
signal \N__61767\ : std_logic;
signal \N__61764\ : std_logic;
signal \N__61763\ : std_logic;
signal \N__61760\ : std_logic;
signal \N__61757\ : std_logic;
signal \N__61754\ : std_logic;
signal \N__61747\ : std_logic;
signal \N__61746\ : std_logic;
signal \N__61745\ : std_logic;
signal \N__61742\ : std_logic;
signal \N__61741\ : std_logic;
signal \N__61738\ : std_logic;
signal \N__61737\ : std_logic;
signal \N__61734\ : std_logic;
signal \N__61731\ : std_logic;
signal \N__61728\ : std_logic;
signal \N__61725\ : std_logic;
signal \N__61722\ : std_logic;
signal \N__61715\ : std_logic;
signal \N__61708\ : std_logic;
signal \N__61705\ : std_logic;
signal \N__61702\ : std_logic;
signal \N__61699\ : std_logic;
signal \N__61696\ : std_logic;
signal \N__61695\ : std_logic;
signal \N__61694\ : std_logic;
signal \N__61691\ : std_logic;
signal \N__61688\ : std_logic;
signal \N__61685\ : std_logic;
signal \N__61682\ : std_logic;
signal \N__61679\ : std_logic;
signal \N__61672\ : std_logic;
signal \N__61669\ : std_logic;
signal \N__61668\ : std_logic;
signal \N__61667\ : std_logic;
signal \N__61666\ : std_logic;
signal \N__61663\ : std_logic;
signal \N__61660\ : std_logic;
signal \N__61655\ : std_logic;
signal \N__61652\ : std_logic;
signal \N__61647\ : std_logic;
signal \N__61642\ : std_logic;
signal \N__61641\ : std_logic;
signal \N__61638\ : std_logic;
signal \N__61635\ : std_logic;
signal \N__61632\ : std_logic;
signal \N__61629\ : std_logic;
signal \N__61626\ : std_logic;
signal \N__61623\ : std_logic;
signal \N__61618\ : std_logic;
signal \N__61617\ : std_logic;
signal \N__61616\ : std_logic;
signal \N__61615\ : std_logic;
signal \N__61612\ : std_logic;
signal \N__61609\ : std_logic;
signal \N__61604\ : std_logic;
signal \N__61603\ : std_logic;
signal \N__61600\ : std_logic;
signal \N__61597\ : std_logic;
signal \N__61594\ : std_logic;
signal \N__61591\ : std_logic;
signal \N__61588\ : std_logic;
signal \N__61579\ : std_logic;
signal \N__61578\ : std_logic;
signal \N__61575\ : std_logic;
signal \N__61572\ : std_logic;
signal \N__61569\ : std_logic;
signal \N__61566\ : std_logic;
signal \N__61561\ : std_logic;
signal \N__61558\ : std_logic;
signal \N__61555\ : std_logic;
signal \N__61552\ : std_logic;
signal \N__61549\ : std_logic;
signal \N__61546\ : std_logic;
signal \N__61543\ : std_logic;
signal \N__61542\ : std_logic;
signal \N__61539\ : std_logic;
signal \N__61536\ : std_logic;
signal \N__61533\ : std_logic;
signal \N__61530\ : std_logic;
signal \N__61525\ : std_logic;
signal \N__61522\ : std_logic;
signal \N__61519\ : std_logic;
signal \N__61518\ : std_logic;
signal \N__61517\ : std_logic;
signal \N__61514\ : std_logic;
signal \N__61511\ : std_logic;
signal \N__61508\ : std_logic;
signal \N__61501\ : std_logic;
signal \N__61500\ : std_logic;
signal \N__61497\ : std_logic;
signal \N__61496\ : std_logic;
signal \N__61493\ : std_logic;
signal \N__61488\ : std_logic;
signal \N__61485\ : std_logic;
signal \N__61482\ : std_logic;
signal \N__61481\ : std_logic;
signal \N__61476\ : std_logic;
signal \N__61473\ : std_logic;
signal \N__61468\ : std_logic;
signal \N__61467\ : std_logic;
signal \N__61464\ : std_logic;
signal \N__61461\ : std_logic;
signal \N__61458\ : std_logic;
signal \N__61455\ : std_logic;
signal \N__61452\ : std_logic;
signal \N__61449\ : std_logic;
signal \N__61448\ : std_logic;
signal \N__61443\ : std_logic;
signal \N__61440\ : std_logic;
signal \N__61435\ : std_logic;
signal \N__61434\ : std_logic;
signal \N__61431\ : std_logic;
signal \N__61430\ : std_logic;
signal \N__61427\ : std_logic;
signal \N__61424\ : std_logic;
signal \N__61421\ : std_logic;
signal \N__61420\ : std_logic;
signal \N__61417\ : std_logic;
signal \N__61416\ : std_logic;
signal \N__61415\ : std_logic;
signal \N__61410\ : std_logic;
signal \N__61407\ : std_logic;
signal \N__61404\ : std_logic;
signal \N__61399\ : std_logic;
signal \N__61390\ : std_logic;
signal \N__61389\ : std_logic;
signal \N__61386\ : std_logic;
signal \N__61383\ : std_logic;
signal \N__61382\ : std_logic;
signal \N__61379\ : std_logic;
signal \N__61376\ : std_logic;
signal \N__61373\ : std_logic;
signal \N__61370\ : std_logic;
signal \N__61367\ : std_logic;
signal \N__61360\ : std_logic;
signal \N__61359\ : std_logic;
signal \N__61356\ : std_logic;
signal \N__61353\ : std_logic;
signal \N__61350\ : std_logic;
signal \N__61347\ : std_logic;
signal \N__61344\ : std_logic;
signal \N__61343\ : std_logic;
signal \N__61338\ : std_logic;
signal \N__61335\ : std_logic;
signal \N__61330\ : std_logic;
signal \N__61329\ : std_logic;
signal \N__61326\ : std_logic;
signal \N__61323\ : std_logic;
signal \N__61322\ : std_logic;
signal \N__61319\ : std_logic;
signal \N__61316\ : std_logic;
signal \N__61313\ : std_logic;
signal \N__61312\ : std_logic;
signal \N__61307\ : std_logic;
signal \N__61304\ : std_logic;
signal \N__61301\ : std_logic;
signal \N__61294\ : std_logic;
signal \N__61291\ : std_logic;
signal \N__61290\ : std_logic;
signal \N__61289\ : std_logic;
signal \N__61286\ : std_logic;
signal \N__61285\ : std_logic;
signal \N__61284\ : std_logic;
signal \N__61281\ : std_logic;
signal \N__61278\ : std_logic;
signal \N__61275\ : std_logic;
signal \N__61268\ : std_logic;
signal \N__61261\ : std_logic;
signal \N__61258\ : std_logic;
signal \N__61255\ : std_logic;
signal \N__61254\ : std_logic;
signal \N__61251\ : std_logic;
signal \N__61248\ : std_logic;
signal \N__61243\ : std_logic;
signal \N__61242\ : std_logic;
signal \N__61239\ : std_logic;
signal \N__61236\ : std_logic;
signal \N__61235\ : std_logic;
signal \N__61232\ : std_logic;
signal \N__61229\ : std_logic;
signal \N__61226\ : std_logic;
signal \N__61219\ : std_logic;
signal \N__61216\ : std_logic;
signal \N__61213\ : std_logic;
signal \N__61210\ : std_logic;
signal \N__61209\ : std_logic;
signal \N__61206\ : std_logic;
signal \N__61203\ : std_logic;
signal \N__61202\ : std_logic;
signal \N__61199\ : std_logic;
signal \N__61196\ : std_logic;
signal \N__61193\ : std_logic;
signal \N__61188\ : std_logic;
signal \N__61185\ : std_logic;
signal \N__61182\ : std_logic;
signal \N__61177\ : std_logic;
signal \N__61176\ : std_logic;
signal \N__61173\ : std_logic;
signal \N__61172\ : std_logic;
signal \N__61169\ : std_logic;
signal \N__61166\ : std_logic;
signal \N__61163\ : std_logic;
signal \N__61156\ : std_logic;
signal \N__61153\ : std_logic;
signal \N__61150\ : std_logic;
signal \N__61149\ : std_logic;
signal \N__61146\ : std_logic;
signal \N__61143\ : std_logic;
signal \N__61138\ : std_logic;
signal \N__61135\ : std_logic;
signal \N__61132\ : std_logic;
signal \N__61131\ : std_logic;
signal \N__61128\ : std_logic;
signal \N__61125\ : std_logic;
signal \N__61124\ : std_logic;
signal \N__61119\ : std_logic;
signal \N__61116\ : std_logic;
signal \N__61111\ : std_logic;
signal \N__61108\ : std_logic;
signal \N__61107\ : std_logic;
signal \N__61104\ : std_logic;
signal \N__61103\ : std_logic;
signal \N__61100\ : std_logic;
signal \N__61097\ : std_logic;
signal \N__61094\ : std_logic;
signal \N__61093\ : std_logic;
signal \N__61092\ : std_logic;
signal \N__61089\ : std_logic;
signal \N__61084\ : std_logic;
signal \N__61079\ : std_logic;
signal \N__61072\ : std_logic;
signal \N__61069\ : std_logic;
signal \N__61066\ : std_logic;
signal \N__61063\ : std_logic;
signal \N__61062\ : std_logic;
signal \N__61059\ : std_logic;
signal \N__61056\ : std_logic;
signal \N__61051\ : std_logic;
signal \N__61048\ : std_logic;
signal \N__61045\ : std_logic;
signal \N__61044\ : std_logic;
signal \N__61041\ : std_logic;
signal \N__61040\ : std_logic;
signal \N__61037\ : std_logic;
signal \N__61032\ : std_logic;
signal \N__61027\ : std_logic;
signal \N__61024\ : std_logic;
signal \N__61023\ : std_logic;
signal \N__61020\ : std_logic;
signal \N__61017\ : std_logic;
signal \N__61014\ : std_logic;
signal \N__61011\ : std_logic;
signal \N__61008\ : std_logic;
signal \N__61003\ : std_logic;
signal \N__61000\ : std_logic;
signal \N__60997\ : std_logic;
signal \N__60996\ : std_logic;
signal \N__60993\ : std_logic;
signal \N__60990\ : std_logic;
signal \N__60989\ : std_logic;
signal \N__60986\ : std_logic;
signal \N__60983\ : std_logic;
signal \N__60980\ : std_logic;
signal \N__60973\ : std_logic;
signal \N__60972\ : std_logic;
signal \N__60969\ : std_logic;
signal \N__60966\ : std_logic;
signal \N__60963\ : std_logic;
signal \N__60958\ : std_logic;
signal \N__60955\ : std_logic;
signal \N__60952\ : std_logic;
signal \N__60949\ : std_logic;
signal \N__60948\ : std_logic;
signal \N__60947\ : std_logic;
signal \N__60944\ : std_logic;
signal \N__60941\ : std_logic;
signal \N__60938\ : std_logic;
signal \N__60937\ : std_logic;
signal \N__60934\ : std_logic;
signal \N__60931\ : std_logic;
signal \N__60928\ : std_logic;
signal \N__60925\ : std_logic;
signal \N__60922\ : std_logic;
signal \N__60915\ : std_logic;
signal \N__60912\ : std_logic;
signal \N__60907\ : std_logic;
signal \N__60904\ : std_logic;
signal \N__60901\ : std_logic;
signal \N__60898\ : std_logic;
signal \N__60897\ : std_logic;
signal \N__60896\ : std_logic;
signal \N__60895\ : std_logic;
signal \N__60894\ : std_logic;
signal \N__60893\ : std_logic;
signal \N__60892\ : std_logic;
signal \N__60891\ : std_logic;
signal \N__60890\ : std_logic;
signal \N__60889\ : std_logic;
signal \N__60888\ : std_logic;
signal \N__60887\ : std_logic;
signal \N__60884\ : std_logic;
signal \N__60883\ : std_logic;
signal \N__60882\ : std_logic;
signal \N__60881\ : std_logic;
signal \N__60878\ : std_logic;
signal \N__60871\ : std_logic;
signal \N__60870\ : std_logic;
signal \N__60869\ : std_logic;
signal \N__60868\ : std_logic;
signal \N__60867\ : std_logic;
signal \N__60864\ : std_logic;
signal \N__60863\ : std_logic;
signal \N__60856\ : std_logic;
signal \N__60853\ : std_logic;
signal \N__60852\ : std_logic;
signal \N__60851\ : std_logic;
signal \N__60850\ : std_logic;
signal \N__60849\ : std_logic;
signal \N__60848\ : std_logic;
signal \N__60847\ : std_logic;
signal \N__60846\ : std_logic;
signal \N__60845\ : std_logic;
signal \N__60844\ : std_logic;
signal \N__60843\ : std_logic;
signal \N__60842\ : std_logic;
signal \N__60839\ : std_logic;
signal \N__60836\ : std_logic;
signal \N__60835\ : std_logic;
signal \N__60834\ : std_logic;
signal \N__60831\ : std_logic;
signal \N__60824\ : std_logic;
signal \N__60823\ : std_logic;
signal \N__60820\ : std_logic;
signal \N__60817\ : std_logic;
signal \N__60808\ : std_logic;
signal \N__60807\ : std_logic;
signal \N__60806\ : std_logic;
signal \N__60803\ : std_logic;
signal \N__60800\ : std_logic;
signal \N__60795\ : std_logic;
signal \N__60784\ : std_logic;
signal \N__60777\ : std_logic;
signal \N__60770\ : std_logic;
signal \N__60767\ : std_logic;
signal \N__60766\ : std_logic;
signal \N__60765\ : std_logic;
signal \N__60764\ : std_logic;
signal \N__60763\ : std_logic;
signal \N__60762\ : std_logic;
signal \N__60761\ : std_logic;
signal \N__60760\ : std_logic;
signal \N__60759\ : std_logic;
signal \N__60758\ : std_logic;
signal \N__60757\ : std_logic;
signal \N__60756\ : std_logic;
signal \N__60755\ : std_logic;
signal \N__60752\ : std_logic;
signal \N__60747\ : std_logic;
signal \N__60742\ : std_logic;
signal \N__60739\ : std_logic;
signal \N__60734\ : std_logic;
signal \N__60731\ : std_logic;
signal \N__60728\ : std_logic;
signal \N__60727\ : std_logic;
signal \N__60724\ : std_logic;
signal \N__60719\ : std_logic;
signal \N__60716\ : std_logic;
signal \N__60715\ : std_logic;
signal \N__60714\ : std_logic;
signal \N__60713\ : std_logic;
signal \N__60708\ : std_logic;
signal \N__60703\ : std_logic;
signal \N__60688\ : std_logic;
signal \N__60685\ : std_logic;
signal \N__60676\ : std_logic;
signal \N__60673\ : std_logic;
signal \N__60668\ : std_logic;
signal \N__60661\ : std_logic;
signal \N__60658\ : std_logic;
signal \N__60655\ : std_logic;
signal \N__60652\ : std_logic;
signal \N__60649\ : std_logic;
signal \N__60646\ : std_logic;
signal \N__60645\ : std_logic;
signal \N__60644\ : std_logic;
signal \N__60643\ : std_logic;
signal \N__60642\ : std_logic;
signal \N__60639\ : std_logic;
signal \N__60634\ : std_logic;
signal \N__60629\ : std_logic;
signal \N__60624\ : std_logic;
signal \N__60617\ : std_logic;
signal \N__60614\ : std_logic;
signal \N__60611\ : std_logic;
signal \N__60602\ : std_logic;
signal \N__60593\ : std_logic;
signal \N__60574\ : std_logic;
signal \N__60571\ : std_logic;
signal \N__60568\ : std_logic;
signal \N__60567\ : std_logic;
signal \N__60566\ : std_logic;
signal \N__60563\ : std_logic;
signal \N__60558\ : std_logic;
signal \N__60553\ : std_logic;
signal \N__60550\ : std_logic;
signal \N__60547\ : std_logic;
signal \N__60546\ : std_logic;
signal \N__60543\ : std_logic;
signal \N__60540\ : std_logic;
signal \N__60535\ : std_logic;
signal \N__60532\ : std_logic;
signal \N__60531\ : std_logic;
signal \N__60528\ : std_logic;
signal \N__60525\ : std_logic;
signal \N__60520\ : std_logic;
signal \N__60519\ : std_logic;
signal \N__60516\ : std_logic;
signal \N__60513\ : std_logic;
signal \N__60512\ : std_logic;
signal \N__60511\ : std_logic;
signal \N__60508\ : std_logic;
signal \N__60503\ : std_logic;
signal \N__60500\ : std_logic;
signal \N__60497\ : std_logic;
signal \N__60490\ : std_logic;
signal \N__60489\ : std_logic;
signal \N__60486\ : std_logic;
signal \N__60483\ : std_logic;
signal \N__60482\ : std_logic;
signal \N__60479\ : std_logic;
signal \N__60476\ : std_logic;
signal \N__60473\ : std_logic;
signal \N__60470\ : std_logic;
signal \N__60467\ : std_logic;
signal \N__60464\ : std_logic;
signal \N__60461\ : std_logic;
signal \N__60458\ : std_logic;
signal \N__60451\ : std_logic;
signal \N__60450\ : std_logic;
signal \N__60447\ : std_logic;
signal \N__60444\ : std_logic;
signal \N__60441\ : std_logic;
signal \N__60436\ : std_logic;
signal \N__60435\ : std_logic;
signal \N__60432\ : std_logic;
signal \N__60429\ : std_logic;
signal \N__60426\ : std_logic;
signal \N__60421\ : std_logic;
signal \N__60418\ : std_logic;
signal \N__60415\ : std_logic;
signal \N__60412\ : std_logic;
signal \N__60409\ : std_logic;
signal \N__60406\ : std_logic;
signal \N__60403\ : std_logic;
signal \N__60400\ : std_logic;
signal \N__60399\ : std_logic;
signal \N__60398\ : std_logic;
signal \N__60395\ : std_logic;
signal \N__60392\ : std_logic;
signal \N__60389\ : std_logic;
signal \N__60384\ : std_logic;
signal \N__60383\ : std_logic;
signal \N__60380\ : std_logic;
signal \N__60377\ : std_logic;
signal \N__60374\ : std_logic;
signal \N__60367\ : std_logic;
signal \N__60364\ : std_logic;
signal \N__60363\ : std_logic;
signal \N__60360\ : std_logic;
signal \N__60357\ : std_logic;
signal \N__60356\ : std_logic;
signal \N__60351\ : std_logic;
signal \N__60348\ : std_logic;
signal \N__60345\ : std_logic;
signal \N__60340\ : std_logic;
signal \N__60337\ : std_logic;
signal \N__60334\ : std_logic;
signal \N__60333\ : std_logic;
signal \N__60330\ : std_logic;
signal \N__60329\ : std_logic;
signal \N__60326\ : std_logic;
signal \N__60323\ : std_logic;
signal \N__60320\ : std_logic;
signal \N__60313\ : std_logic;
signal \N__60312\ : std_logic;
signal \N__60311\ : std_logic;
signal \N__60310\ : std_logic;
signal \N__60305\ : std_logic;
signal \N__60302\ : std_logic;
signal \N__60299\ : std_logic;
signal \N__60296\ : std_logic;
signal \N__60293\ : std_logic;
signal \N__60290\ : std_logic;
signal \N__60287\ : std_logic;
signal \N__60284\ : std_logic;
signal \N__60277\ : std_logic;
signal \N__60274\ : std_logic;
signal \N__60271\ : std_logic;
signal \N__60268\ : std_logic;
signal \N__60265\ : std_logic;
signal \N__60262\ : std_logic;
signal \N__60259\ : std_logic;
signal \N__60256\ : std_logic;
signal \N__60255\ : std_logic;
signal \N__60254\ : std_logic;
signal \N__60253\ : std_logic;
signal \N__60250\ : std_logic;
signal \N__60245\ : std_logic;
signal \N__60242\ : std_logic;
signal \N__60235\ : std_logic;
signal \N__60234\ : std_logic;
signal \N__60233\ : std_logic;
signal \N__60232\ : std_logic;
signal \N__60229\ : std_logic;
signal \N__60226\ : std_logic;
signal \N__60223\ : std_logic;
signal \N__60220\ : std_logic;
signal \N__60211\ : std_logic;
signal \N__60208\ : std_logic;
signal \N__60207\ : std_logic;
signal \N__60204\ : std_logic;
signal \N__60201\ : std_logic;
signal \N__60196\ : std_logic;
signal \N__60195\ : std_logic;
signal \N__60192\ : std_logic;
signal \N__60191\ : std_logic;
signal \N__60188\ : std_logic;
signal \N__60185\ : std_logic;
signal \N__60182\ : std_logic;
signal \N__60179\ : std_logic;
signal \N__60176\ : std_logic;
signal \N__60173\ : std_logic;
signal \N__60172\ : std_logic;
signal \N__60169\ : std_logic;
signal \N__60164\ : std_logic;
signal \N__60161\ : std_logic;
signal \N__60154\ : std_logic;
signal \N__60151\ : std_logic;
signal \N__60150\ : std_logic;
signal \N__60147\ : std_logic;
signal \N__60144\ : std_logic;
signal \N__60143\ : std_logic;
signal \N__60140\ : std_logic;
signal \N__60139\ : std_logic;
signal \N__60134\ : std_logic;
signal \N__60131\ : std_logic;
signal \N__60128\ : std_logic;
signal \N__60121\ : std_logic;
signal \N__60118\ : std_logic;
signal \N__60117\ : std_logic;
signal \N__60114\ : std_logic;
signal \N__60111\ : std_logic;
signal \N__60108\ : std_logic;
signal \N__60103\ : std_logic;
signal \N__60102\ : std_logic;
signal \N__60101\ : std_logic;
signal \N__60098\ : std_logic;
signal \N__60095\ : std_logic;
signal \N__60094\ : std_logic;
signal \N__60091\ : std_logic;
signal \N__60088\ : std_logic;
signal \N__60085\ : std_logic;
signal \N__60082\ : std_logic;
signal \N__60081\ : std_logic;
signal \N__60078\ : std_logic;
signal \N__60073\ : std_logic;
signal \N__60068\ : std_logic;
signal \N__60061\ : std_logic;
signal \N__60058\ : std_logic;
signal \N__60055\ : std_logic;
signal \N__60054\ : std_logic;
signal \N__60051\ : std_logic;
signal \N__60048\ : std_logic;
signal \N__60045\ : std_logic;
signal \N__60042\ : std_logic;
signal \N__60037\ : std_logic;
signal \N__60034\ : std_logic;
signal \N__60031\ : std_logic;
signal \N__60030\ : std_logic;
signal \N__60027\ : std_logic;
signal \N__60024\ : std_logic;
signal \N__60021\ : std_logic;
signal \N__60018\ : std_logic;
signal \N__60015\ : std_logic;
signal \N__60012\ : std_logic;
signal \N__60007\ : std_logic;
signal \N__60004\ : std_logic;
signal \N__60003\ : std_logic;
signal \N__60002\ : std_logic;
signal \N__59999\ : std_logic;
signal \N__59996\ : std_logic;
signal \N__59993\ : std_logic;
signal \N__59990\ : std_logic;
signal \N__59983\ : std_logic;
signal \N__59980\ : std_logic;
signal \N__59977\ : std_logic;
signal \N__59976\ : std_logic;
signal \N__59973\ : std_logic;
signal \N__59970\ : std_logic;
signal \N__59965\ : std_logic;
signal \N__59962\ : std_logic;
signal \N__59959\ : std_logic;
signal \N__59958\ : std_logic;
signal \N__59957\ : std_logic;
signal \N__59954\ : std_logic;
signal \N__59949\ : std_logic;
signal \N__59944\ : std_logic;
signal \N__59941\ : std_logic;
signal \N__59940\ : std_logic;
signal \N__59939\ : std_logic;
signal \N__59936\ : std_logic;
signal \N__59933\ : std_logic;
signal \N__59930\ : std_logic;
signal \N__59925\ : std_logic;
signal \N__59922\ : std_logic;
signal \N__59919\ : std_logic;
signal \N__59914\ : std_logic;
signal \N__59911\ : std_logic;
signal \N__59910\ : std_logic;
signal \N__59907\ : std_logic;
signal \N__59904\ : std_logic;
signal \N__59899\ : std_logic;
signal \N__59898\ : std_logic;
signal \N__59897\ : std_logic;
signal \N__59894\ : std_logic;
signal \N__59889\ : std_logic;
signal \N__59884\ : std_logic;
signal \N__59883\ : std_logic;
signal \N__59880\ : std_logic;
signal \N__59877\ : std_logic;
signal \N__59874\ : std_logic;
signal \N__59869\ : std_logic;
signal \N__59868\ : std_logic;
signal \N__59865\ : std_logic;
signal \N__59864\ : std_logic;
signal \N__59863\ : std_logic;
signal \N__59860\ : std_logic;
signal \N__59859\ : std_logic;
signal \N__59856\ : std_logic;
signal \N__59853\ : std_logic;
signal \N__59850\ : std_logic;
signal \N__59845\ : std_logic;
signal \N__59842\ : std_logic;
signal \N__59833\ : std_logic;
signal \N__59832\ : std_logic;
signal \N__59829\ : std_logic;
signal \N__59826\ : std_logic;
signal \N__59823\ : std_logic;
signal \N__59820\ : std_logic;
signal \N__59817\ : std_logic;
signal \N__59812\ : std_logic;
signal \N__59811\ : std_logic;
signal \N__59808\ : std_logic;
signal \N__59805\ : std_logic;
signal \N__59802\ : std_logic;
signal \N__59797\ : std_logic;
signal \N__59794\ : std_logic;
signal \N__59791\ : std_logic;
signal \N__59788\ : std_logic;
signal \N__59787\ : std_logic;
signal \N__59784\ : std_logic;
signal \N__59781\ : std_logic;
signal \N__59778\ : std_logic;
signal \N__59775\ : std_logic;
signal \N__59770\ : std_logic;
signal \N__59767\ : std_logic;
signal \N__59764\ : std_logic;
signal \N__59761\ : std_logic;
signal \N__59758\ : std_logic;
signal \N__59757\ : std_logic;
signal \N__59756\ : std_logic;
signal \N__59753\ : std_logic;
signal \N__59752\ : std_logic;
signal \N__59751\ : std_logic;
signal \N__59750\ : std_logic;
signal \N__59749\ : std_logic;
signal \N__59748\ : std_logic;
signal \N__59747\ : std_logic;
signal \N__59740\ : std_logic;
signal \N__59733\ : std_logic;
signal \N__59728\ : std_logic;
signal \N__59725\ : std_logic;
signal \N__59716\ : std_logic;
signal \N__59715\ : std_logic;
signal \N__59712\ : std_logic;
signal \N__59711\ : std_logic;
signal \N__59710\ : std_logic;
signal \N__59709\ : std_logic;
signal \N__59708\ : std_logic;
signal \N__59705\ : std_logic;
signal \N__59700\ : std_logic;
signal \N__59699\ : std_logic;
signal \N__59698\ : std_logic;
signal \N__59695\ : std_logic;
signal \N__59694\ : std_logic;
signal \N__59691\ : std_logic;
signal \N__59690\ : std_logic;
signal \N__59685\ : std_logic;
signal \N__59682\ : std_logic;
signal \N__59677\ : std_logic;
signal \N__59672\ : std_logic;
signal \N__59669\ : std_logic;
signal \N__59666\ : std_logic;
signal \N__59659\ : std_logic;
signal \N__59656\ : std_logic;
signal \N__59655\ : std_logic;
signal \N__59654\ : std_logic;
signal \N__59653\ : std_logic;
signal \N__59650\ : std_logic;
signal \N__59647\ : std_logic;
signal \N__59644\ : std_logic;
signal \N__59641\ : std_logic;
signal \N__59634\ : std_logic;
signal \N__59631\ : std_logic;
signal \N__59628\ : std_logic;
signal \N__59625\ : std_logic;
signal \N__59620\ : std_logic;
signal \N__59617\ : std_logic;
signal \N__59610\ : std_logic;
signal \N__59607\ : std_logic;
signal \N__59604\ : std_logic;
signal \N__59601\ : std_logic;
signal \N__59598\ : std_logic;
signal \N__59593\ : std_logic;
signal \N__59592\ : std_logic;
signal \N__59589\ : std_logic;
signal \N__59584\ : std_logic;
signal \N__59581\ : std_logic;
signal \N__59580\ : std_logic;
signal \N__59579\ : std_logic;
signal \N__59578\ : std_logic;
signal \N__59575\ : std_logic;
signal \N__59572\ : std_logic;
signal \N__59569\ : std_logic;
signal \N__59566\ : std_logic;
signal \N__59563\ : std_logic;
signal \N__59558\ : std_logic;
signal \N__59555\ : std_logic;
signal \N__59552\ : std_logic;
signal \N__59549\ : std_logic;
signal \N__59542\ : std_logic;
signal \N__59541\ : std_logic;
signal \N__59538\ : std_logic;
signal \N__59535\ : std_logic;
signal \N__59534\ : std_logic;
signal \N__59533\ : std_logic;
signal \N__59528\ : std_logic;
signal \N__59523\ : std_logic;
signal \N__59522\ : std_logic;
signal \N__59517\ : std_logic;
signal \N__59514\ : std_logic;
signal \N__59511\ : std_logic;
signal \N__59508\ : std_logic;
signal \N__59505\ : std_logic;
signal \N__59500\ : std_logic;
signal \N__59499\ : std_logic;
signal \N__59496\ : std_logic;
signal \N__59493\ : std_logic;
signal \N__59490\ : std_logic;
signal \N__59489\ : std_logic;
signal \N__59488\ : std_logic;
signal \N__59485\ : std_logic;
signal \N__59482\ : std_logic;
signal \N__59477\ : std_logic;
signal \N__59470\ : std_logic;
signal \N__59467\ : std_logic;
signal \N__59464\ : std_logic;
signal \N__59461\ : std_logic;
signal \N__59458\ : std_logic;
signal \N__59455\ : std_logic;
signal \N__59452\ : std_logic;
signal \N__59449\ : std_logic;
signal \N__59446\ : std_logic;
signal \N__59445\ : std_logic;
signal \N__59440\ : std_logic;
signal \N__59439\ : std_logic;
signal \N__59436\ : std_logic;
signal \N__59433\ : std_logic;
signal \N__59430\ : std_logic;
signal \N__59427\ : std_logic;
signal \N__59424\ : std_logic;
signal \N__59419\ : std_logic;
signal \N__59416\ : std_logic;
signal \N__59413\ : std_logic;
signal \N__59410\ : std_logic;
signal \N__59409\ : std_logic;
signal \N__59408\ : std_logic;
signal \N__59407\ : std_logic;
signal \N__59402\ : std_logic;
signal \N__59401\ : std_logic;
signal \N__59400\ : std_logic;
signal \N__59397\ : std_logic;
signal \N__59394\ : std_logic;
signal \N__59393\ : std_logic;
signal \N__59390\ : std_logic;
signal \N__59385\ : std_logic;
signal \N__59382\ : std_logic;
signal \N__59377\ : std_logic;
signal \N__59372\ : std_logic;
signal \N__59365\ : std_logic;
signal \N__59362\ : std_logic;
signal \N__59359\ : std_logic;
signal \N__59356\ : std_logic;
signal \N__59353\ : std_logic;
signal \N__59352\ : std_logic;
signal \N__59349\ : std_logic;
signal \N__59346\ : std_logic;
signal \N__59343\ : std_logic;
signal \N__59340\ : std_logic;
signal \N__59337\ : std_logic;
signal \N__59336\ : std_logic;
signal \N__59335\ : std_logic;
signal \N__59332\ : std_logic;
signal \N__59329\ : std_logic;
signal \N__59324\ : std_logic;
signal \N__59317\ : std_logic;
signal \N__59314\ : std_logic;
signal \N__59311\ : std_logic;
signal \N__59310\ : std_logic;
signal \N__59307\ : std_logic;
signal \N__59306\ : std_logic;
signal \N__59303\ : std_logic;
signal \N__59300\ : std_logic;
signal \N__59297\ : std_logic;
signal \N__59290\ : std_logic;
signal \N__59289\ : std_logic;
signal \N__59286\ : std_logic;
signal \N__59283\ : std_logic;
signal \N__59280\ : std_logic;
signal \N__59279\ : std_logic;
signal \N__59278\ : std_logic;
signal \N__59275\ : std_logic;
signal \N__59272\ : std_logic;
signal \N__59269\ : std_logic;
signal \N__59266\ : std_logic;
signal \N__59257\ : std_logic;
signal \N__59256\ : std_logic;
signal \N__59253\ : std_logic;
signal \N__59250\ : std_logic;
signal \N__59245\ : std_logic;
signal \N__59244\ : std_logic;
signal \N__59241\ : std_logic;
signal \N__59238\ : std_logic;
signal \N__59235\ : std_logic;
signal \N__59232\ : std_logic;
signal \N__59227\ : std_logic;
signal \N__59226\ : std_logic;
signal \N__59223\ : std_logic;
signal \N__59220\ : std_logic;
signal \N__59217\ : std_logic;
signal \N__59212\ : std_logic;
signal \N__59211\ : std_logic;
signal \N__59210\ : std_logic;
signal \N__59207\ : std_logic;
signal \N__59204\ : std_logic;
signal \N__59201\ : std_logic;
signal \N__59200\ : std_logic;
signal \N__59199\ : std_logic;
signal \N__59198\ : std_logic;
signal \N__59195\ : std_logic;
signal \N__59190\ : std_logic;
signal \N__59187\ : std_logic;
signal \N__59184\ : std_logic;
signal \N__59181\ : std_logic;
signal \N__59178\ : std_logic;
signal \N__59173\ : std_logic;
signal \N__59170\ : std_logic;
signal \N__59169\ : std_logic;
signal \N__59168\ : std_logic;
signal \N__59165\ : std_logic;
signal \N__59162\ : std_logic;
signal \N__59157\ : std_logic;
signal \N__59154\ : std_logic;
signal \N__59151\ : std_logic;
signal \N__59148\ : std_logic;
signal \N__59141\ : std_logic;
signal \N__59138\ : std_logic;
signal \N__59135\ : std_logic;
signal \N__59130\ : std_logic;
signal \N__59125\ : std_logic;
signal \N__59122\ : std_logic;
signal \N__59119\ : std_logic;
signal \N__59118\ : std_logic;
signal \N__59117\ : std_logic;
signal \N__59114\ : std_logic;
signal \N__59109\ : std_logic;
signal \N__59104\ : std_logic;
signal \N__59101\ : std_logic;
signal \N__59098\ : std_logic;
signal \N__59095\ : std_logic;
signal \N__59092\ : std_logic;
signal \N__59089\ : std_logic;
signal \N__59086\ : std_logic;
signal \N__59083\ : std_logic;
signal \N__59080\ : std_logic;
signal \N__59079\ : std_logic;
signal \N__59074\ : std_logic;
signal \N__59071\ : std_logic;
signal \N__59068\ : std_logic;
signal \N__59067\ : std_logic;
signal \N__59066\ : std_logic;
signal \N__59065\ : std_logic;
signal \N__59062\ : std_logic;
signal \N__59059\ : std_logic;
signal \N__59054\ : std_logic;
signal \N__59047\ : std_logic;
signal \N__59044\ : std_logic;
signal \N__59043\ : std_logic;
signal \N__59038\ : std_logic;
signal \N__59035\ : std_logic;
signal \N__59032\ : std_logic;
signal \N__59031\ : std_logic;
signal \N__59026\ : std_logic;
signal \N__59023\ : std_logic;
signal \N__59020\ : std_logic;
signal \N__59019\ : std_logic;
signal \N__59016\ : std_logic;
signal \N__59013\ : std_logic;
signal \N__59008\ : std_logic;
signal \N__59007\ : std_logic;
signal \N__59006\ : std_logic;
signal \N__59003\ : std_logic;
signal \N__59000\ : std_logic;
signal \N__58997\ : std_logic;
signal \N__58996\ : std_logic;
signal \N__58993\ : std_logic;
signal \N__58990\ : std_logic;
signal \N__58987\ : std_logic;
signal \N__58984\ : std_logic;
signal \N__58979\ : std_logic;
signal \N__58972\ : std_logic;
signal \N__58969\ : std_logic;
signal \N__58966\ : std_logic;
signal \N__58963\ : std_logic;
signal \N__58960\ : std_logic;
signal \N__58957\ : std_logic;
signal \N__58954\ : std_logic;
signal \N__58953\ : std_logic;
signal \N__58952\ : std_logic;
signal \N__58949\ : std_logic;
signal \N__58944\ : std_logic;
signal \N__58939\ : std_logic;
signal \N__58938\ : std_logic;
signal \N__58935\ : std_logic;
signal \N__58932\ : std_logic;
signal \N__58929\ : std_logic;
signal \N__58926\ : std_logic;
signal \N__58923\ : std_logic;
signal \N__58918\ : std_logic;
signal \N__58915\ : std_logic;
signal \N__58912\ : std_logic;
signal \N__58909\ : std_logic;
signal \N__58906\ : std_logic;
signal \N__58903\ : std_logic;
signal \N__58900\ : std_logic;
signal \N__58899\ : std_logic;
signal \N__58898\ : std_logic;
signal \N__58897\ : std_logic;
signal \N__58896\ : std_logic;
signal \N__58893\ : std_logic;
signal \N__58890\ : std_logic;
signal \N__58885\ : std_logic;
signal \N__58882\ : std_logic;
signal \N__58873\ : std_logic;
signal \N__58870\ : std_logic;
signal \N__58867\ : std_logic;
signal \N__58866\ : std_logic;
signal \N__58861\ : std_logic;
signal \N__58858\ : std_logic;
signal \N__58855\ : std_logic;
signal \N__58852\ : std_logic;
signal \N__58849\ : std_logic;
signal \N__58846\ : std_logic;
signal \N__58845\ : std_logic;
signal \N__58842\ : std_logic;
signal \N__58839\ : std_logic;
signal \N__58838\ : std_logic;
signal \N__58837\ : std_logic;
signal \N__58836\ : std_logic;
signal \N__58835\ : std_logic;
signal \N__58832\ : std_logic;
signal \N__58829\ : std_logic;
signal \N__58826\ : std_logic;
signal \N__58823\ : std_logic;
signal \N__58822\ : std_logic;
signal \N__58819\ : std_logic;
signal \N__58816\ : std_logic;
signal \N__58813\ : std_logic;
signal \N__58810\ : std_logic;
signal \N__58807\ : std_logic;
signal \N__58804\ : std_logic;
signal \N__58799\ : std_logic;
signal \N__58796\ : std_logic;
signal \N__58793\ : std_logic;
signal \N__58788\ : std_logic;
signal \N__58783\ : std_logic;
signal \N__58774\ : std_logic;
signal \N__58771\ : std_logic;
signal \N__58770\ : std_logic;
signal \N__58767\ : std_logic;
signal \N__58766\ : std_logic;
signal \N__58763\ : std_logic;
signal \N__58760\ : std_logic;
signal \N__58757\ : std_logic;
signal \N__58754\ : std_logic;
signal \N__58751\ : std_logic;
signal \N__58746\ : std_logic;
signal \N__58741\ : std_logic;
signal \N__58740\ : std_logic;
signal \N__58737\ : std_logic;
signal \N__58734\ : std_logic;
signal \N__58729\ : std_logic;
signal \N__58726\ : std_logic;
signal \N__58723\ : std_logic;
signal \N__58720\ : std_logic;
signal \N__58717\ : std_logic;
signal \N__58714\ : std_logic;
signal \N__58713\ : std_logic;
signal \N__58712\ : std_logic;
signal \N__58709\ : std_logic;
signal \N__58706\ : std_logic;
signal \N__58703\ : std_logic;
signal \N__58696\ : std_logic;
signal \N__58693\ : std_logic;
signal \N__58692\ : std_logic;
signal \N__58691\ : std_logic;
signal \N__58688\ : std_logic;
signal \N__58685\ : std_logic;
signal \N__58682\ : std_logic;
signal \N__58675\ : std_logic;
signal \N__58672\ : std_logic;
signal \N__58669\ : std_logic;
signal \N__58666\ : std_logic;
signal \N__58663\ : std_logic;
signal \N__58660\ : std_logic;
signal \N__58657\ : std_logic;
signal \N__58654\ : std_logic;
signal \N__58651\ : std_logic;
signal \N__58648\ : std_logic;
signal \N__58645\ : std_logic;
signal \N__58644\ : std_logic;
signal \N__58643\ : std_logic;
signal \N__58638\ : std_logic;
signal \N__58637\ : std_logic;
signal \N__58634\ : std_logic;
signal \N__58631\ : std_logic;
signal \N__58628\ : std_logic;
signal \N__58623\ : std_logic;
signal \N__58618\ : std_logic;
signal \N__58615\ : std_logic;
signal \N__58614\ : std_logic;
signal \N__58611\ : std_logic;
signal \N__58610\ : std_logic;
signal \N__58609\ : std_logic;
signal \N__58606\ : std_logic;
signal \N__58603\ : std_logic;
signal \N__58600\ : std_logic;
signal \N__58597\ : std_logic;
signal \N__58594\ : std_logic;
signal \N__58591\ : std_logic;
signal \N__58588\ : std_logic;
signal \N__58583\ : std_logic;
signal \N__58580\ : std_logic;
signal \N__58573\ : std_logic;
signal \N__58570\ : std_logic;
signal \N__58567\ : std_logic;
signal \N__58564\ : std_logic;
signal \N__58561\ : std_logic;
signal \N__58560\ : std_logic;
signal \N__58557\ : std_logic;
signal \N__58554\ : std_logic;
signal \N__58551\ : std_logic;
signal \N__58548\ : std_logic;
signal \N__58543\ : std_logic;
signal \N__58542\ : std_logic;
signal \N__58541\ : std_logic;
signal \N__58536\ : std_logic;
signal \N__58533\ : std_logic;
signal \N__58528\ : std_logic;
signal \N__58525\ : std_logic;
signal \N__58522\ : std_logic;
signal \N__58519\ : std_logic;
signal \N__58516\ : std_logic;
signal \N__58513\ : std_logic;
signal \N__58510\ : std_logic;
signal \N__58507\ : std_logic;
signal \N__58504\ : std_logic;
signal \N__58501\ : std_logic;
signal \N__58498\ : std_logic;
signal \N__58497\ : std_logic;
signal \N__58494\ : std_logic;
signal \N__58491\ : std_logic;
signal \N__58490\ : std_logic;
signal \N__58487\ : std_logic;
signal \N__58484\ : std_logic;
signal \N__58483\ : std_logic;
signal \N__58480\ : std_logic;
signal \N__58475\ : std_logic;
signal \N__58472\ : std_logic;
signal \N__58469\ : std_logic;
signal \N__58466\ : std_logic;
signal \N__58459\ : std_logic;
signal \N__58458\ : std_logic;
signal \N__58455\ : std_logic;
signal \N__58452\ : std_logic;
signal \N__58447\ : std_logic;
signal \N__58446\ : std_logic;
signal \N__58441\ : std_logic;
signal \N__58438\ : std_logic;
signal \N__58435\ : std_logic;
signal \N__58432\ : std_logic;
signal \N__58429\ : std_logic;
signal \N__58428\ : std_logic;
signal \N__58427\ : std_logic;
signal \N__58426\ : std_logic;
signal \N__58423\ : std_logic;
signal \N__58420\ : std_logic;
signal \N__58417\ : std_logic;
signal \N__58414\ : std_logic;
signal \N__58409\ : std_logic;
signal \N__58404\ : std_logic;
signal \N__58401\ : std_logic;
signal \N__58396\ : std_logic;
signal \N__58393\ : std_logic;
signal \N__58390\ : std_logic;
signal \N__58387\ : std_logic;
signal \N__58384\ : std_logic;
signal \N__58381\ : std_logic;
signal \N__58378\ : std_logic;
signal \N__58377\ : std_logic;
signal \N__58374\ : std_logic;
signal \N__58371\ : std_logic;
signal \N__58368\ : std_logic;
signal \N__58365\ : std_logic;
signal \N__58362\ : std_logic;
signal \N__58357\ : std_logic;
signal \N__58354\ : std_logic;
signal \N__58351\ : std_logic;
signal \N__58348\ : std_logic;
signal \N__58345\ : std_logic;
signal \N__58342\ : std_logic;
signal \N__58341\ : std_logic;
signal \N__58338\ : std_logic;
signal \N__58337\ : std_logic;
signal \N__58334\ : std_logic;
signal \N__58331\ : std_logic;
signal \N__58328\ : std_logic;
signal \N__58327\ : std_logic;
signal \N__58324\ : std_logic;
signal \N__58321\ : std_logic;
signal \N__58318\ : std_logic;
signal \N__58315\ : std_logic;
signal \N__58312\ : std_logic;
signal \N__58309\ : std_logic;
signal \N__58300\ : std_logic;
signal \N__58297\ : std_logic;
signal \N__58294\ : std_logic;
signal \N__58291\ : std_logic;
signal \N__58288\ : std_logic;
signal \N__58285\ : std_logic;
signal \N__58282\ : std_logic;
signal \N__58279\ : std_logic;
signal \N__58278\ : std_logic;
signal \N__58275\ : std_logic;
signal \N__58272\ : std_logic;
signal \N__58269\ : std_logic;
signal \N__58266\ : std_logic;
signal \N__58261\ : std_logic;
signal \N__58258\ : std_logic;
signal \N__58257\ : std_logic;
signal \N__58256\ : std_logic;
signal \N__58253\ : std_logic;
signal \N__58248\ : std_logic;
signal \N__58243\ : std_logic;
signal \N__58240\ : std_logic;
signal \N__58237\ : std_logic;
signal \N__58236\ : std_logic;
signal \N__58233\ : std_logic;
signal \N__58230\ : std_logic;
signal \N__58227\ : std_logic;
signal \N__58224\ : std_logic;
signal \N__58221\ : std_logic;
signal \N__58216\ : std_logic;
signal \N__58213\ : std_logic;
signal \N__58212\ : std_logic;
signal \N__58209\ : std_logic;
signal \N__58206\ : std_logic;
signal \N__58205\ : std_logic;
signal \N__58200\ : std_logic;
signal \N__58197\ : std_logic;
signal \N__58194\ : std_logic;
signal \N__58189\ : std_logic;
signal \N__58186\ : std_logic;
signal \N__58185\ : std_logic;
signal \N__58182\ : std_logic;
signal \N__58179\ : std_logic;
signal \N__58174\ : std_logic;
signal \N__58173\ : std_logic;
signal \N__58172\ : std_logic;
signal \N__58169\ : std_logic;
signal \N__58166\ : std_logic;
signal \N__58163\ : std_logic;
signal \N__58162\ : std_logic;
signal \N__58159\ : std_logic;
signal \N__58156\ : std_logic;
signal \N__58153\ : std_logic;
signal \N__58150\ : std_logic;
signal \N__58141\ : std_logic;
signal \N__58138\ : std_logic;
signal \N__58137\ : std_logic;
signal \N__58134\ : std_logic;
signal \N__58131\ : std_logic;
signal \N__58130\ : std_logic;
signal \N__58127\ : std_logic;
signal \N__58124\ : std_logic;
signal \N__58121\ : std_logic;
signal \N__58118\ : std_logic;
signal \N__58115\ : std_logic;
signal \N__58112\ : std_logic;
signal \N__58109\ : std_logic;
signal \N__58106\ : std_logic;
signal \N__58099\ : std_logic;
signal \N__58098\ : std_logic;
signal \N__58095\ : std_logic;
signal \N__58094\ : std_logic;
signal \N__58091\ : std_logic;
signal \N__58088\ : std_logic;
signal \N__58085\ : std_logic;
signal \N__58082\ : std_logic;
signal \N__58075\ : std_logic;
signal \N__58072\ : std_logic;
signal \N__58069\ : std_logic;
signal \N__58068\ : std_logic;
signal \N__58067\ : std_logic;
signal \N__58064\ : std_logic;
signal \N__58063\ : std_logic;
signal \N__58062\ : std_logic;
signal \N__58061\ : std_logic;
signal \N__58056\ : std_logic;
signal \N__58051\ : std_logic;
signal \N__58046\ : std_logic;
signal \N__58043\ : std_logic;
signal \N__58036\ : std_logic;
signal \N__58033\ : std_logic;
signal \N__58030\ : std_logic;
signal \N__58029\ : std_logic;
signal \N__58028\ : std_logic;
signal \N__58025\ : std_logic;
signal \N__58022\ : std_logic;
signal \N__58019\ : std_logic;
signal \N__58018\ : std_logic;
signal \N__58013\ : std_logic;
signal \N__58010\ : std_logic;
signal \N__58007\ : std_logic;
signal \N__58004\ : std_logic;
signal \N__57997\ : std_logic;
signal \N__57994\ : std_logic;
signal \N__57991\ : std_logic;
signal \N__57988\ : std_logic;
signal \N__57987\ : std_logic;
signal \N__57984\ : std_logic;
signal \N__57981\ : std_logic;
signal \N__57978\ : std_logic;
signal \N__57973\ : std_logic;
signal \N__57972\ : std_logic;
signal \N__57969\ : std_logic;
signal \N__57966\ : std_logic;
signal \N__57963\ : std_logic;
signal \N__57960\ : std_logic;
signal \N__57955\ : std_logic;
signal \N__57952\ : std_logic;
signal \N__57949\ : std_logic;
signal \N__57946\ : std_logic;
signal \N__57943\ : std_logic;
signal \N__57940\ : std_logic;
signal \N__57937\ : std_logic;
signal \N__57936\ : std_logic;
signal \N__57933\ : std_logic;
signal \N__57930\ : std_logic;
signal \N__57925\ : std_logic;
signal \N__57924\ : std_logic;
signal \N__57921\ : std_logic;
signal \N__57918\ : std_logic;
signal \N__57915\ : std_logic;
signal \N__57910\ : std_logic;
signal \N__57909\ : std_logic;
signal \N__57908\ : std_logic;
signal \N__57905\ : std_logic;
signal \N__57902\ : std_logic;
signal \N__57899\ : std_logic;
signal \N__57896\ : std_logic;
signal \N__57893\ : std_logic;
signal \N__57890\ : std_logic;
signal \N__57889\ : std_logic;
signal \N__57882\ : std_logic;
signal \N__57879\ : std_logic;
signal \N__57874\ : std_logic;
signal \N__57871\ : std_logic;
signal \N__57870\ : std_logic;
signal \N__57869\ : std_logic;
signal \N__57866\ : std_logic;
signal \N__57863\ : std_logic;
signal \N__57860\ : std_logic;
signal \N__57857\ : std_logic;
signal \N__57850\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57844\ : std_logic;
signal \N__57843\ : std_logic;
signal \N__57842\ : std_logic;
signal \N__57839\ : std_logic;
signal \N__57834\ : std_logic;
signal \N__57829\ : std_logic;
signal \N__57826\ : std_logic;
signal \N__57823\ : std_logic;
signal \N__57820\ : std_logic;
signal \N__57817\ : std_logic;
signal \N__57814\ : std_logic;
signal \N__57811\ : std_logic;
signal \N__57810\ : std_logic;
signal \N__57809\ : std_logic;
signal \N__57806\ : std_logic;
signal \N__57801\ : std_logic;
signal \N__57796\ : std_logic;
signal \N__57795\ : std_logic;
signal \N__57792\ : std_logic;
signal \N__57789\ : std_logic;
signal \N__57786\ : std_logic;
signal \N__57783\ : std_logic;
signal \N__57778\ : std_logic;
signal \N__57775\ : std_logic;
signal \N__57772\ : std_logic;
signal \N__57769\ : std_logic;
signal \N__57766\ : std_logic;
signal \N__57763\ : std_logic;
signal \N__57760\ : std_logic;
signal \N__57757\ : std_logic;
signal \N__57756\ : std_logic;
signal \N__57753\ : std_logic;
signal \N__57750\ : std_logic;
signal \N__57747\ : std_logic;
signal \N__57742\ : std_logic;
signal \N__57739\ : std_logic;
signal \N__57736\ : std_logic;
signal \N__57733\ : std_logic;
signal \N__57732\ : std_logic;
signal \N__57731\ : std_logic;
signal \N__57730\ : std_logic;
signal \N__57727\ : std_logic;
signal \N__57724\ : std_logic;
signal \N__57721\ : std_logic;
signal \N__57718\ : std_logic;
signal \N__57713\ : std_logic;
signal \N__57712\ : std_logic;
signal \N__57709\ : std_logic;
signal \N__57706\ : std_logic;
signal \N__57703\ : std_logic;
signal \N__57700\ : std_logic;
signal \N__57691\ : std_logic;
signal \N__57688\ : std_logic;
signal \N__57685\ : std_logic;
signal \N__57682\ : std_logic;
signal \N__57679\ : std_logic;
signal \N__57676\ : std_logic;
signal \N__57675\ : std_logic;
signal \N__57674\ : std_logic;
signal \N__57671\ : std_logic;
signal \N__57668\ : std_logic;
signal \N__57665\ : std_logic;
signal \N__57658\ : std_logic;
signal \N__57655\ : std_logic;
signal \N__57652\ : std_logic;
signal \N__57649\ : std_logic;
signal \N__57646\ : std_logic;
signal \N__57643\ : std_logic;
signal \N__57640\ : std_logic;
signal \N__57639\ : std_logic;
signal \N__57636\ : std_logic;
signal \N__57633\ : std_logic;
signal \N__57632\ : std_logic;
signal \N__57629\ : std_logic;
signal \N__57624\ : std_logic;
signal \N__57619\ : std_logic;
signal \N__57616\ : std_logic;
signal \N__57615\ : std_logic;
signal \N__57614\ : std_logic;
signal \N__57609\ : std_logic;
signal \N__57606\ : std_logic;
signal \N__57605\ : std_logic;
signal \N__57602\ : std_logic;
signal \N__57597\ : std_logic;
signal \N__57592\ : std_logic;
signal \N__57589\ : std_logic;
signal \N__57586\ : std_logic;
signal \N__57585\ : std_logic;
signal \N__57584\ : std_logic;
signal \N__57583\ : std_logic;
signal \N__57582\ : std_logic;
signal \N__57581\ : std_logic;
signal \N__57578\ : std_logic;
signal \N__57573\ : std_logic;
signal \N__57570\ : std_logic;
signal \N__57567\ : std_logic;
signal \N__57564\ : std_logic;
signal \N__57553\ : std_logic;
signal \N__57550\ : std_logic;
signal \N__57547\ : std_logic;
signal \N__57544\ : std_logic;
signal \N__57541\ : std_logic;
signal \N__57540\ : std_logic;
signal \N__57537\ : std_logic;
signal \N__57534\ : std_logic;
signal \N__57529\ : std_logic;
signal \N__57526\ : std_logic;
signal \N__57523\ : std_logic;
signal \N__57520\ : std_logic;
signal \N__57517\ : std_logic;
signal \N__57514\ : std_logic;
signal \N__57511\ : std_logic;
signal \N__57508\ : std_logic;
signal \N__57505\ : std_logic;
signal \N__57502\ : std_logic;
signal \N__57499\ : std_logic;
signal \N__57498\ : std_logic;
signal \N__57493\ : std_logic;
signal \N__57490\ : std_logic;
signal \N__57489\ : std_logic;
signal \N__57486\ : std_logic;
signal \N__57483\ : std_logic;
signal \N__57480\ : std_logic;
signal \N__57477\ : std_logic;
signal \N__57472\ : std_logic;
signal \N__57469\ : std_logic;
signal \N__57468\ : std_logic;
signal \N__57465\ : std_logic;
signal \N__57462\ : std_logic;
signal \N__57459\ : std_logic;
signal \N__57456\ : std_logic;
signal \N__57451\ : std_logic;
signal \N__57448\ : std_logic;
signal \N__57447\ : std_logic;
signal \N__57446\ : std_logic;
signal \N__57445\ : std_logic;
signal \N__57444\ : std_logic;
signal \N__57441\ : std_logic;
signal \N__57438\ : std_logic;
signal \N__57433\ : std_logic;
signal \N__57430\ : std_logic;
signal \N__57425\ : std_logic;
signal \N__57422\ : std_logic;
signal \N__57419\ : std_logic;
signal \N__57416\ : std_logic;
signal \N__57413\ : std_logic;
signal \N__57406\ : std_logic;
signal \N__57403\ : std_logic;
signal \N__57400\ : std_logic;
signal \N__57397\ : std_logic;
signal \N__57396\ : std_logic;
signal \N__57395\ : std_logic;
signal \N__57392\ : std_logic;
signal \N__57387\ : std_logic;
signal \N__57382\ : std_logic;
signal \N__57379\ : std_logic;
signal \N__57376\ : std_logic;
signal \N__57373\ : std_logic;
signal \N__57370\ : std_logic;
signal \N__57369\ : std_logic;
signal \N__57366\ : std_logic;
signal \N__57365\ : std_logic;
signal \N__57362\ : std_logic;
signal \N__57359\ : std_logic;
signal \N__57356\ : std_logic;
signal \N__57353\ : std_logic;
signal \N__57346\ : std_logic;
signal \N__57345\ : std_logic;
signal \N__57342\ : std_logic;
signal \N__57339\ : std_logic;
signal \N__57336\ : std_logic;
signal \N__57333\ : std_logic;
signal \N__57330\ : std_logic;
signal \N__57325\ : std_logic;
signal \N__57324\ : std_logic;
signal \N__57321\ : std_logic;
signal \N__57318\ : std_logic;
signal \N__57315\ : std_logic;
signal \N__57314\ : std_logic;
signal \N__57313\ : std_logic;
signal \N__57310\ : std_logic;
signal \N__57307\ : std_logic;
signal \N__57304\ : std_logic;
signal \N__57301\ : std_logic;
signal \N__57292\ : std_logic;
signal \N__57291\ : std_logic;
signal \N__57286\ : std_logic;
signal \N__57285\ : std_logic;
signal \N__57284\ : std_logic;
signal \N__57283\ : std_logic;
signal \N__57280\ : std_logic;
signal \N__57277\ : std_logic;
signal \N__57274\ : std_logic;
signal \N__57271\ : std_logic;
signal \N__57266\ : std_logic;
signal \N__57263\ : std_logic;
signal \N__57258\ : std_logic;
signal \N__57253\ : std_logic;
signal \N__57250\ : std_logic;
signal \N__57247\ : std_logic;
signal \N__57244\ : std_logic;
signal \N__57241\ : std_logic;
signal \N__57238\ : std_logic;
signal \N__57235\ : std_logic;
signal \N__57234\ : std_logic;
signal \N__57231\ : std_logic;
signal \N__57228\ : std_logic;
signal \N__57225\ : std_logic;
signal \N__57220\ : std_logic;
signal \N__57217\ : std_logic;
signal \N__57216\ : std_logic;
signal \N__57213\ : std_logic;
signal \N__57210\ : std_logic;
signal \N__57207\ : std_logic;
signal \N__57204\ : std_logic;
signal \N__57199\ : std_logic;
signal \N__57196\ : std_logic;
signal \N__57193\ : std_logic;
signal \N__57190\ : std_logic;
signal \N__57187\ : std_logic;
signal \N__57186\ : std_logic;
signal \N__57183\ : std_logic;
signal \N__57178\ : std_logic;
signal \N__57175\ : std_logic;
signal \N__57172\ : std_logic;
signal \N__57169\ : std_logic;
signal \N__57166\ : std_logic;
signal \N__57163\ : std_logic;
signal \N__57160\ : std_logic;
signal \N__57159\ : std_logic;
signal \N__57158\ : std_logic;
signal \N__57157\ : std_logic;
signal \N__57156\ : std_logic;
signal \N__57155\ : std_logic;
signal \N__57154\ : std_logic;
signal \N__57151\ : std_logic;
signal \N__57146\ : std_logic;
signal \N__57143\ : std_logic;
signal \N__57136\ : std_logic;
signal \N__57127\ : std_logic;
signal \N__57126\ : std_logic;
signal \N__57123\ : std_logic;
signal \N__57120\ : std_logic;
signal \N__57115\ : std_logic;
signal \N__57112\ : std_logic;
signal \N__57109\ : std_logic;
signal \N__57106\ : std_logic;
signal \N__57105\ : std_logic;
signal \N__57102\ : std_logic;
signal \N__57101\ : std_logic;
signal \N__57098\ : std_logic;
signal \N__57095\ : std_logic;
signal \N__57092\ : std_logic;
signal \N__57091\ : std_logic;
signal \N__57090\ : std_logic;
signal \N__57085\ : std_logic;
signal \N__57082\ : std_logic;
signal \N__57079\ : std_logic;
signal \N__57076\ : std_logic;
signal \N__57073\ : std_logic;
signal \N__57064\ : std_logic;
signal \N__57061\ : std_logic;
signal \N__57060\ : std_logic;
signal \N__57059\ : std_logic;
signal \N__57058\ : std_logic;
signal \N__57055\ : std_logic;
signal \N__57054\ : std_logic;
signal \N__57051\ : std_logic;
signal \N__57048\ : std_logic;
signal \N__57045\ : std_logic;
signal \N__57042\ : std_logic;
signal \N__57039\ : std_logic;
signal \N__57028\ : std_logic;
signal \N__57027\ : std_logic;
signal \N__57024\ : std_logic;
signal \N__57021\ : std_logic;
signal \N__57018\ : std_logic;
signal \N__57015\ : std_logic;
signal \N__57012\ : std_logic;
signal \N__57009\ : std_logic;
signal \N__57008\ : std_logic;
signal \N__57007\ : std_logic;
signal \N__57004\ : std_logic;
signal \N__57003\ : std_logic;
signal \N__57002\ : std_logic;
signal \N__56999\ : std_logic;
signal \N__56994\ : std_logic;
signal \N__56993\ : std_logic;
signal \N__56992\ : std_logic;
signal \N__56991\ : std_logic;
signal \N__56988\ : std_logic;
signal \N__56985\ : std_logic;
signal \N__56982\ : std_logic;
signal \N__56979\ : std_logic;
signal \N__56976\ : std_logic;
signal \N__56973\ : std_logic;
signal \N__56970\ : std_logic;
signal \N__56967\ : std_logic;
signal \N__56950\ : std_logic;
signal \N__56947\ : std_logic;
signal \N__56946\ : std_logic;
signal \N__56943\ : std_logic;
signal \N__56940\ : std_logic;
signal \N__56939\ : std_logic;
signal \N__56938\ : std_logic;
signal \N__56935\ : std_logic;
signal \N__56934\ : std_logic;
signal \N__56929\ : std_logic;
signal \N__56928\ : std_logic;
signal \N__56927\ : std_logic;
signal \N__56924\ : std_logic;
signal \N__56921\ : std_logic;
signal \N__56918\ : std_logic;
signal \N__56915\ : std_logic;
signal \N__56914\ : std_logic;
signal \N__56911\ : std_logic;
signal \N__56910\ : std_logic;
signal \N__56905\ : std_logic;
signal \N__56902\ : std_logic;
signal \N__56899\ : std_logic;
signal \N__56898\ : std_logic;
signal \N__56895\ : std_logic;
signal \N__56890\ : std_logic;
signal \N__56889\ : std_logic;
signal \N__56886\ : std_logic;
signal \N__56883\ : std_logic;
signal \N__56878\ : std_logic;
signal \N__56875\ : std_logic;
signal \N__56870\ : std_logic;
signal \N__56867\ : std_logic;
signal \N__56864\ : std_logic;
signal \N__56861\ : std_logic;
signal \N__56858\ : std_logic;
signal \N__56845\ : std_logic;
signal \N__56842\ : std_logic;
signal \N__56839\ : std_logic;
signal \N__56836\ : std_logic;
signal \N__56835\ : std_logic;
signal \N__56832\ : std_logic;
signal \N__56829\ : std_logic;
signal \N__56828\ : std_logic;
signal \N__56827\ : std_logic;
signal \N__56826\ : std_logic;
signal \N__56823\ : std_logic;
signal \N__56822\ : std_logic;
signal \N__56819\ : std_logic;
signal \N__56818\ : std_logic;
signal \N__56811\ : std_logic;
signal \N__56810\ : std_logic;
signal \N__56809\ : std_logic;
signal \N__56808\ : std_logic;
signal \N__56805\ : std_logic;
signal \N__56802\ : std_logic;
signal \N__56799\ : std_logic;
signal \N__56796\ : std_logic;
signal \N__56793\ : std_logic;
signal \N__56788\ : std_logic;
signal \N__56785\ : std_logic;
signal \N__56770\ : std_logic;
signal \N__56767\ : std_logic;
signal \N__56764\ : std_logic;
signal \N__56763\ : std_logic;
signal \N__56760\ : std_logic;
signal \N__56757\ : std_logic;
signal \N__56754\ : std_logic;
signal \N__56749\ : std_logic;
signal \N__56748\ : std_logic;
signal \N__56745\ : std_logic;
signal \N__56744\ : std_logic;
signal \N__56743\ : std_logic;
signal \N__56742\ : std_logic;
signal \N__56739\ : std_logic;
signal \N__56736\ : std_logic;
signal \N__56733\ : std_logic;
signal \N__56730\ : std_logic;
signal \N__56729\ : std_logic;
signal \N__56726\ : std_logic;
signal \N__56723\ : std_logic;
signal \N__56720\ : std_logic;
signal \N__56719\ : std_logic;
signal \N__56718\ : std_logic;
signal \N__56715\ : std_logic;
signal \N__56712\ : std_logic;
signal \N__56709\ : std_logic;
signal \N__56708\ : std_logic;
signal \N__56705\ : std_logic;
signal \N__56700\ : std_logic;
signal \N__56699\ : std_logic;
signal \N__56696\ : std_logic;
signal \N__56693\ : std_logic;
signal \N__56692\ : std_logic;
signal \N__56691\ : std_logic;
signal \N__56688\ : std_logic;
signal \N__56683\ : std_logic;
signal \N__56680\ : std_logic;
signal \N__56675\ : std_logic;
signal \N__56672\ : std_logic;
signal \N__56669\ : std_logic;
signal \N__56666\ : std_logic;
signal \N__56661\ : std_logic;
signal \N__56658\ : std_logic;
signal \N__56653\ : std_logic;
signal \N__56648\ : std_logic;
signal \N__56645\ : std_logic;
signal \N__56642\ : std_logic;
signal \N__56639\ : std_logic;
signal \N__56636\ : std_logic;
signal \N__56631\ : std_logic;
signal \N__56630\ : std_logic;
signal \N__56625\ : std_logic;
signal \N__56620\ : std_logic;
signal \N__56617\ : std_logic;
signal \N__56614\ : std_logic;
signal \N__56605\ : std_logic;
signal \N__56602\ : std_logic;
signal \N__56601\ : std_logic;
signal \N__56600\ : std_logic;
signal \N__56599\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56597\ : std_logic;
signal \N__56596\ : std_logic;
signal \N__56593\ : std_logic;
signal \N__56590\ : std_logic;
signal \N__56589\ : std_logic;
signal \N__56586\ : std_logic;
signal \N__56583\ : std_logic;
signal \N__56582\ : std_logic;
signal \N__56579\ : std_logic;
signal \N__56574\ : std_logic;
signal \N__56573\ : std_logic;
signal \N__56570\ : std_logic;
signal \N__56569\ : std_logic;
signal \N__56568\ : std_logic;
signal \N__56565\ : std_logic;
signal \N__56562\ : std_logic;
signal \N__56557\ : std_logic;
signal \N__56554\ : std_logic;
signal \N__56551\ : std_logic;
signal \N__56548\ : std_logic;
signal \N__56545\ : std_logic;
signal \N__56544\ : std_logic;
signal \N__56541\ : std_logic;
signal \N__56538\ : std_logic;
signal \N__56535\ : std_logic;
signal \N__56530\ : std_logic;
signal \N__56527\ : std_logic;
signal \N__56520\ : std_logic;
signal \N__56517\ : std_logic;
signal \N__56514\ : std_logic;
signal \N__56507\ : std_logic;
signal \N__56504\ : std_logic;
signal \N__56501\ : std_logic;
signal \N__56496\ : std_logic;
signal \N__56495\ : std_logic;
signal \N__56492\ : std_logic;
signal \N__56487\ : std_logic;
signal \N__56484\ : std_logic;
signal \N__56481\ : std_logic;
signal \N__56478\ : std_logic;
signal \N__56467\ : std_logic;
signal \N__56466\ : std_logic;
signal \N__56465\ : std_logic;
signal \N__56462\ : std_logic;
signal \N__56459\ : std_logic;
signal \N__56458\ : std_logic;
signal \N__56457\ : std_logic;
signal \N__56456\ : std_logic;
signal \N__56455\ : std_logic;
signal \N__56452\ : std_logic;
signal \N__56449\ : std_logic;
signal \N__56446\ : std_logic;
signal \N__56443\ : std_logic;
signal \N__56440\ : std_logic;
signal \N__56439\ : std_logic;
signal \N__56436\ : std_logic;
signal \N__56435\ : std_logic;
signal \N__56434\ : std_logic;
signal \N__56431\ : std_logic;
signal \N__56428\ : std_logic;
signal \N__56423\ : std_logic;
signal \N__56420\ : std_logic;
signal \N__56419\ : std_logic;
signal \N__56416\ : std_logic;
signal \N__56413\ : std_logic;
signal \N__56410\ : std_logic;
signal \N__56407\ : std_logic;
signal \N__56404\ : std_logic;
signal \N__56403\ : std_logic;
signal \N__56400\ : std_logic;
signal \N__56395\ : std_logic;
signal \N__56394\ : std_logic;
signal \N__56391\ : std_logic;
signal \N__56388\ : std_logic;
signal \N__56383\ : std_logic;
signal \N__56376\ : std_logic;
signal \N__56373\ : std_logic;
signal \N__56370\ : std_logic;
signal \N__56367\ : std_logic;
signal \N__56364\ : std_logic;
signal \N__56357\ : std_logic;
signal \N__56354\ : std_logic;
signal \N__56353\ : std_logic;
signal \N__56350\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56338\ : std_logic;
signal \N__56335\ : std_logic;
signal \N__56326\ : std_logic;
signal \N__56323\ : std_logic;
signal \N__56322\ : std_logic;
signal \N__56319\ : std_logic;
signal \N__56316\ : std_logic;
signal \N__56311\ : std_logic;
signal \N__56308\ : std_logic;
signal \N__56305\ : std_logic;
signal \N__56304\ : std_logic;
signal \N__56301\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56293\ : std_logic;
signal \N__56290\ : std_logic;
signal \N__56287\ : std_logic;
signal \N__56284\ : std_logic;
signal \N__56283\ : std_logic;
signal \N__56280\ : std_logic;
signal \N__56279\ : std_logic;
signal \N__56278\ : std_logic;
signal \N__56275\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56269\ : std_logic;
signal \N__56266\ : std_logic;
signal \N__56263\ : std_logic;
signal \N__56258\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56248\ : std_logic;
signal \N__56245\ : std_logic;
signal \N__56242\ : std_logic;
signal \N__56239\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56230\ : std_logic;
signal \N__56227\ : std_logic;
signal \N__56224\ : std_logic;
signal \N__56221\ : std_logic;
signal \N__56220\ : std_logic;
signal \N__56217\ : std_logic;
signal \N__56214\ : std_logic;
signal \N__56211\ : std_logic;
signal \N__56208\ : std_logic;
signal \N__56207\ : std_logic;
signal \N__56204\ : std_logic;
signal \N__56201\ : std_logic;
signal \N__56198\ : std_logic;
signal \N__56195\ : std_logic;
signal \N__56188\ : std_logic;
signal \N__56187\ : std_logic;
signal \N__56186\ : std_logic;
signal \N__56181\ : std_logic;
signal \N__56178\ : std_logic;
signal \N__56175\ : std_logic;
signal \N__56172\ : std_logic;
signal \N__56169\ : std_logic;
signal \N__56164\ : std_logic;
signal \N__56161\ : std_logic;
signal \N__56160\ : std_logic;
signal \N__56157\ : std_logic;
signal \N__56154\ : std_logic;
signal \N__56149\ : std_logic;
signal \N__56146\ : std_logic;
signal \N__56143\ : std_logic;
signal \N__56142\ : std_logic;
signal \N__56139\ : std_logic;
signal \N__56138\ : std_logic;
signal \N__56135\ : std_logic;
signal \N__56132\ : std_logic;
signal \N__56129\ : std_logic;
signal \N__56126\ : std_logic;
signal \N__56123\ : std_logic;
signal \N__56120\ : std_logic;
signal \N__56117\ : std_logic;
signal \N__56114\ : std_logic;
signal \N__56107\ : std_logic;
signal \N__56104\ : std_logic;
signal \N__56101\ : std_logic;
signal \N__56098\ : std_logic;
signal \N__56095\ : std_logic;
signal \N__56092\ : std_logic;
signal \N__56089\ : std_logic;
signal \N__56086\ : std_logic;
signal \N__56083\ : std_logic;
signal \N__56080\ : std_logic;
signal \N__56077\ : std_logic;
signal \N__56074\ : std_logic;
signal \N__56071\ : std_logic;
signal \N__56068\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56062\ : std_logic;
signal \N__56059\ : std_logic;
signal \N__56058\ : std_logic;
signal \N__56057\ : std_logic;
signal \N__56054\ : std_logic;
signal \N__56053\ : std_logic;
signal \N__56050\ : std_logic;
signal \N__56047\ : std_logic;
signal \N__56044\ : std_logic;
signal \N__56041\ : std_logic;
signal \N__56038\ : std_logic;
signal \N__56035\ : std_logic;
signal \N__56032\ : std_logic;
signal \N__56029\ : std_logic;
signal \N__56020\ : std_logic;
signal \N__56017\ : std_logic;
signal \N__56014\ : std_logic;
signal \N__56011\ : std_logic;
signal \N__56010\ : std_logic;
signal \N__56007\ : std_logic;
signal \N__56006\ : std_logic;
signal \N__56003\ : std_logic;
signal \N__56000\ : std_logic;
signal \N__55999\ : std_logic;
signal \N__55996\ : std_logic;
signal \N__55993\ : std_logic;
signal \N__55990\ : std_logic;
signal \N__55987\ : std_logic;
signal \N__55984\ : std_logic;
signal \N__55981\ : std_logic;
signal \N__55978\ : std_logic;
signal \N__55975\ : std_logic;
signal \N__55966\ : std_logic;
signal \N__55965\ : std_logic;
signal \N__55964\ : std_logic;
signal \N__55959\ : std_logic;
signal \N__55956\ : std_logic;
signal \N__55953\ : std_logic;
signal \N__55948\ : std_logic;
signal \N__55945\ : std_logic;
signal \N__55942\ : std_logic;
signal \N__55939\ : std_logic;
signal \N__55938\ : std_logic;
signal \N__55935\ : std_logic;
signal \N__55932\ : std_logic;
signal \N__55929\ : std_logic;
signal \N__55924\ : std_logic;
signal \N__55921\ : std_logic;
signal \N__55920\ : std_logic;
signal \N__55919\ : std_logic;
signal \N__55916\ : std_logic;
signal \N__55911\ : std_logic;
signal \N__55908\ : std_logic;
signal \N__55905\ : std_logic;
signal \N__55900\ : std_logic;
signal \N__55897\ : std_logic;
signal \N__55896\ : std_logic;
signal \N__55895\ : std_logic;
signal \N__55894\ : std_logic;
signal \N__55891\ : std_logic;
signal \N__55890\ : std_logic;
signal \N__55887\ : std_logic;
signal \N__55884\ : std_logic;
signal \N__55877\ : std_logic;
signal \N__55876\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55870\ : std_logic;
signal \N__55867\ : std_logic;
signal \N__55864\ : std_logic;
signal \N__55861\ : std_logic;
signal \N__55858\ : std_logic;
signal \N__55855\ : std_logic;
signal \N__55846\ : std_logic;
signal \N__55843\ : std_logic;
signal \N__55840\ : std_logic;
signal \N__55839\ : std_logic;
signal \N__55836\ : std_logic;
signal \N__55833\ : std_logic;
signal \N__55830\ : std_logic;
signal \N__55829\ : std_logic;
signal \N__55826\ : std_logic;
signal \N__55823\ : std_logic;
signal \N__55820\ : std_logic;
signal \N__55815\ : std_logic;
signal \N__55810\ : std_logic;
signal \N__55807\ : std_logic;
signal \N__55804\ : std_logic;
signal \N__55801\ : std_logic;
signal \N__55798\ : std_logic;
signal \N__55795\ : std_logic;
signal \N__55794\ : std_logic;
signal \N__55791\ : std_logic;
signal \N__55788\ : std_logic;
signal \N__55783\ : std_logic;
signal \N__55780\ : std_logic;
signal \N__55777\ : std_logic;
signal \N__55774\ : std_logic;
signal \N__55771\ : std_logic;
signal \N__55768\ : std_logic;
signal \N__55765\ : std_logic;
signal \N__55762\ : std_logic;
signal \N__55759\ : std_logic;
signal \N__55756\ : std_logic;
signal \N__55753\ : std_logic;
signal \N__55750\ : std_logic;
signal \N__55749\ : std_logic;
signal \N__55746\ : std_logic;
signal \N__55743\ : std_logic;
signal \N__55738\ : std_logic;
signal \N__55735\ : std_logic;
signal \N__55732\ : std_logic;
signal \N__55729\ : std_logic;
signal \N__55728\ : std_logic;
signal \N__55725\ : std_logic;
signal \N__55724\ : std_logic;
signal \N__55721\ : std_logic;
signal \N__55718\ : std_logic;
signal \N__55715\ : std_logic;
signal \N__55712\ : std_logic;
signal \N__55709\ : std_logic;
signal \N__55706\ : std_logic;
signal \N__55703\ : std_logic;
signal \N__55700\ : std_logic;
signal \N__55697\ : std_logic;
signal \N__55690\ : std_logic;
signal \N__55687\ : std_logic;
signal \N__55684\ : std_logic;
signal \N__55681\ : std_logic;
signal \N__55678\ : std_logic;
signal \N__55675\ : std_logic;
signal \N__55672\ : std_logic;
signal \N__55669\ : std_logic;
signal \N__55668\ : std_logic;
signal \N__55665\ : std_logic;
signal \N__55662\ : std_logic;
signal \N__55659\ : std_logic;
signal \N__55656\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55645\ : std_logic;
signal \N__55642\ : std_logic;
signal \N__55641\ : std_logic;
signal \N__55638\ : std_logic;
signal \N__55635\ : std_logic;
signal \N__55630\ : std_logic;
signal \N__55627\ : std_logic;
signal \N__55626\ : std_logic;
signal \N__55625\ : std_logic;
signal \N__55624\ : std_logic;
signal \N__55623\ : std_logic;
signal \N__55620\ : std_logic;
signal \N__55617\ : std_logic;
signal \N__55614\ : std_logic;
signal \N__55609\ : std_logic;
signal \N__55606\ : std_logic;
signal \N__55603\ : std_logic;
signal \N__55600\ : std_logic;
signal \N__55597\ : std_logic;
signal \N__55594\ : std_logic;
signal \N__55591\ : std_logic;
signal \N__55588\ : std_logic;
signal \N__55585\ : std_logic;
signal \N__55576\ : std_logic;
signal \N__55573\ : std_logic;
signal \N__55570\ : std_logic;
signal \N__55567\ : std_logic;
signal \N__55564\ : std_logic;
signal \N__55563\ : std_logic;
signal \N__55558\ : std_logic;
signal \N__55557\ : std_logic;
signal \N__55554\ : std_logic;
signal \N__55551\ : std_logic;
signal \N__55548\ : std_logic;
signal \N__55543\ : std_logic;
signal \N__55540\ : std_logic;
signal \N__55539\ : std_logic;
signal \N__55536\ : std_logic;
signal \N__55535\ : std_logic;
signal \N__55534\ : std_logic;
signal \N__55531\ : std_logic;
signal \N__55528\ : std_logic;
signal \N__55525\ : std_logic;
signal \N__55522\ : std_logic;
signal \N__55513\ : std_logic;
signal \N__55510\ : std_logic;
signal \N__55509\ : std_logic;
signal \N__55506\ : std_logic;
signal \N__55503\ : std_logic;
signal \N__55498\ : std_logic;
signal \N__55497\ : std_logic;
signal \N__55494\ : std_logic;
signal \N__55491\ : std_logic;
signal \N__55486\ : std_logic;
signal \N__55485\ : std_logic;
signal \N__55482\ : std_logic;
signal \N__55479\ : std_logic;
signal \N__55476\ : std_logic;
signal \N__55471\ : std_logic;
signal \N__55468\ : std_logic;
signal \N__55465\ : std_logic;
signal \N__55462\ : std_logic;
signal \N__55459\ : std_logic;
signal \N__55456\ : std_logic;
signal \N__55453\ : std_logic;
signal \N__55450\ : std_logic;
signal \N__55447\ : std_logic;
signal \N__55444\ : std_logic;
signal \N__55441\ : std_logic;
signal \N__55438\ : std_logic;
signal \N__55435\ : std_logic;
signal \N__55432\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55429\ : std_logic;
signal \N__55426\ : std_logic;
signal \N__55421\ : std_logic;
signal \N__55418\ : std_logic;
signal \N__55417\ : std_logic;
signal \N__55412\ : std_logic;
signal \N__55409\ : std_logic;
signal \N__55406\ : std_logic;
signal \N__55403\ : std_logic;
signal \N__55396\ : std_logic;
signal \N__55395\ : std_logic;
signal \N__55394\ : std_logic;
signal \N__55389\ : std_logic;
signal \N__55386\ : std_logic;
signal \N__55385\ : std_logic;
signal \N__55382\ : std_logic;
signal \N__55379\ : std_logic;
signal \N__55376\ : std_logic;
signal \N__55375\ : std_logic;
signal \N__55372\ : std_logic;
signal \N__55367\ : std_logic;
signal \N__55364\ : std_logic;
signal \N__55361\ : std_logic;
signal \N__55358\ : std_logic;
signal \N__55351\ : std_logic;
signal \N__55350\ : std_logic;
signal \N__55345\ : std_logic;
signal \N__55342\ : std_logic;
signal \N__55339\ : std_logic;
signal \N__55338\ : std_logic;
signal \N__55335\ : std_logic;
signal \N__55332\ : std_logic;
signal \N__55329\ : std_logic;
signal \N__55328\ : std_logic;
signal \N__55327\ : std_logic;
signal \N__55326\ : std_logic;
signal \N__55323\ : std_logic;
signal \N__55320\ : std_logic;
signal \N__55317\ : std_logic;
signal \N__55312\ : std_logic;
signal \N__55303\ : std_logic;
signal \N__55302\ : std_logic;
signal \N__55299\ : std_logic;
signal \N__55296\ : std_logic;
signal \N__55293\ : std_logic;
signal \N__55290\ : std_logic;
signal \N__55287\ : std_logic;
signal \N__55282\ : std_logic;
signal \N__55279\ : std_logic;
signal \N__55276\ : std_logic;
signal \N__55273\ : std_logic;
signal \N__55270\ : std_logic;
signal \N__55267\ : std_logic;
signal \N__55264\ : std_logic;
signal \N__55261\ : std_logic;
signal \N__55258\ : std_logic;
signal \N__55255\ : std_logic;
signal \N__55252\ : std_logic;
signal \N__55249\ : std_logic;
signal \N__55246\ : std_logic;
signal \N__55243\ : std_logic;
signal \N__55240\ : std_logic;
signal \N__55237\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55231\ : std_logic;
signal \N__55228\ : std_logic;
signal \N__55225\ : std_logic;
signal \N__55222\ : std_logic;
signal \N__55219\ : std_logic;
signal \N__55218\ : std_logic;
signal \N__55217\ : std_logic;
signal \N__55214\ : std_logic;
signal \N__55211\ : std_logic;
signal \N__55210\ : std_logic;
signal \N__55207\ : std_logic;
signal \N__55204\ : std_logic;
signal \N__55201\ : std_logic;
signal \N__55198\ : std_logic;
signal \N__55195\ : std_logic;
signal \N__55192\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55177\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55171\ : std_logic;
signal \N__55168\ : std_logic;
signal \N__55165\ : std_logic;
signal \N__55162\ : std_logic;
signal \N__55159\ : std_logic;
signal \N__55156\ : std_logic;
signal \N__55155\ : std_logic;
signal \N__55152\ : std_logic;
signal \N__55149\ : std_logic;
signal \N__55144\ : std_logic;
signal \N__55141\ : std_logic;
signal \N__55138\ : std_logic;
signal \N__55137\ : std_logic;
signal \N__55134\ : std_logic;
signal \N__55131\ : std_logic;
signal \N__55126\ : std_logic;
signal \N__55123\ : std_logic;
signal \N__55120\ : std_logic;
signal \N__55119\ : std_logic;
signal \N__55118\ : std_logic;
signal \N__55115\ : std_logic;
signal \N__55112\ : std_logic;
signal \N__55109\ : std_logic;
signal \N__55102\ : std_logic;
signal \N__55101\ : std_logic;
signal \N__55098\ : std_logic;
signal \N__55097\ : std_logic;
signal \N__55096\ : std_logic;
signal \N__55095\ : std_logic;
signal \N__55092\ : std_logic;
signal \N__55089\ : std_logic;
signal \N__55084\ : std_logic;
signal \N__55081\ : std_logic;
signal \N__55078\ : std_logic;
signal \N__55073\ : std_logic;
signal \N__55066\ : std_logic;
signal \N__55065\ : std_logic;
signal \N__55064\ : std_logic;
signal \N__55061\ : std_logic;
signal \N__55058\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55054\ : std_logic;
signal \N__55051\ : std_logic;
signal \N__55048\ : std_logic;
signal \N__55047\ : std_logic;
signal \N__55044\ : std_logic;
signal \N__55037\ : std_logic;
signal \N__55034\ : std_logic;
signal \N__55027\ : std_logic;
signal \N__55024\ : std_logic;
signal \N__55021\ : std_logic;
signal \N__55018\ : std_logic;
signal \N__55015\ : std_logic;
signal \N__55012\ : std_logic;
signal \N__55011\ : std_logic;
signal \N__55008\ : std_logic;
signal \N__55005\ : std_logic;
signal \N__55000\ : std_logic;
signal \N__54999\ : std_logic;
signal \N__54996\ : std_logic;
signal \N__54993\ : std_logic;
signal \N__54988\ : std_logic;
signal \N__54985\ : std_logic;
signal \N__54982\ : std_logic;
signal \N__54979\ : std_logic;
signal \N__54976\ : std_logic;
signal \N__54973\ : std_logic;
signal \N__54970\ : std_logic;
signal \N__54967\ : std_logic;
signal \N__54964\ : std_logic;
signal \N__54961\ : std_logic;
signal \N__54958\ : std_logic;
signal \N__54955\ : std_logic;
signal \N__54952\ : std_logic;
signal \N__54951\ : std_logic;
signal \N__54948\ : std_logic;
signal \N__54945\ : std_logic;
signal \N__54942\ : std_logic;
signal \N__54937\ : std_logic;
signal \N__54936\ : std_logic;
signal \N__54931\ : std_logic;
signal \N__54928\ : std_logic;
signal \N__54927\ : std_logic;
signal \N__54924\ : std_logic;
signal \N__54921\ : std_logic;
signal \N__54916\ : std_logic;
signal \N__54913\ : std_logic;
signal \N__54910\ : std_logic;
signal \N__54907\ : std_logic;
signal \N__54906\ : std_logic;
signal \N__54903\ : std_logic;
signal \N__54900\ : std_logic;
signal \N__54895\ : std_logic;
signal \N__54894\ : std_logic;
signal \N__54893\ : std_logic;
signal \N__54890\ : std_logic;
signal \N__54889\ : std_logic;
signal \N__54886\ : std_logic;
signal \N__54883\ : std_logic;
signal \N__54880\ : std_logic;
signal \N__54877\ : std_logic;
signal \N__54874\ : std_logic;
signal \N__54871\ : std_logic;
signal \N__54866\ : std_logic;
signal \N__54859\ : std_logic;
signal \N__54856\ : std_logic;
signal \N__54853\ : std_logic;
signal \N__54850\ : std_logic;
signal \N__54847\ : std_logic;
signal \N__54844\ : std_logic;
signal \N__54841\ : std_logic;
signal \N__54838\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54832\ : std_logic;
signal \N__54829\ : std_logic;
signal \N__54828\ : std_logic;
signal \N__54825\ : std_logic;
signal \N__54822\ : std_logic;
signal \N__54819\ : std_logic;
signal \N__54816\ : std_logic;
signal \N__54815\ : std_logic;
signal \N__54812\ : std_logic;
signal \N__54809\ : std_logic;
signal \N__54806\ : std_logic;
signal \N__54799\ : std_logic;
signal \N__54796\ : std_logic;
signal \N__54795\ : std_logic;
signal \N__54792\ : std_logic;
signal \N__54789\ : std_logic;
signal \N__54784\ : std_logic;
signal \N__54781\ : std_logic;
signal \N__54778\ : std_logic;
signal \N__54777\ : std_logic;
signal \N__54776\ : std_logic;
signal \N__54773\ : std_logic;
signal \N__54768\ : std_logic;
signal \N__54767\ : std_logic;
signal \N__54766\ : std_logic;
signal \N__54761\ : std_logic;
signal \N__54756\ : std_logic;
signal \N__54751\ : std_logic;
signal \N__54748\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54746\ : std_logic;
signal \N__54743\ : std_logic;
signal \N__54740\ : std_logic;
signal \N__54737\ : std_logic;
signal \N__54734\ : std_logic;
signal \N__54731\ : std_logic;
signal \N__54726\ : std_logic;
signal \N__54723\ : std_logic;
signal \N__54718\ : std_logic;
signal \N__54715\ : std_logic;
signal \N__54714\ : std_logic;
signal \N__54711\ : std_logic;
signal \N__54710\ : std_logic;
signal \N__54709\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54703\ : std_logic;
signal \N__54700\ : std_logic;
signal \N__54697\ : std_logic;
signal \N__54688\ : std_logic;
signal \N__54685\ : std_logic;
signal \N__54684\ : std_logic;
signal \N__54683\ : std_logic;
signal \N__54682\ : std_logic;
signal \N__54679\ : std_logic;
signal \N__54676\ : std_logic;
signal \N__54673\ : std_logic;
signal \N__54670\ : std_logic;
signal \N__54667\ : std_logic;
signal \N__54664\ : std_logic;
signal \N__54663\ : std_logic;
signal \N__54660\ : std_logic;
signal \N__54657\ : std_logic;
signal \N__54654\ : std_logic;
signal \N__54651\ : std_logic;
signal \N__54648\ : std_logic;
signal \N__54643\ : std_logic;
signal \N__54634\ : std_logic;
signal \N__54633\ : std_logic;
signal \N__54630\ : std_logic;
signal \N__54627\ : std_logic;
signal \N__54626\ : std_logic;
signal \N__54623\ : std_logic;
signal \N__54618\ : std_logic;
signal \N__54613\ : std_logic;
signal \N__54610\ : std_logic;
signal \N__54607\ : std_logic;
signal \N__54604\ : std_logic;
signal \N__54601\ : std_logic;
signal \N__54600\ : std_logic;
signal \N__54595\ : std_logic;
signal \N__54592\ : std_logic;
signal \N__54589\ : std_logic;
signal \N__54588\ : std_logic;
signal \N__54587\ : std_logic;
signal \N__54584\ : std_logic;
signal \N__54581\ : std_logic;
signal \N__54578\ : std_logic;
signal \N__54571\ : std_logic;
signal \N__54568\ : std_logic;
signal \N__54565\ : std_logic;
signal \N__54562\ : std_logic;
signal \N__54561\ : std_logic;
signal \N__54558\ : std_logic;
signal \N__54555\ : std_logic;
signal \N__54552\ : std_logic;
signal \N__54549\ : std_logic;
signal \N__54544\ : std_logic;
signal \N__54541\ : std_logic;
signal \N__54538\ : std_logic;
signal \N__54535\ : std_logic;
signal \N__54532\ : std_logic;
signal \N__54529\ : std_logic;
signal \N__54528\ : std_logic;
signal \N__54525\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54519\ : std_logic;
signal \N__54514\ : std_logic;
signal \N__54511\ : std_logic;
signal \N__54508\ : std_logic;
signal \N__54507\ : std_logic;
signal \N__54504\ : std_logic;
signal \N__54501\ : std_logic;
signal \N__54500\ : std_logic;
signal \N__54497\ : std_logic;
signal \N__54494\ : std_logic;
signal \N__54491\ : std_logic;
signal \N__54488\ : std_logic;
signal \N__54481\ : std_logic;
signal \N__54478\ : std_logic;
signal \N__54477\ : std_logic;
signal \N__54474\ : std_logic;
signal \N__54471\ : std_logic;
signal \N__54468\ : std_logic;
signal \N__54467\ : std_logic;
signal \N__54464\ : std_logic;
signal \N__54461\ : std_logic;
signal \N__54458\ : std_logic;
signal \N__54453\ : std_logic;
signal \N__54448\ : std_logic;
signal \N__54447\ : std_logic;
signal \N__54444\ : std_logic;
signal \N__54441\ : std_logic;
signal \N__54436\ : std_logic;
signal \N__54433\ : std_logic;
signal \N__54432\ : std_logic;
signal \N__54429\ : std_logic;
signal \N__54426\ : std_logic;
signal \N__54421\ : std_logic;
signal \N__54420\ : std_logic;
signal \N__54417\ : std_logic;
signal \N__54414\ : std_logic;
signal \N__54411\ : std_logic;
signal \N__54408\ : std_logic;
signal \N__54407\ : std_logic;
signal \N__54404\ : std_logic;
signal \N__54401\ : std_logic;
signal \N__54400\ : std_logic;
signal \N__54399\ : std_logic;
signal \N__54396\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54390\ : std_logic;
signal \N__54387\ : std_logic;
signal \N__54384\ : std_logic;
signal \N__54379\ : std_logic;
signal \N__54374\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54364\ : std_logic;
signal \N__54363\ : std_logic;
signal \N__54360\ : std_logic;
signal \N__54357\ : std_logic;
signal \N__54352\ : std_logic;
signal \N__54349\ : std_logic;
signal \N__54346\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54340\ : std_logic;
signal \N__54337\ : std_logic;
signal \N__54334\ : std_logic;
signal \N__54331\ : std_logic;
signal \N__54328\ : std_logic;
signal \N__54325\ : std_logic;
signal \N__54322\ : std_logic;
signal \N__54321\ : std_logic;
signal \N__54320\ : std_logic;
signal \N__54319\ : std_logic;
signal \N__54316\ : std_logic;
signal \N__54313\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54301\ : std_logic;
signal \N__54300\ : std_logic;
signal \N__54297\ : std_logic;
signal \N__54294\ : std_logic;
signal \N__54289\ : std_logic;
signal \N__54286\ : std_logic;
signal \N__54285\ : std_logic;
signal \N__54284\ : std_logic;
signal \N__54283\ : std_logic;
signal \N__54280\ : std_logic;
signal \N__54277\ : std_logic;
signal \N__54274\ : std_logic;
signal \N__54271\ : std_logic;
signal \N__54262\ : std_logic;
signal \N__54261\ : std_logic;
signal \N__54258\ : std_logic;
signal \N__54255\ : std_logic;
signal \N__54250\ : std_logic;
signal \N__54247\ : std_logic;
signal \N__54244\ : std_logic;
signal \N__54241\ : std_logic;
signal \N__54238\ : std_logic;
signal \N__54235\ : std_logic;
signal \N__54232\ : std_logic;
signal \N__54229\ : std_logic;
signal \N__54226\ : std_logic;
signal \N__54223\ : std_logic;
signal \N__54220\ : std_logic;
signal \N__54217\ : std_logic;
signal \N__54214\ : std_logic;
signal \N__54213\ : std_logic;
signal \N__54210\ : std_logic;
signal \N__54207\ : std_logic;
signal \N__54204\ : std_logic;
signal \N__54201\ : std_logic;
signal \N__54198\ : std_logic;
signal \N__54193\ : std_logic;
signal \N__54190\ : std_logic;
signal \N__54189\ : std_logic;
signal \N__54188\ : std_logic;
signal \N__54185\ : std_logic;
signal \N__54180\ : std_logic;
signal \N__54175\ : std_logic;
signal \N__54174\ : std_logic;
signal \N__54171\ : std_logic;
signal \N__54168\ : std_logic;
signal \N__54165\ : std_logic;
signal \N__54164\ : std_logic;
signal \N__54161\ : std_logic;
signal \N__54158\ : std_logic;
signal \N__54155\ : std_logic;
signal \N__54148\ : std_logic;
signal \N__54145\ : std_logic;
signal \N__54142\ : std_logic;
signal \N__54139\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54135\ : std_logic;
signal \N__54132\ : std_logic;
signal \N__54131\ : std_logic;
signal \N__54130\ : std_logic;
signal \N__54127\ : std_logic;
signal \N__54124\ : std_logic;
signal \N__54119\ : std_logic;
signal \N__54112\ : std_logic;
signal \N__54111\ : std_logic;
signal \N__54108\ : std_logic;
signal \N__54105\ : std_logic;
signal \N__54100\ : std_logic;
signal \N__54097\ : std_logic;
signal \N__54094\ : std_logic;
signal \N__54093\ : std_logic;
signal \N__54090\ : std_logic;
signal \N__54087\ : std_logic;
signal \N__54084\ : std_logic;
signal \N__54079\ : std_logic;
signal \N__54076\ : std_logic;
signal \N__54073\ : std_logic;
signal \N__54070\ : std_logic;
signal \N__54067\ : std_logic;
signal \N__54064\ : std_logic;
signal \N__54061\ : std_logic;
signal \N__54058\ : std_logic;
signal \N__54055\ : std_logic;
signal \N__54054\ : std_logic;
signal \N__54051\ : std_logic;
signal \N__54048\ : std_logic;
signal \N__54043\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54039\ : std_logic;
signal \N__54036\ : std_logic;
signal \N__54031\ : std_logic;
signal \N__54030\ : std_logic;
signal \N__54027\ : std_logic;
signal \N__54024\ : std_logic;
signal \N__54019\ : std_logic;
signal \N__54016\ : std_logic;
signal \N__54015\ : std_logic;
signal \N__54012\ : std_logic;
signal \N__54009\ : std_logic;
signal \N__54008\ : std_logic;
signal \N__54007\ : std_logic;
signal \N__54004\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__53998\ : std_logic;
signal \N__53995\ : std_logic;
signal \N__53986\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53980\ : std_logic;
signal \N__53979\ : std_logic;
signal \N__53976\ : std_logic;
signal \N__53973\ : std_logic;
signal \N__53968\ : std_logic;
signal \N__53965\ : std_logic;
signal \N__53962\ : std_logic;
signal \N__53959\ : std_logic;
signal \N__53956\ : std_logic;
signal \N__53953\ : std_logic;
signal \N__53950\ : std_logic;
signal \N__53947\ : std_logic;
signal \N__53944\ : std_logic;
signal \N__53941\ : std_logic;
signal \N__53940\ : std_logic;
signal \N__53937\ : std_logic;
signal \N__53934\ : std_logic;
signal \N__53931\ : std_logic;
signal \N__53928\ : std_logic;
signal \N__53925\ : std_logic;
signal \N__53920\ : std_logic;
signal \N__53917\ : std_logic;
signal \N__53916\ : std_logic;
signal \N__53913\ : std_logic;
signal \N__53910\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53902\ : std_logic;
signal \N__53901\ : std_logic;
signal \N__53898\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53892\ : std_logic;
signal \N__53889\ : std_logic;
signal \N__53886\ : std_logic;
signal \N__53883\ : std_logic;
signal \N__53880\ : std_logic;
signal \N__53877\ : std_logic;
signal \N__53874\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53866\ : std_logic;
signal \N__53863\ : std_logic;
signal \N__53862\ : std_logic;
signal \N__53859\ : std_logic;
signal \N__53856\ : std_logic;
signal \N__53851\ : std_logic;
signal \N__53848\ : std_logic;
signal \N__53845\ : std_logic;
signal \N__53842\ : std_logic;
signal \N__53839\ : std_logic;
signal \N__53836\ : std_logic;
signal \N__53833\ : std_logic;
signal \N__53830\ : std_logic;
signal \N__53827\ : std_logic;
signal \N__53824\ : std_logic;
signal \N__53821\ : std_logic;
signal \N__53818\ : std_logic;
signal \N__53817\ : std_logic;
signal \N__53814\ : std_logic;
signal \N__53811\ : std_logic;
signal \N__53810\ : std_logic;
signal \N__53809\ : std_logic;
signal \N__53806\ : std_logic;
signal \N__53803\ : std_logic;
signal \N__53800\ : std_logic;
signal \N__53797\ : std_logic;
signal \N__53788\ : std_logic;
signal \N__53787\ : std_logic;
signal \N__53786\ : std_logic;
signal \N__53783\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53777\ : std_logic;
signal \N__53770\ : std_logic;
signal \N__53767\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53763\ : std_logic;
signal \N__53762\ : std_logic;
signal \N__53759\ : std_logic;
signal \N__53756\ : std_logic;
signal \N__53751\ : std_logic;
signal \N__53746\ : std_logic;
signal \N__53743\ : std_logic;
signal \N__53740\ : std_logic;
signal \N__53737\ : std_logic;
signal \N__53734\ : std_logic;
signal \N__53731\ : std_logic;
signal \N__53728\ : std_logic;
signal \N__53727\ : std_logic;
signal \N__53724\ : std_logic;
signal \N__53721\ : std_logic;
signal \N__53720\ : std_logic;
signal \N__53719\ : std_logic;
signal \N__53716\ : std_logic;
signal \N__53713\ : std_logic;
signal \N__53710\ : std_logic;
signal \N__53707\ : std_logic;
signal \N__53700\ : std_logic;
signal \N__53695\ : std_logic;
signal \N__53694\ : std_logic;
signal \N__53691\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53689\ : std_logic;
signal \N__53686\ : std_logic;
signal \N__53683\ : std_logic;
signal \N__53678\ : std_logic;
signal \N__53675\ : std_logic;
signal \N__53672\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53664\ : std_logic;
signal \N__53661\ : std_logic;
signal \N__53656\ : std_logic;
signal \N__53655\ : std_logic;
signal \N__53654\ : std_logic;
signal \N__53651\ : std_logic;
signal \N__53650\ : std_logic;
signal \N__53647\ : std_logic;
signal \N__53644\ : std_logic;
signal \N__53641\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53633\ : std_logic;
signal \N__53630\ : std_logic;
signal \N__53627\ : std_logic;
signal \N__53626\ : std_logic;
signal \N__53623\ : std_logic;
signal \N__53618\ : std_logic;
signal \N__53615\ : std_logic;
signal \N__53612\ : std_logic;
signal \N__53609\ : std_logic;
signal \N__53602\ : std_logic;
signal \N__53601\ : std_logic;
signal \N__53600\ : std_logic;
signal \N__53599\ : std_logic;
signal \N__53598\ : std_logic;
signal \N__53595\ : std_logic;
signal \N__53590\ : std_logic;
signal \N__53587\ : std_logic;
signal \N__53584\ : std_logic;
signal \N__53581\ : std_logic;
signal \N__53576\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53570\ : std_logic;
signal \N__53567\ : std_logic;
signal \N__53560\ : std_logic;
signal \N__53557\ : std_logic;
signal \N__53554\ : std_logic;
signal \N__53551\ : std_logic;
signal \N__53548\ : std_logic;
signal \N__53545\ : std_logic;
signal \N__53542\ : std_logic;
signal \N__53539\ : std_logic;
signal \N__53536\ : std_logic;
signal \N__53533\ : std_logic;
signal \N__53532\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53524\ : std_logic;
signal \N__53521\ : std_logic;
signal \N__53518\ : std_logic;
signal \N__53515\ : std_logic;
signal \N__53512\ : std_logic;
signal \N__53509\ : std_logic;
signal \N__53506\ : std_logic;
signal \N__53503\ : std_logic;
signal \N__53502\ : std_logic;
signal \N__53499\ : std_logic;
signal \N__53496\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53490\ : std_logic;
signal \N__53487\ : std_logic;
signal \N__53482\ : std_logic;
signal \N__53479\ : std_logic;
signal \N__53476\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53472\ : std_logic;
signal \N__53469\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53465\ : std_logic;
signal \N__53464\ : std_logic;
signal \N__53461\ : std_logic;
signal \N__53458\ : std_logic;
signal \N__53457\ : std_logic;
signal \N__53452\ : std_logic;
signal \N__53449\ : std_logic;
signal \N__53448\ : std_logic;
signal \N__53445\ : std_logic;
signal \N__53442\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53436\ : std_logic;
signal \N__53433\ : std_logic;
signal \N__53426\ : std_logic;
signal \N__53423\ : std_logic;
signal \N__53416\ : std_logic;
signal \N__53413\ : std_logic;
signal \N__53410\ : std_logic;
signal \N__53409\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53403\ : std_logic;
signal \N__53400\ : std_logic;
signal \N__53397\ : std_logic;
signal \N__53392\ : std_logic;
signal \N__53389\ : std_logic;
signal \N__53388\ : std_logic;
signal \N__53387\ : std_logic;
signal \N__53386\ : std_logic;
signal \N__53383\ : std_logic;
signal \N__53380\ : std_logic;
signal \N__53375\ : std_logic;
signal \N__53372\ : std_logic;
signal \N__53369\ : std_logic;
signal \N__53368\ : std_logic;
signal \N__53365\ : std_logic;
signal \N__53360\ : std_logic;
signal \N__53357\ : std_logic;
signal \N__53354\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53346\ : std_logic;
signal \N__53343\ : std_logic;
signal \N__53340\ : std_logic;
signal \N__53335\ : std_logic;
signal \N__53332\ : std_logic;
signal \N__53329\ : std_logic;
signal \N__53328\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53322\ : std_logic;
signal \N__53321\ : std_logic;
signal \N__53318\ : std_logic;
signal \N__53315\ : std_logic;
signal \N__53312\ : std_logic;
signal \N__53307\ : std_logic;
signal \N__53302\ : std_logic;
signal \N__53299\ : std_logic;
signal \N__53296\ : std_logic;
signal \N__53293\ : std_logic;
signal \N__53292\ : std_logic;
signal \N__53287\ : std_logic;
signal \N__53286\ : std_logic;
signal \N__53283\ : std_logic;
signal \N__53280\ : std_logic;
signal \N__53279\ : std_logic;
signal \N__53274\ : std_logic;
signal \N__53271\ : std_logic;
signal \N__53268\ : std_logic;
signal \N__53265\ : std_logic;
signal \N__53262\ : std_logic;
signal \N__53257\ : std_logic;
signal \N__53256\ : std_logic;
signal \N__53251\ : std_logic;
signal \N__53248\ : std_logic;
signal \N__53245\ : std_logic;
signal \N__53242\ : std_logic;
signal \N__53241\ : std_logic;
signal \N__53238\ : std_logic;
signal \N__53235\ : std_logic;
signal \N__53232\ : std_logic;
signal \N__53227\ : std_logic;
signal \N__53224\ : std_logic;
signal \N__53221\ : std_logic;
signal \N__53218\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53214\ : std_logic;
signal \N__53211\ : std_logic;
signal \N__53206\ : std_logic;
signal \N__53203\ : std_logic;
signal \N__53200\ : std_logic;
signal \N__53197\ : std_logic;
signal \N__53196\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53194\ : std_logic;
signal \N__53193\ : std_logic;
signal \N__53190\ : std_logic;
signal \N__53189\ : std_logic;
signal \N__53188\ : std_logic;
signal \N__53185\ : std_logic;
signal \N__53182\ : std_logic;
signal \N__53181\ : std_logic;
signal \N__53178\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53175\ : std_logic;
signal \N__53174\ : std_logic;
signal \N__53171\ : std_logic;
signal \N__53170\ : std_logic;
signal \N__53169\ : std_logic;
signal \N__53168\ : std_logic;
signal \N__53165\ : std_logic;
signal \N__53162\ : std_logic;
signal \N__53159\ : std_logic;
signal \N__53156\ : std_logic;
signal \N__53153\ : std_logic;
signal \N__53150\ : std_logic;
signal \N__53147\ : std_logic;
signal \N__53144\ : std_logic;
signal \N__53141\ : std_logic;
signal \N__53138\ : std_logic;
signal \N__53137\ : std_logic;
signal \N__53136\ : std_logic;
signal \N__53135\ : std_logic;
signal \N__53132\ : std_logic;
signal \N__53131\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53128\ : std_logic;
signal \N__53125\ : std_logic;
signal \N__53120\ : std_logic;
signal \N__53117\ : std_logic;
signal \N__53116\ : std_logic;
signal \N__53115\ : std_logic;
signal \N__53110\ : std_logic;
signal \N__53105\ : std_logic;
signal \N__53098\ : std_logic;
signal \N__53093\ : std_logic;
signal \N__53090\ : std_logic;
signal \N__53087\ : std_logic;
signal \N__53084\ : std_logic;
signal \N__53077\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53065\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53053\ : std_logic;
signal \N__53046\ : std_logic;
signal \N__53029\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53027\ : std_logic;
signal \N__53026\ : std_logic;
signal \N__53023\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53021\ : std_logic;
signal \N__53020\ : std_logic;
signal \N__53019\ : std_logic;
signal \N__53016\ : std_logic;
signal \N__53013\ : std_logic;
signal \N__53012\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53006\ : std_logic;
signal \N__53003\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52988\ : std_logic;
signal \N__52985\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52981\ : std_logic;
signal \N__52978\ : std_logic;
signal \N__52975\ : std_logic;
signal \N__52974\ : std_logic;
signal \N__52973\ : std_logic;
signal \N__52972\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52967\ : std_logic;
signal \N__52964\ : std_logic;
signal \N__52961\ : std_logic;
signal \N__52958\ : std_logic;
signal \N__52951\ : std_logic;
signal \N__52948\ : std_logic;
signal \N__52947\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52929\ : std_logic;
signal \N__52924\ : std_logic;
signal \N__52919\ : std_logic;
signal \N__52914\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52902\ : std_logic;
signal \N__52891\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52888\ : std_logic;
signal \N__52887\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52885\ : std_logic;
signal \N__52884\ : std_logic;
signal \N__52881\ : std_logic;
signal \N__52878\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52873\ : std_logic;
signal \N__52872\ : std_logic;
signal \N__52871\ : std_logic;
signal \N__52870\ : std_logic;
signal \N__52869\ : std_logic;
signal \N__52868\ : std_logic;
signal \N__52867\ : std_logic;
signal \N__52864\ : std_logic;
signal \N__52861\ : std_logic;
signal \N__52860\ : std_logic;
signal \N__52859\ : std_logic;
signal \N__52858\ : std_logic;
signal \N__52855\ : std_logic;
signal \N__52852\ : std_logic;
signal \N__52849\ : std_logic;
signal \N__52848\ : std_logic;
signal \N__52847\ : std_logic;
signal \N__52846\ : std_logic;
signal \N__52845\ : std_logic;
signal \N__52844\ : std_logic;
signal \N__52843\ : std_logic;
signal \N__52840\ : std_logic;
signal \N__52837\ : std_logic;
signal \N__52834\ : std_logic;
signal \N__52831\ : std_logic;
signal \N__52828\ : std_logic;
signal \N__52825\ : std_logic;
signal \N__52822\ : std_logic;
signal \N__52819\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52815\ : std_logic;
signal \N__52812\ : std_logic;
signal \N__52809\ : std_logic;
signal \N__52804\ : std_logic;
signal \N__52801\ : std_logic;
signal \N__52798\ : std_logic;
signal \N__52795\ : std_logic;
signal \N__52792\ : std_logic;
signal \N__52787\ : std_logic;
signal \N__52784\ : std_logic;
signal \N__52781\ : std_logic;
signal \N__52778\ : std_logic;
signal \N__52775\ : std_logic;
signal \N__52772\ : std_logic;
signal \N__52769\ : std_logic;
signal \N__52764\ : std_logic;
signal \N__52749\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52744\ : std_logic;
signal \N__52741\ : std_logic;
signal \N__52738\ : std_logic;
signal \N__52731\ : std_logic;
signal \N__52728\ : std_logic;
signal \N__52725\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52703\ : std_logic;
signal \N__52700\ : std_logic;
signal \N__52697\ : std_logic;
signal \N__52694\ : std_logic;
signal \N__52691\ : std_logic;
signal \N__52686\ : std_logic;
signal \N__52679\ : std_logic;
signal \N__52674\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52660\ : std_logic;
signal \N__52659\ : std_logic;
signal \N__52654\ : std_logic;
signal \N__52651\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52649\ : std_logic;
signal \N__52646\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52638\ : std_logic;
signal \N__52633\ : std_logic;
signal \N__52630\ : std_logic;
signal \N__52629\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52623\ : std_logic;
signal \N__52618\ : std_logic;
signal \N__52615\ : std_logic;
signal \N__52612\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52608\ : std_logic;
signal \N__52605\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52597\ : std_logic;
signal \N__52596\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52590\ : std_logic;
signal \N__52585\ : std_logic;
signal \N__52582\ : std_logic;
signal \N__52579\ : std_logic;
signal \N__52576\ : std_logic;
signal \N__52573\ : std_logic;
signal \N__52570\ : std_logic;
signal \N__52567\ : std_logic;
signal \N__52564\ : std_logic;
signal \N__52561\ : std_logic;
signal \N__52558\ : std_logic;
signal \N__52555\ : std_logic;
signal \N__52552\ : std_logic;
signal \N__52549\ : std_logic;
signal \N__52546\ : std_logic;
signal \N__52543\ : std_logic;
signal \N__52540\ : std_logic;
signal \N__52539\ : std_logic;
signal \N__52536\ : std_logic;
signal \N__52535\ : std_logic;
signal \N__52534\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52528\ : std_logic;
signal \N__52525\ : std_logic;
signal \N__52522\ : std_logic;
signal \N__52513\ : std_logic;
signal \N__52510\ : std_logic;
signal \N__52509\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52505\ : std_logic;
signal \N__52502\ : std_logic;
signal \N__52499\ : std_logic;
signal \N__52496\ : std_logic;
signal \N__52493\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52480\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52476\ : std_logic;
signal \N__52475\ : std_logic;
signal \N__52470\ : std_logic;
signal \N__52467\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52461\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52453\ : std_logic;
signal \N__52450\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52443\ : std_logic;
signal \N__52440\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52429\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52414\ : std_logic;
signal \N__52411\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52404\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52392\ : std_logic;
signal \N__52391\ : std_logic;
signal \N__52386\ : std_logic;
signal \N__52383\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52377\ : std_logic;
signal \N__52376\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52367\ : std_logic;
signal \N__52364\ : std_logic;
signal \N__52361\ : std_logic;
signal \N__52358\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52343\ : std_logic;
signal \N__52340\ : std_logic;
signal \N__52335\ : std_logic;
signal \N__52330\ : std_logic;
signal \N__52329\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52323\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52317\ : std_logic;
signal \N__52314\ : std_logic;
signal \N__52309\ : std_logic;
signal \N__52306\ : std_logic;
signal \N__52303\ : std_logic;
signal \N__52300\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52288\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52282\ : std_logic;
signal \N__52279\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52274\ : std_logic;
signal \N__52271\ : std_logic;
signal \N__52268\ : std_logic;
signal \N__52265\ : std_logic;
signal \N__52262\ : std_logic;
signal \N__52259\ : std_logic;
signal \N__52256\ : std_logic;
signal \N__52253\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52229\ : std_logic;
signal \N__52226\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52217\ : std_logic;
signal \N__52210\ : std_logic;
signal \N__52207\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52203\ : std_logic;
signal \N__52202\ : std_logic;
signal \N__52199\ : std_logic;
signal \N__52196\ : std_logic;
signal \N__52193\ : std_logic;
signal \N__52190\ : std_logic;
signal \N__52183\ : std_logic;
signal \N__52180\ : std_logic;
signal \N__52179\ : std_logic;
signal \N__52178\ : std_logic;
signal \N__52175\ : std_logic;
signal \N__52172\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52156\ : std_logic;
signal \N__52149\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52143\ : std_logic;
signal \N__52138\ : std_logic;
signal \N__52135\ : std_logic;
signal \N__52134\ : std_logic;
signal \N__52133\ : std_logic;
signal \N__52132\ : std_logic;
signal \N__52129\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52116\ : std_logic;
signal \N__52111\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52107\ : std_logic;
signal \N__52106\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52098\ : std_logic;
signal \N__52095\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52089\ : std_logic;
signal \N__52086\ : std_logic;
signal \N__52083\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52069\ : std_logic;
signal \N__52068\ : std_logic;
signal \N__52065\ : std_logic;
signal \N__52062\ : std_logic;
signal \N__52059\ : std_logic;
signal \N__52058\ : std_logic;
signal \N__52055\ : std_logic;
signal \N__52054\ : std_logic;
signal \N__52051\ : std_logic;
signal \N__52050\ : std_logic;
signal \N__52047\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52041\ : std_logic;
signal \N__52038\ : std_logic;
signal \N__52035\ : std_logic;
signal \N__52034\ : std_logic;
signal \N__52031\ : std_logic;
signal \N__52028\ : std_logic;
signal \N__52025\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51991\ : std_logic;
signal \N__51990\ : std_logic;
signal \N__51987\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51979\ : std_logic;
signal \N__51978\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51971\ : std_logic;
signal \N__51970\ : std_logic;
signal \N__51967\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51961\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51953\ : std_logic;
signal \N__51950\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51942\ : std_logic;
signal \N__51939\ : std_logic;
signal \N__51938\ : std_logic;
signal \N__51935\ : std_logic;
signal \N__51932\ : std_logic;
signal \N__51927\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51915\ : std_logic;
signal \N__51914\ : std_logic;
signal \N__51911\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51907\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51899\ : std_logic;
signal \N__51892\ : std_logic;
signal \N__51889\ : std_logic;
signal \N__51886\ : std_logic;
signal \N__51883\ : std_logic;
signal \N__51880\ : std_logic;
signal \N__51877\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51865\ : std_logic;
signal \N__51862\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51855\ : std_logic;
signal \N__51854\ : std_logic;
signal \N__51851\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51841\ : std_logic;
signal \N__51838\ : std_logic;
signal \N__51837\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51820\ : std_logic;
signal \N__51819\ : std_logic;
signal \N__51816\ : std_logic;
signal \N__51813\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51802\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51791\ : std_logic;
signal \N__51788\ : std_logic;
signal \N__51785\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51777\ : std_logic;
signal \N__51776\ : std_logic;
signal \N__51775\ : std_logic;
signal \N__51774\ : std_logic;
signal \N__51773\ : std_logic;
signal \N__51768\ : std_logic;
signal \N__51765\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51759\ : std_logic;
signal \N__51756\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51754\ : std_logic;
signal \N__51753\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51744\ : std_logic;
signal \N__51741\ : std_logic;
signal \N__51738\ : std_logic;
signal \N__51733\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51721\ : std_logic;
signal \N__51712\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51710\ : std_logic;
signal \N__51707\ : std_logic;
signal \N__51704\ : std_logic;
signal \N__51701\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51697\ : std_logic;
signal \N__51694\ : std_logic;
signal \N__51691\ : std_logic;
signal \N__51688\ : std_logic;
signal \N__51687\ : std_logic;
signal \N__51686\ : std_logic;
signal \N__51685\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51683\ : std_logic;
signal \N__51680\ : std_logic;
signal \N__51673\ : std_logic;
signal \N__51670\ : std_logic;
signal \N__51665\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51634\ : std_logic;
signal \N__51631\ : std_logic;
signal \N__51630\ : std_logic;
signal \N__51627\ : std_logic;
signal \N__51624\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51622\ : std_logic;
signal \N__51619\ : std_logic;
signal \N__51616\ : std_logic;
signal \N__51613\ : std_logic;
signal \N__51610\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51598\ : std_logic;
signal \N__51597\ : std_logic;
signal \N__51596\ : std_logic;
signal \N__51593\ : std_logic;
signal \N__51592\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51586\ : std_logic;
signal \N__51581\ : std_logic;
signal \N__51578\ : std_logic;
signal \N__51571\ : std_logic;
signal \N__51568\ : std_logic;
signal \N__51567\ : std_logic;
signal \N__51566\ : std_logic;
signal \N__51563\ : std_logic;
signal \N__51560\ : std_logic;
signal \N__51557\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51547\ : std_logic;
signal \N__51544\ : std_logic;
signal \N__51543\ : std_logic;
signal \N__51540\ : std_logic;
signal \N__51537\ : std_logic;
signal \N__51534\ : std_logic;
signal \N__51531\ : std_logic;
signal \N__51526\ : std_logic;
signal \N__51523\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51517\ : std_logic;
signal \N__51514\ : std_logic;
signal \N__51511\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51493\ : std_logic;
signal \N__51490\ : std_logic;
signal \N__51487\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51474\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51471\ : std_logic;
signal \N__51470\ : std_logic;
signal \N__51467\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51464\ : std_logic;
signal \N__51463\ : std_logic;
signal \N__51458\ : std_logic;
signal \N__51455\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51451\ : std_logic;
signal \N__51450\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51448\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51444\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51433\ : std_logic;
signal \N__51426\ : std_logic;
signal \N__51423\ : std_logic;
signal \N__51420\ : std_logic;
signal \N__51417\ : std_logic;
signal \N__51414\ : std_logic;
signal \N__51413\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51411\ : std_logic;
signal \N__51410\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51404\ : std_logic;
signal \N__51403\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51398\ : std_logic;
signal \N__51395\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51388\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51373\ : std_logic;
signal \N__51372\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51367\ : std_logic;
signal \N__51366\ : std_logic;
signal \N__51363\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51351\ : std_logic;
signal \N__51348\ : std_logic;
signal \N__51343\ : std_logic;
signal \N__51340\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51326\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51322\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51304\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51290\ : std_logic;
signal \N__51287\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51267\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51257\ : std_logic;
signal \N__51250\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51239\ : std_logic;
signal \N__51236\ : std_logic;
signal \N__51231\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51193\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51175\ : std_logic;
signal \N__51174\ : std_logic;
signal \N__51173\ : std_logic;
signal \N__51172\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51166\ : std_logic;
signal \N__51163\ : std_logic;
signal \N__51162\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51160\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51151\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51132\ : std_logic;
signal \N__51131\ : std_logic;
signal \N__51130\ : std_logic;
signal \N__51127\ : std_logic;
signal \N__51124\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51122\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51114\ : std_logic;
signal \N__51113\ : std_logic;
signal \N__51112\ : std_logic;
signal \N__51111\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51099\ : std_logic;
signal \N__51098\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51096\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51090\ : std_logic;
signal \N__51089\ : std_logic;
signal \N__51088\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51086\ : std_logic;
signal \N__51085\ : std_logic;
signal \N__51082\ : std_logic;
signal \N__51079\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51071\ : std_logic;
signal \N__51070\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51068\ : std_logic;
signal \N__51067\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51065\ : std_logic;
signal \N__51064\ : std_logic;
signal \N__51061\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51055\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51053\ : std_logic;
signal \N__51052\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51046\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51042\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51036\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51016\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51011\ : std_logic;
signal \N__51010\ : std_logic;
signal \N__51007\ : std_logic;
signal \N__51004\ : std_logic;
signal \N__51001\ : std_logic;
signal \N__50998\ : std_logic;
signal \N__50995\ : std_logic;
signal \N__50988\ : std_logic;
signal \N__50987\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50981\ : std_logic;
signal \N__50980\ : std_logic;
signal \N__50975\ : std_logic;
signal \N__50974\ : std_logic;
signal \N__50973\ : std_logic;
signal \N__50970\ : std_logic;
signal \N__50969\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50963\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50961\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50955\ : std_logic;
signal \N__50954\ : std_logic;
signal \N__50951\ : std_logic;
signal \N__50948\ : std_logic;
signal \N__50945\ : std_logic;
signal \N__50942\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50929\ : std_logic;
signal \N__50924\ : std_logic;
signal \N__50919\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50911\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50888\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50880\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50861\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50846\ : std_logic;
signal \N__50843\ : std_logic;
signal \N__50830\ : std_logic;
signal \N__50827\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50803\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50791\ : std_logic;
signal \N__50784\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50780\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50777\ : std_logic;
signal \N__50768\ : std_logic;
signal \N__50765\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50752\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50739\ : std_logic;
signal \N__50732\ : std_logic;
signal \N__50729\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50709\ : std_logic;
signal \N__50706\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50700\ : std_logic;
signal \N__50699\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50690\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50680\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50674\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50665\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50662\ : std_logic;
signal \N__50661\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50658\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50652\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50643\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50632\ : std_logic;
signal \N__50629\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50620\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50610\ : std_logic;
signal \N__50609\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50591\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50564\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50504\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50475\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50186\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50167\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50139\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50116\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50103\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50080\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50072\ : std_logic;
signal \N__50065\ : std_logic;
signal \N__50062\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50056\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49972\ : std_logic;
signal \N__49969\ : std_logic;
signal \N__49966\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49870\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49664\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49654\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49641\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49635\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49622\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49475\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49472\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49449\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49391\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49275\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49271\ : std_logic;
signal \N__49270\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49256\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49223\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49190\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49166\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49048\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49022\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49006\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49002\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48974\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48938\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48892\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48890\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48847\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48380\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48249\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48058\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48028\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47946\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47557\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47522\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47213\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47186\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47177\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47168\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47159\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47023\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46496\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45601\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45109\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44380\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44287\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42386\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41287\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41048\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \VCCG0\ : std_logic;
signal \CLK_c\ : std_logic;
signal tx_enable : std_logic;
signal \GB_BUFFER_PIN_9_c_THRU_CO\ : std_logic;
signal \LED_c\ : std_logic;
signal \quad_counter1.n26_adj_4207_cascade_\ : std_logic;
signal \quad_counter1.n25_adj_4209\ : std_logic;
signal n12907 : std_logic;
signal \quadB_delayed_adj_4543\ : std_logic;
signal \PIN_13_c\ : std_logic;
signal \n12907_cascade_\ : std_logic;
signal \quad_counter1.n27_adj_4208\ : std_logic;
signal \quad_counter1.n28_adj_4206\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \c0.n19612\ : std_logic;
signal \c0.n19613\ : std_logic;
signal \c0.n19614\ : std_logic;
signal \c0.n19615\ : std_logic;
signal \c0.n19616\ : std_logic;
signal \c0.n19617\ : std_logic;
signal \c0.n19618\ : std_logic;
signal \n23768_cascade_\ : std_logic;
signal \n23897_cascade_\ : std_logic;
signal \n10_adj_4532_cascade_\ : std_logic;
signal \c0.n21322\ : std_logic;
signal rx_i : std_logic;
signal \quad_counter1.n27\ : std_logic;
signal \quad_counter1.n28_cascade_\ : std_logic;
signal \quad_counter1.n25\ : std_logic;
signal \n9818_cascade_\ : std_logic;
signal b_delay_counter_0_adj_4541 : std_logic;
signal n187_adj_4546 : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \quad_counter1.b_delay_counter_1\ : std_logic;
signal \quad_counter1.n19503\ : std_logic;
signal \quad_counter1.b_delay_counter_2\ : std_logic;
signal \quad_counter1.n19504\ : std_logic;
signal \quad_counter1.b_delay_counter_3\ : std_logic;
signal \quad_counter1.n19505\ : std_logic;
signal \quad_counter1.b_delay_counter_4\ : std_logic;
signal \quad_counter1.n19506\ : std_logic;
signal \quad_counter1.b_delay_counter_5\ : std_logic;
signal \quad_counter1.n19507\ : std_logic;
signal \quad_counter1.b_delay_counter_6\ : std_logic;
signal \quad_counter1.n19508\ : std_logic;
signal \quad_counter1.b_delay_counter_7\ : std_logic;
signal \quad_counter1.n19509\ : std_logic;
signal \quad_counter1.n19510\ : std_logic;
signal \quad_counter1.b_delay_counter_8\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \quad_counter1.b_delay_counter_9\ : std_logic;
signal \quad_counter1.n19511\ : std_logic;
signal \quad_counter1.b_delay_counter_10\ : std_logic;
signal \quad_counter1.n19512\ : std_logic;
signal \quad_counter1.b_delay_counter_11\ : std_logic;
signal \quad_counter1.n19513\ : std_logic;
signal \quad_counter1.b_delay_counter_12\ : std_logic;
signal \quad_counter1.n19514\ : std_logic;
signal \quad_counter1.b_delay_counter_13\ : std_logic;
signal \quad_counter1.n19515\ : std_logic;
signal \quad_counter1.b_delay_counter_14\ : std_logic;
signal \quad_counter1.n19516\ : std_logic;
signal \quad_counter1.n19517\ : std_logic;
signal \quad_counter1.b_delay_counter_15\ : std_logic;
signal n14377 : std_logic;
signal \b_delay_counter_15__N_4141_adj_4548\ : std_logic;
signal \quad_counter1.A_delayed\ : std_logic;
signal \B_filtered_adj_4539\ : std_logic;
signal \count_enable_adj_4544_cascade_\ : std_logic;
signal data_out_frame_10_6 : std_logic;
signal n26 : std_logic;
signal \n24118_cascade_\ : std_logic;
signal \c0.n23950_cascade_\ : std_logic;
signal \c0.n24147_cascade_\ : std_logic;
signal \c0.n23882\ : std_logic;
signal n24150 : std_logic;
signal \n24097_cascade_\ : std_logic;
signal n24117 : std_logic;
signal n24112 : std_logic;
signal \n23849_cascade_\ : std_logic;
signal data_out_frame_10_3 : std_logic;
signal \c0.n24159_cascade_\ : std_logic;
signal \c0.n24162\ : std_logic;
signal \c0.n11_adj_4355\ : std_logic;
signal n23846 : std_logic;
signal \n24114_cascade_\ : std_logic;
signal n10 : std_logic;
signal \c0.n23895\ : std_logic;
signal \c0.n24051_cascade_\ : std_logic;
signal \c0.n23844\ : std_logic;
signal \c0.n23847\ : std_logic;
signal \c0.n11_adj_4348\ : std_logic;
signal n24102 : std_logic;
signal \c0.n24047\ : std_logic;
signal \c0.n5_adj_4358\ : std_logic;
signal data_out_frame_6_7 : std_logic;
signal data_out_frame_0_3 : std_logic;
signal \c0.n24011\ : std_logic;
signal data_out_frame_0_2 : std_logic;
signal \c0.n6_adj_4521\ : std_logic;
signal \c0.n23859_cascade_\ : std_logic;
signal \n23861_cascade_\ : std_logic;
signal n10_adj_4534 : std_logic;
signal \c0.n5_adj_4522\ : std_logic;
signal data_out_frame_6_2 : std_logic;
signal \c0.n24007\ : std_logic;
signal \c0.n6\ : std_logic;
signal \r_Tx_Data_6\ : std_logic;
signal \r_Tx_Data_2\ : std_logic;
signal \b_delay_counter_15__N_4141_cascade_\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \quad_counter1.a_delay_counter_1\ : std_logic;
signal \quad_counter1.n19518\ : std_logic;
signal \quad_counter1.a_delay_counter_2\ : std_logic;
signal \quad_counter1.n19519\ : std_logic;
signal \quad_counter1.a_delay_counter_3\ : std_logic;
signal \quad_counter1.n19520\ : std_logic;
signal \quad_counter1.a_delay_counter_4\ : std_logic;
signal \quad_counter1.n19521\ : std_logic;
signal \quad_counter1.a_delay_counter_5\ : std_logic;
signal \quad_counter1.n19522\ : std_logic;
signal \quad_counter1.n19523\ : std_logic;
signal \quad_counter1.a_delay_counter_7\ : std_logic;
signal \quad_counter1.n19524\ : std_logic;
signal \quad_counter1.n19525\ : std_logic;
signal \quad_counter1.a_delay_counter_8\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \quad_counter1.n19526\ : std_logic;
signal \quad_counter1.a_delay_counter_10\ : std_logic;
signal \quad_counter1.n19527\ : std_logic;
signal \quad_counter1.a_delay_counter_11\ : std_logic;
signal \quad_counter1.n19528\ : std_logic;
signal \quad_counter1.n19529\ : std_logic;
signal \quad_counter1.n19530\ : std_logic;
signal \quad_counter1.a_delay_counter_14\ : std_logic;
signal \quad_counter1.n19531\ : std_logic;
signal \quad_counter1.n19532\ : std_logic;
signal \quad_counter1.a_delay_counter_15\ : std_logic;
signal data_out_frame_11_6 : std_logic;
signal \A_filtered_adj_4538\ : std_logic;
signal \quad_counter1.B_delayed\ : std_logic;
signal n39_adj_4545 : std_logic;
signal a_delay_counter_0_adj_4540 : std_logic;
signal \c0.n22048_cascade_\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal encoder1_position_0 : std_logic;
signal \quad_counter1.count_direction\ : std_logic;
signal n2205 : std_logic;
signal \quad_counter1.n19548\ : std_logic;
signal \quad_counter1.n19549\ : std_logic;
signal n2203 : std_logic;
signal \quad_counter1.n19550\ : std_logic;
signal n2202 : std_logic;
signal \quad_counter1.n19551\ : std_logic;
signal \quad_counter1.n19552\ : std_logic;
signal n2200 : std_logic;
signal \quad_counter1.n19553\ : std_logic;
signal n2199 : std_logic;
signal \quad_counter1.n19554\ : std_logic;
signal \quad_counter1.n19555\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \quad_counter1.n19556\ : std_logic;
signal \quad_counter1.n19557\ : std_logic;
signal \quad_counter1.n19558\ : std_logic;
signal \quad_counter1.n19559\ : std_logic;
signal \quad_counter1.n19560\ : std_logic;
signal \quad_counter1.n19561\ : std_logic;
signal n2191 : std_logic;
signal \quad_counter1.n19562\ : std_logic;
signal \quad_counter1.n19563\ : std_logic;
signal n2190 : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \quad_counter1.n19564\ : std_logic;
signal \quad_counter1.n19565\ : std_logic;
signal n2187 : std_logic;
signal \quad_counter1.n19566\ : std_logic;
signal \quad_counter1.n19567\ : std_logic;
signal \quad_counter1.n19568\ : std_logic;
signal \quad_counter1.n19569\ : std_logic;
signal n2183 : std_logic;
signal \quad_counter1.n19570\ : std_logic;
signal \quad_counter1.n19571\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \quad_counter1.n19572\ : std_logic;
signal \quad_counter1.n19573\ : std_logic;
signal n2179 : std_logic;
signal \quad_counter1.n19574\ : std_logic;
signal \quad_counter1.n19575\ : std_logic;
signal n2177 : std_logic;
signal \quad_counter1.n19576\ : std_logic;
signal \quad_counter1.n19577\ : std_logic;
signal \quad_counter1.n19578\ : std_logic;
signal \quad_counter1.n19579\ : std_logic;
signal \quad_counter1.n2140\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal n2174 : std_logic;
signal data_out_frame_0_4 : std_logic;
signal data_out_frame_13_5 : std_logic;
signal data_out_frame_9_3 : std_logic;
signal \c0.n24171\ : std_logic;
signal \c0.n24174\ : std_logic;
signal \c0.n23856\ : std_logic;
signal n24108 : std_logic;
signal \n23858_cascade_\ : std_logic;
signal \r_Tx_Data_5\ : std_logic;
signal \r_Tx_Data_4\ : std_logic;
signal n10_adj_4533 : std_logic;
signal data_out_frame_9_2 : std_logic;
signal \c0.n24180_cascade_\ : std_logic;
signal n24106 : std_logic;
signal data_out_frame_7_0 : std_logic;
signal data_out_frame_6_0 : std_logic;
signal n10_adj_4536 : std_logic;
signal \c0.n5_adj_4422\ : std_logic;
signal \c0.n24059\ : std_logic;
signal \c0.n23850_cascade_\ : std_logic;
signal \n23852_cascade_\ : std_logic;
signal byte_transmit_counter_3 : std_logic;
signal \n10_adj_4537_cascade_\ : std_logic;
signal n24110 : std_logic;
signal \r_Tx_Data_0\ : std_logic;
signal n24195 : std_logic;
signal \n24100_cascade_\ : std_logic;
signal n16706 : std_logic;
signal \c0.tx.n23985_cascade_\ : std_logic;
signal \c0.tx.n31_adj_4216_cascade_\ : std_logic;
signal n187 : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \quad_counter0.n19473\ : std_logic;
signal \quad_counter0.n19474\ : std_logic;
signal \quad_counter0.n19475\ : std_logic;
signal \quad_counter0.n19476\ : std_logic;
signal \quad_counter0.n19477\ : std_logic;
signal \quad_counter0.n19478\ : std_logic;
signal \quad_counter0.n19479\ : std_logic;
signal \quad_counter0.n19480\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \quad_counter0.n19481\ : std_logic;
signal \quad_counter0.n19482\ : std_logic;
signal \quad_counter0.n19483\ : std_logic;
signal \quad_counter0.n19484\ : std_logic;
signal \quad_counter0.n19485\ : std_logic;
signal \quad_counter0.n19486\ : std_logic;
signal \quad_counter0.n19487\ : std_logic;
signal n14198 : std_logic;
signal \b_delay_counter_15__N_4141\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \quad_counter0.n19488\ : std_logic;
signal \quad_counter0.n19489\ : std_logic;
signal \quad_counter0.n19490\ : std_logic;
signal \quad_counter0.n19491\ : std_logic;
signal \quad_counter0.n19492\ : std_logic;
signal \quad_counter0.n19493\ : std_logic;
signal \quad_counter0.n19494\ : std_logic;
signal \quad_counter0.n19495\ : std_logic;
signal \bfn_10_25_0_\ : std_logic;
signal \quad_counter0.n19496\ : std_logic;
signal \quad_counter0.n19497\ : std_logic;
signal \quad_counter0.n19498\ : std_logic;
signal \quad_counter0.n19499\ : std_logic;
signal \quad_counter0.n19500\ : std_logic;
signal \quad_counter0.n19501\ : std_logic;
signal \quad_counter0.n19502\ : std_logic;
signal \c0.n24_adj_4502\ : std_logic;
signal \c0.n18_adj_4414_cascade_\ : std_logic;
signal \c0.n13360\ : std_logic;
signal \c0.n23550_cascade_\ : std_logic;
signal \c0.n22_adj_4503_cascade_\ : std_logic;
signal \c0.n26_adj_4504\ : std_logic;
signal \c0.n26_adj_4517\ : std_logic;
signal \c0.n21305_cascade_\ : std_logic;
signal \c0.data_out_frame_28_2\ : std_logic;
signal \c0.n6_adj_4515\ : std_logic;
signal \c0.n12532_cascade_\ : std_logic;
signal \c0.n22126_cascade_\ : std_logic;
signal \c0.data_out_frame_28_4\ : std_logic;
signal \quad_counter1.a_delay_counter_12\ : std_logic;
signal \quad_counter1.a_delay_counter_13\ : std_logic;
signal \quad_counter1.a_delay_counter_9\ : std_logic;
signal \quad_counter1.a_delay_counter_6\ : std_logic;
signal \quad_counter1.n26\ : std_logic;
signal \a_delay_counter_15__N_4124_adj_4547\ : std_logic;
signal \quadA_delayed_adj_4542\ : std_logic;
signal \PIN_12_c\ : std_logic;
signal \a_delay_counter_15__N_4124_adj_4547_cascade_\ : std_logic;
signal n9818 : std_logic;
signal n14228 : std_logic;
signal data_out_frame_29_2 : std_logic;
signal n2196 : std_logic;
signal \c0.n13079_cascade_\ : std_logic;
signal \c0.n22116\ : std_logic;
signal \c0.n6_adj_4308\ : std_logic;
signal data_out_frame_13_0 : std_logic;
signal \c0.n11_adj_4424\ : std_logic;
signal \c0.n6_adj_4335_cascade_\ : std_logic;
signal \c0.n21229_cascade_\ : std_logic;
signal n2193 : std_logic;
signal \c0.n6_adj_4309\ : std_logic;
signal n2204 : std_logic;
signal \c0.n6_adj_4310_cascade_\ : std_logic;
signal \c0.n22037\ : std_logic;
signal encoder1_position_15 : std_logic;
signal data_out_frame_12_7 : std_logic;
signal \c0.n11_adj_4360\ : std_logic;
signal n2197 : std_logic;
signal \c0.n5_adj_4227\ : std_logic;
signal data_out_frame_7_4 : std_logic;
signal \c0.data_out_frame_29__7__N_850\ : std_logic;
signal data_out_frame_11_4 : std_logic;
signal \c0.n23881\ : std_logic;
signal n2189 : std_logic;
signal encoder1_position_16 : std_logic;
signal data_out_frame_10_4 : std_logic;
signal data_out_frame_7_2 : std_logic;
signal n2188 : std_logic;
signal n2184 : std_logic;
signal n2182 : std_logic;
signal n2176 : std_logic;
signal data_out_frame_29_3 : std_logic;
signal data_out_frame_28_3 : std_logic;
signal \c0.n26\ : std_logic;
signal n2175 : std_logic;
signal data_out_frame_7_5 : std_logic;
signal \c0.n5_adj_4346\ : std_logic;
signal data_out_frame_9_7 : std_logic;
signal tx_o : std_logic;
signal \c0.n6_adj_4392\ : std_logic;
signal \c0.byte_transmit_counter_6\ : std_logic;
signal \c0.n23574_cascade_\ : std_logic;
signal \c0.byte_transmit_counter_7\ : std_logic;
signal \c0.n38_adj_4387_cascade_\ : std_logic;
signal data_out_frame_5_2 : std_logic;
signal n23768 : std_logic;
signal byte_transmit_counter_4 : std_logic;
signal n23864 : std_logic;
signal data_out_frame_5_6 : std_logic;
signal data_out_frame_13_3 : std_logic;
signal \c0.n11_adj_4218\ : std_logic;
signal data_out_frame_11_5 : std_logic;
signal data_out_frame_9_5 : std_logic;
signal \c0.n24141_cascade_\ : std_logic;
signal data_out_frame_8_5 : std_logic;
signal \c0.n24144\ : std_logic;
signal \r_Tx_Data_7\ : std_logic;
signal \r_Tx_Data_3\ : std_logic;
signal \r_Bit_Index_2_adj_4551\ : std_logic;
signal n4_adj_4554 : std_logic;
signal \n24189_cascade_\ : std_logic;
signal \r_Bit_Index_1_adj_4552\ : std_logic;
signal n10_adj_4535 : std_logic;
signal byte_transmit_counter_5 : std_logic;
signal \r_Tx_Data_1\ : std_logic;
signal data_in_0_7 : std_logic;
signal data_out_frame_5_3 : std_logic;
signal data_out_frame_6_3 : std_logic;
signal \c0.n5\ : std_logic;
signal data_out_frame_5_5 : std_logic;
signal data_out_frame_11_0 : std_logic;
signal \c0.n24165_cascade_\ : std_logic;
signal \c0.n24168\ : std_logic;
signal \quad_counter0.b_delay_counter_3\ : std_logic;
signal \quad_counter0.b_delay_counter_9\ : std_logic;
signal \quad_counter0.b_delay_counter_4\ : std_logic;
signal b_delay_counter_0 : std_logic;
signal \PIN_8_c\ : std_logic;
signal \quadB_delayed\ : std_logic;
signal \B_filtered\ : std_logic;
signal \quad_counter0.b_delay_counter_13\ : std_logic;
signal \quad_counter0.b_delay_counter_1\ : std_logic;
signal \quad_counter0.b_delay_counter_2\ : std_logic;
signal \quad_counter0.b_delay_counter_5\ : std_logic;
signal \quad_counter0.b_delay_counter_11\ : std_logic;
signal \quad_counter0.b_delay_counter_10\ : std_logic;
signal \quad_counter0.b_delay_counter_8\ : std_logic;
signal \quad_counter0.b_delay_counter_6\ : std_logic;
signal \quad_counter0.n28_adj_4198\ : std_logic;
signal \quad_counter0.n26_adj_4199_cascade_\ : std_logic;
signal \quad_counter0.n25_adj_4201\ : std_logic;
signal n12909 : std_logic;
signal \quad_counter0.A_delayed\ : std_logic;
signal \quad_counter0.B_delayed\ : std_logic;
signal \quad_counter0.a_delay_counter_3\ : std_logic;
signal \quad_counter0.a_delay_counter_8\ : std_logic;
signal \quad_counter0.a_delay_counter_2\ : std_logic;
signal \quad_counter0.a_delay_counter_1\ : std_logic;
signal \quad_counter0.a_delay_counter_5\ : std_logic;
signal \quad_counter0.a_delay_counter_11\ : std_logic;
signal \quad_counter0.a_delay_counter_4\ : std_logic;
signal \A_filtered\ : std_logic;
signal \PIN_7_c\ : std_logic;
signal \quadA_delayed\ : std_logic;
signal n14421 : std_logic;
signal \a_delay_counter_15__N_4124\ : std_logic;
signal n39 : std_logic;
signal \n14421_cascade_\ : std_logic;
signal a_delay_counter_0 : std_logic;
signal \quad_counter0.a_delay_counter_14\ : std_logic;
signal \quad_counter0.a_delay_counter_15\ : std_logic;
signal \quad_counter0.a_delay_counter_7\ : std_logic;
signal \quad_counter0.a_delay_counter_10\ : std_logic;
signal \quad_counter0.n28_adj_4202\ : std_logic;
signal \quad_counter0.n27_adj_4204_cascade_\ : std_logic;
signal \quad_counter0.n25_adj_4205\ : std_logic;
signal n9821 : std_logic;
signal \quad_counter0.a_delay_counter_12\ : std_logic;
signal \quad_counter0.a_delay_counter_13\ : std_logic;
signal \quad_counter0.a_delay_counter_6\ : std_logic;
signal \quad_counter0.a_delay_counter_9\ : std_logic;
signal \quad_counter0.n26_adj_4203\ : std_logic;
signal \data_out_frame_28__3__N_1881\ : std_logic;
signal \c0.n20257\ : std_logic;
signal \c0.n21062\ : std_logic;
signal \c0.data_out_frame_28_1\ : std_logic;
signal \c0.data_out_frame_29_1\ : std_logic;
signal \c0.n26_adj_4519\ : std_logic;
signal \c0.n12542_cascade_\ : std_logic;
signal \c0.n14_adj_4340_cascade_\ : std_logic;
signal \c0.n20320\ : std_logic;
signal \c0.n20320_cascade_\ : std_logic;
signal \c0.n22180_cascade_\ : std_logic;
signal \c0.n10498_cascade_\ : std_logic;
signal \c0.n20253_cascade_\ : std_logic;
signal \c0.n21229\ : std_logic;
signal \c0.n15_adj_4513\ : std_logic;
signal \c0.n22066\ : std_logic;
signal encoder1_position_3 : std_logic;
signal \c0.n21071_cascade_\ : std_logic;
signal \data_out_frame_29__2__N_1749\ : std_logic;
signal \c0.n17_adj_4501\ : std_logic;
signal \c0.data_out_frame_29_0\ : std_logic;
signal \c0.n26_adj_4423\ : std_logic;
signal \c0.n16_adj_4500\ : std_logic;
signal \c0.n10422\ : std_logic;
signal \c0.n6_adj_4313_cascade_\ : std_logic;
signal \c0.n21156_cascade_\ : std_logic;
signal \c0.n21175_cascade_\ : std_logic;
signal \c0.n20276_cascade_\ : std_logic;
signal \c0.n21110_cascade_\ : std_logic;
signal \c0.n14_adj_4514\ : std_logic;
signal encoder1_position_22 : std_logic;
signal n2201 : std_logic;
signal \c0.n22277\ : std_logic;
signal \c0.n22102_cascade_\ : std_logic;
signal \c0.n22293\ : std_logic;
signal \c0.n15_adj_4325_cascade_\ : std_logic;
signal \c0.n21041\ : std_logic;
signal \c0.n21041_cascade_\ : std_logic;
signal \c0.n22102\ : std_logic;
signal \c0.n22361_cascade_\ : std_logic;
signal \c0.n10_adj_4314\ : std_logic;
signal encoder1_position_21 : std_logic;
signal \c0.n24153\ : std_logic;
signal data_out_frame_8_6 : std_logic;
signal \c0.n24156\ : std_logic;
signal data_out_frame_12_6 : std_logic;
signal data_out_frame_11_3 : std_logic;
signal n2181 : std_logic;
signal \c0.n22224\ : std_logic;
signal \c0.n22224_cascade_\ : std_logic;
signal \c0.n13349_cascade_\ : std_logic;
signal \c0.n6_adj_4334\ : std_logic;
signal n24104 : std_logic;
signal \c0.n22405\ : std_logic;
signal encoder1_position_31 : std_logic;
signal data_out_frame_10_7 : std_logic;
signal data_out_frame_8_7 : std_logic;
signal data_out_frame_11_7 : std_logic;
signal data_out_frame_12_3 : std_logic;
signal \c0.n7_adj_4492_cascade_\ : std_logic;
signal data_in_1_5 : std_logic;
signal \c0.n9_adj_4493\ : std_logic;
signal \c0.n23600\ : std_logic;
signal data_in_0_6 : std_logic;
signal data_in_2_2 : std_logic;
signal data_in_0_3 : std_logic;
signal \c0.n14_adj_4495_cascade_\ : std_logic;
signal \c0.n15_adj_4496\ : std_logic;
signal \c0.n10_adj_4231_cascade_\ : std_logic;
signal \c0.n14\ : std_logic;
signal n9539 : std_logic;
signal data_out_frame_10_0 : std_logic;
signal data_in_3_3 : std_logic;
signal encoder1_position_18 : std_logic;
signal data_out_frame_11_2 : std_logic;
signal \c0.n24177\ : std_logic;
signal data_out_frame_5_0 : std_logic;
signal encoder1_position_29 : std_logic;
signal data_out_frame_10_5 : std_logic;
signal \c0.tx.n16631_cascade_\ : std_logic;
signal n14442 : std_logic;
signal \c0.n21370\ : std_logic;
signal \c0.n21376\ : std_logic;
signal \c0.n21362\ : std_logic;
signal \c0.n21128\ : std_logic;
signal \c0.n12_adj_4516\ : std_logic;
signal \c0.n9_adj_4339\ : std_logic;
signal \c0.n22018_cascade_\ : std_logic;
signal \c0.n21946\ : std_logic;
signal \c0.n21946_cascade_\ : std_logic;
signal \c0.n12532\ : std_logic;
signal \c0.n12491_cascade_\ : std_logic;
signal \c0.data_out_frame_28_6\ : std_logic;
signal \c0.n26_adj_4351\ : std_logic;
signal \c0.n7_adj_4307_cascade_\ : std_logic;
signal \data_out_frame_29__3__N_1662\ : std_logic;
signal \c0.n22024\ : std_logic;
signal \c0.data_out_frame_29_4\ : std_logic;
signal \c0.n22151\ : std_logic;
signal \c0.n22151_cascade_\ : std_logic;
signal \c0.n6_adj_4397_cascade_\ : std_logic;
signal \c0.data_out_frame_28_0\ : std_logic;
signal \c0.n22018\ : std_logic;
signal \c0.data_out_frame_29_5\ : std_logic;
signal \c0.data_out_frame_28_5\ : std_logic;
signal \c0.n26_adj_4347\ : std_logic;
signal \c0.n20376\ : std_logic;
signal \c0.n6_adj_4509_cascade_\ : std_logic;
signal \c0.n22393\ : std_logic;
signal \c0.n10498\ : std_logic;
signal \c0.n22393_cascade_\ : std_logic;
signal \c0.n14_adj_4510_cascade_\ : std_logic;
signal \c0.n10462\ : std_logic;
signal \c0.n21150\ : std_logic;
signal \c0.n10_adj_4511\ : std_logic;
signal \c0.n10_adj_4330\ : std_logic;
signal \c0.n21192_cascade_\ : std_logic;
signal \c0.n20931_cascade_\ : std_logic;
signal \c0.n21175\ : std_logic;
signal \c0.n21156\ : std_logic;
signal \c0.n12554\ : std_logic;
signal \c0.n20931\ : std_logic;
signal \c0.n22991\ : std_logic;
signal \c0.n21189_cascade_\ : std_logic;
signal \c0.n21058\ : std_logic;
signal \c0.n21192\ : std_logic;
signal \c0.n13349\ : std_logic;
signal \c0.n13480_cascade_\ : std_logic;
signal \c0.n21122_cascade_\ : std_logic;
signal encoder1_position_14 : std_logic;
signal \c0.n20767\ : std_logic;
signal \c0.n20767_cascade_\ : std_logic;
signal encoder1_position_24 : std_logic;
signal n2195 : std_logic;
signal data_out_frame_9_6 : std_logic;
signal data_out_frame_13_6 : std_logic;
signal n2194 : std_logic;
signal \c0.n11\ : std_logic;
signal \c0.n14_adj_4329\ : std_logic;
signal n2198 : std_logic;
signal n2192 : std_logic;
signal n2186 : std_logic;
signal encoder1_position_19 : std_logic;
signal \c0.n19_adj_4319\ : std_logic;
signal \c0.n23557\ : std_logic;
signal n2180 : std_logic;
signal \c0.n21914_cascade_\ : std_logic;
signal \c0.n21_adj_4320\ : std_logic;
signal data_out_frame_8_4 : std_logic;
signal \c0.n23880\ : std_logic;
signal data_out_frame_9_4 : std_logic;
signal n2178 : std_logic;
signal encoder1_position_27 : std_logic;
signal data_out_frame_10_2 : std_logic;
signal data_out_frame_5_4 : std_logic;
signal data_out_frame_6_4 : std_logic;
signal \c0.n13003\ : std_logic;
signal \c0.n19_adj_4367\ : std_logic;
signal \c0.n20_adj_4362_cascade_\ : std_logic;
signal \c0.n23834\ : std_logic;
signal data_in_1_2 : std_logic;
signal data_in_0_5 : std_logic;
signal data_in_1_6 : std_logic;
signal \c0.n17_adj_4479_cascade_\ : std_logic;
signal \c0.n13023\ : std_logic;
signal data_in_0_2 : std_logic;
signal \c0.n13006\ : std_logic;
signal \c0.n21767\ : std_logic;
signal \c0.tx.n14296\ : std_logic;
signal data_in_1_0 : std_logic;
signal data_in_0_0 : std_logic;
signal data_in_0_4 : std_logic;
signal data_in_1_7 : std_logic;
signal \c0.n10_adj_4494\ : std_logic;
signal \c0.n16_adj_4476\ : std_logic;
signal \c0.n17_adj_4477\ : std_logic;
signal \r_Bit_Index_0_adj_4553\ : std_logic;
signal n24192 : std_logic;
signal n24198 : std_logic;
signal \o_Tx_Serial_N_3783_cascade_\ : std_logic;
signal \c0.tx.n12\ : std_logic;
signal \r_SM_Main_1_adj_4550\ : std_logic;
signal \c0.tx.n6_adj_4214_cascade_\ : std_logic;
signal \c0.tx.n16630\ : std_logic;
signal \n8_cascade_\ : std_logic;
signal \c0.tx.n6_cascade_\ : std_logic;
signal \c0.tx.n31\ : std_logic;
signal \c0.tx.n31_cascade_\ : std_logic;
signal \c0.tx.n47\ : std_logic;
signal \c0.tx.n10\ : std_logic;
signal \c0.tx.r_Clock_Count_0\ : std_logic;
signal \c0.tx.n23960\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \c0.tx.r_Clock_Count_1\ : std_logic;
signal \c0.tx.n23961\ : std_logic;
signal \c0.tx.n19540\ : std_logic;
signal \c0.tx.r_Clock_Count_2\ : std_logic;
signal \c0.tx.n23958\ : std_logic;
signal \c0.tx.n19541\ : std_logic;
signal \c0.tx.r_Clock_Count_3\ : std_logic;
signal \c0.tx.n23963\ : std_logic;
signal \c0.tx.n19542\ : std_logic;
signal \c0.tx.r_Clock_Count_4\ : std_logic;
signal \c0.tx.n23953\ : std_logic;
signal \c0.tx.n19543\ : std_logic;
signal \r_Clock_Count_5\ : std_logic;
signal n316 : std_logic;
signal \c0.tx.n19544\ : std_logic;
signal \c0.tx.n19545\ : std_logic;
signal \r_Clock_Count_7\ : std_logic;
signal n314 : std_logic;
signal \c0.tx.n19546\ : std_logic;
signal \c0.tx.n19547\ : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal \c0.n12878\ : std_logic;
signal \c0.n21360\ : std_logic;
signal \c0.n21356\ : std_logic;
signal \c0.n22317\ : std_logic;
signal \c0.n6_adj_4305\ : std_logic;
signal \c0.n24119\ : std_logic;
signal \c0.n21050\ : std_logic;
signal \c0.n6_adj_4402\ : std_logic;
signal \c0.n22188\ : std_logic;
signal \c0.n20658_cascade_\ : std_logic;
signal \c0.n22166\ : std_logic;
signal \c0.n10467\ : std_logic;
signal \c0.n22180\ : std_logic;
signal \c0.n20330\ : std_logic;
signal \c0.n10434\ : std_logic;
signal \c0.n10513\ : std_logic;
signal \c0.n21189\ : std_logic;
signal \c0.n21135\ : std_logic;
signal \c0.n21219\ : std_logic;
signal \c0.n21811\ : std_logic;
signal \c0.n21135_cascade_\ : std_logic;
signal \c0.n6_adj_4497_cascade_\ : std_logic;
signal \c0.n20151\ : std_logic;
signal \c0.data_out_frame_29_6\ : std_logic;
signal \c0.n21848\ : std_logic;
signal \c0.n20253\ : std_logic;
signal \c0.n21852_cascade_\ : std_logic;
signal \c0.n22346\ : std_logic;
signal \c0.n22126\ : std_logic;
signal \c0.n20298\ : std_logic;
signal \c0.n10_adj_4512_cascade_\ : std_logic;
signal \c0.n10496\ : std_logic;
signal \c0.n20274\ : std_logic;
signal \c0.n21231\ : std_logic;
signal \c0.n22736\ : std_logic;
signal \c0.n21162_cascade_\ : std_logic;
signal \c0.n12526\ : std_logic;
signal \c0.n20201\ : std_logic;
signal \c0.n21876\ : std_logic;
signal data_out_frame_13_7 : std_logic;
signal \c0.n21056\ : std_logic;
signal \c0.n22177\ : std_logic;
signal \c0.n22072\ : std_logic;
signal \c0.n22072_cascade_\ : std_logic;
signal \c0.n22073\ : std_logic;
signal \c0.n20175\ : std_logic;
signal \c0.n20249_cascade_\ : std_logic;
signal \c0.n12528\ : std_logic;
signal \c0.n21065\ : std_logic;
signal \c0.n21842\ : std_logic;
signal \c0.n20230\ : std_logic;
signal \c0.n6_adj_4394\ : std_logic;
signal encoder1_position_5 : std_logic;
signal \c0.n22163_cascade_\ : std_logic;
signal \c0.n20_adj_4505\ : std_logic;
signal \c0.n19_adj_4506_cascade_\ : std_logic;
signal \c0.n21283\ : std_logic;
signal \c0.n6_adj_4508\ : std_logic;
signal \c0.n21116\ : std_logic;
signal \c0.n20819\ : std_logic;
signal \c0.n21_adj_4507\ : std_logic;
signal \c0.n20276\ : std_logic;
signal \c0.n21122\ : std_logic;
signal \c0.n21166\ : std_logic;
signal \c0.n13480\ : std_logic;
signal \c0.n22078\ : std_logic;
signal encoder1_position_9 : std_logic;
signal \c0.n21112\ : std_logic;
signal \c0.n21253\ : std_logic;
signal \c0.n20180_cascade_\ : std_logic;
signal \c0.data_out_frame_29__7__N_1144\ : std_logic;
signal \c0.n20465\ : std_logic;
signal \c0.n21943\ : std_logic;
signal \c0.n21196\ : std_logic;
signal encoder1_position_25 : std_logic;
signal encoder1_position_11 : std_logic;
signal \c0.n20232_cascade_\ : std_logic;
signal \c0.n21146\ : std_logic;
signal \c0.n21146_cascade_\ : std_logic;
signal encoder1_position_23 : std_logic;
signal \c0.n20232\ : std_logic;
signal \c0.n20744\ : std_logic;
signal encoder1_position_1 : std_logic;
signal \c0.n20160\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \quad_counter0.count_direction\ : std_logic;
signal \quad_counter0.n19580\ : std_logic;
signal n2270 : std_logic;
signal \quad_counter0.n19581\ : std_logic;
signal n2269 : std_logic;
signal \quad_counter0.n19582\ : std_logic;
signal n2268 : std_logic;
signal \quad_counter0.n19583\ : std_logic;
signal \quad_counter0.n19584\ : std_logic;
signal \quad_counter0.n19585\ : std_logic;
signal \quad_counter0.n19586\ : std_logic;
signal \quad_counter0.n19587\ : std_logic;
signal encoder0_position_7 : std_logic;
signal n2264 : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \quad_counter0.n19588\ : std_logic;
signal \quad_counter0.n19589\ : std_logic;
signal \quad_counter0.n19590\ : std_logic;
signal \quad_counter0.n19591\ : std_logic;
signal \quad_counter0.n19592\ : std_logic;
signal n2258 : std_logic;
signal \quad_counter0.n19593\ : std_logic;
signal n2257 : std_logic;
signal \quad_counter0.n19594\ : std_logic;
signal \quad_counter0.n19595\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \quad_counter0.n19596\ : std_logic;
signal \quad_counter0.n19597\ : std_logic;
signal \quad_counter0.n19598\ : std_logic;
signal n2252 : std_logic;
signal \quad_counter0.n19599\ : std_logic;
signal n2251 : std_logic;
signal \quad_counter0.n19600\ : std_logic;
signal \quad_counter0.n19601\ : std_logic;
signal \quad_counter0.n19602\ : std_logic;
signal \quad_counter0.n19603\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \quad_counter0.n19604\ : std_logic;
signal \quad_counter0.n19605\ : std_logic;
signal \quad_counter0.n19606\ : std_logic;
signal encoder0_position_27 : std_logic;
signal n2244 : std_logic;
signal \quad_counter0.n19607\ : std_logic;
signal \quad_counter0.n19608\ : std_logic;
signal \quad_counter0.n19609\ : std_logic;
signal n2241 : std_logic;
signal \quad_counter0.n19610\ : std_logic;
signal \quad_counter0.n19611\ : std_logic;
signal \quad_counter0.n2227\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \c0.n14474_cascade_\ : std_logic;
signal data_out_frame_9_1 : std_logic;
signal data_out_frame_8_1 : std_logic;
signal \c0.n24186\ : std_logic;
signal n2248 : std_logic;
signal n2240 : std_logic;
signal data_out_frame_7_7 : std_logic;
signal data_out_frame_5_1 : std_logic;
signal data_out_frame_8_0 : std_logic;
signal data_out_frame_7_1 : std_logic;
signal \c0.n24093\ : std_logic;
signal \c0.n5_adj_4518_cascade_\ : std_logic;
signal \c0.n23862\ : std_logic;
signal \c0.byte_transmit_counter_2\ : std_logic;
signal data_out_frame_5_7 : std_logic;
signal \c0.n24054\ : std_logic;
signal \c0.tx.r_SM_Main_0\ : std_logic;
signal \c0.tx.n7086\ : std_logic;
signal data_in_2_3 : std_logic;
signal data_in_2_1 : std_logic;
signal \c0.n13_adj_4388_cascade_\ : std_logic;
signal \c0.n23135\ : std_logic;
signal \quad_counter0.b_delay_counter_14\ : std_logic;
signal \quad_counter0.b_delay_counter_7\ : std_logic;
signal \quad_counter0.b_delay_counter_12\ : std_logic;
signal \quad_counter0.b_delay_counter_15\ : std_logic;
signal \quad_counter0.n27_adj_4200\ : std_logic;
signal \c0.n14457\ : std_logic;
signal \c0.FRAME_MATCHER_state_22\ : std_logic;
signal \c0.n14457_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_27\ : std_logic;
signal \c0.n21330\ : std_logic;
signal \c0.n30_adj_4411_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_8\ : std_logic;
signal \c0.n21344\ : std_logic;
signal \c0.n21336\ : std_logic;
signal \c0.n44_adj_4412\ : std_logic;
signal \c0.FRAME_MATCHER_state_14\ : std_logic;
signal \c0.FRAME_MATCHER_state_21\ : std_logic;
signal \c0.n21368\ : std_logic;
signal \c0.FRAME_MATCHER_state_29\ : std_logic;
signal \c0.n21326\ : std_logic;
signal \c0.n20658\ : std_logic;
signal \c0.n21152\ : std_logic;
signal \c0.n21168\ : std_logic;
signal \c0.n12542\ : std_logic;
signal \c0.n20180\ : std_logic;
signal \c0.n23260\ : std_logic;
signal \c0.n16_adj_4498_cascade_\ : std_logic;
signal \c0.n21998\ : std_logic;
signal \c0.n21852\ : std_logic;
signal \c0.n20249\ : std_logic;
signal \c0.n21210\ : std_logic;
signal \c0.n17_adj_4499\ : std_logic;
signal \c0.data_out_frame_29_7\ : std_logic;
signal \c0.data_out_frame_28_7\ : std_logic;
signal \c0.n26_adj_4359\ : std_logic;
signal data_out_frame_13_1 : std_logic;
signal data_out_frame_12_1 : std_logic;
signal \c0.n11_adj_4520\ : std_logic;
signal data_out_frame_8_3 : std_logic;
signal \c0.n11_adj_4303\ : std_logic;
signal encoder1_position_12 : std_logic;
signal data_out_frame_12_4 : std_logic;
signal encoder1_position_8 : std_logic;
signal data_out_frame_12_0 : std_logic;
signal \c0.n13079\ : std_logic;
signal \c0.n22174\ : std_logic;
signal data_in_3_5 : std_logic;
signal encoder1_position_10 : std_logic;
signal data_out_frame_12_2 : std_logic;
signal \c0.n21918\ : std_logic;
signal encoder1_position_4 : std_logic;
signal data_out_frame_13_4 : std_logic;
signal encoder1_position_2 : std_logic;
signal data_out_frame_13_2 : std_logic;
signal encoder1_position_6 : std_logic;
signal encoder1_position_7 : std_logic;
signal \c0.n21896\ : std_logic;
signal encoder1_position_26 : std_logic;
signal \c0.n20236\ : std_logic;
signal \c0.n22449\ : std_logic;
signal \c0.n22474\ : std_logic;
signal \c0.n22483\ : std_logic;
signal encoder1_position_30 : std_logic;
signal \c0.n16_adj_4321_cascade_\ : std_logic;
signal \c0.n18_adj_4322_cascade_\ : std_logic;
signal \c0.n17_adj_4323\ : std_logic;
signal \c0.n14_adj_4324\ : std_logic;
signal \c0.n22376\ : std_logic;
signal \c0.n13619\ : std_logic;
signal \c0.n13619_cascade_\ : std_logic;
signal \c0.n22412\ : std_logic;
signal \c0.n13524_cascade_\ : std_logic;
signal \c0.n10_adj_4317\ : std_logic;
signal \c0.n20328\ : std_logic;
signal encoder0_position_14 : std_logic;
signal \c0.n20328_cascade_\ : std_logic;
signal \c0.n22367\ : std_logic;
signal \c0.n22367_cascade_\ : std_logic;
signal \c0.n23569\ : std_logic;
signal n2271 : std_logic;
signal \c0.n10_adj_4331\ : std_logic;
signal \c0.n22230\ : std_logic;
signal encoder0_position_1 : std_logic;
signal \c0.n22461_cascade_\ : std_logic;
signal encoder0_position_13 : std_logic;
signal \c0.n20_adj_4318\ : std_logic;
signal n2265 : std_logic;
signal encoder0_position_6 : std_logic;
signal encoder0_position_20 : std_logic;
signal n2266 : std_logic;
signal encoder0_position_5 : std_logic;
signal \c0.n21808\ : std_logic;
signal n2250 : std_logic;
signal encoder0_position_21 : std_logic;
signal n2262 : std_logic;
signal n2260 : std_logic;
signal n2254 : std_logic;
signal \c0.n10394\ : std_logic;
signal encoder0_position_17 : std_logic;
signal encoder1_position_28 : std_logic;
signal \c0.n13338\ : std_logic;
signal data_in_2_5 : std_logic;
signal data_in_1_3 : std_logic;
signal \c0.n16_adj_4478\ : std_logic;
signal data_in_1_1 : std_logic;
signal data_in_0_1 : std_logic;
signal data_out_frame_6_5 : std_logic;
signal n2256 : std_logic;
signal encoder0_position_15 : std_logic;
signal data_in_2_0 : std_logic;
signal n2247 : std_logic;
signal n2242 : std_logic;
signal data_in_3_6 : std_logic;
signal data_in_2_6 : std_logic;
signal data_out_frame_10_1 : std_logic;
signal \c0.byte_transmit_counter_1\ : std_logic;
signal \c0.n24183\ : std_logic;
signal data_in_3_7 : std_logic;
signal data_in_2_7 : std_logic;
signal data_in_3_2 : std_logic;
signal encoder1_position_17 : std_logic;
signal data_out_frame_11_1 : std_logic;
signal \c0.n9_adj_4415_cascade_\ : std_logic;
signal n14252 : std_logic;
signal \c0.n38_adj_4387\ : std_logic;
signal \c0.tx_active\ : std_logic;
signal \c0.n22651\ : std_logic;
signal \n22661_cascade_\ : std_logic;
signal data_out_frame_7_3 : std_logic;
signal data_out_frame_6_1 : std_logic;
signal encoder0_position_0 : std_logic;
signal data_out_frame_9_0 : std_logic;
signal \c0.n21789\ : std_logic;
signal \c0.n12996_cascade_\ : std_logic;
signal \c0.n13020_cascade_\ : std_logic;
signal \c0.data_out_frame_29_7_N_1483_1_cascade_\ : std_logic;
signal \c0.n6650\ : std_logic;
signal \c0.n6650_cascade_\ : std_logic;
signal \c0.n6_adj_4270\ : std_logic;
signal \c0.n117\ : std_logic;
signal \c0.n63_adj_4301\ : std_logic;
signal \c0.n16958_cascade_\ : std_logic;
signal \c0.n63\ : std_logic;
signal \c0.n22695_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_2\ : std_logic;
signal \c0.n13_adj_4388\ : std_logic;
signal \c0.n9207\ : std_logic;
signal \c0.n14_adj_4337\ : std_logic;
signal \c0.n7_adj_4352_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_26\ : std_logic;
signal \c0.n48_cascade_\ : std_logic;
signal \c0.n45_adj_4413\ : std_logic;
signal \c0.FRAME_MATCHER_state_23\ : std_logic;
signal \c0.n14_adj_4316\ : std_logic;
signal \c0.FRAME_MATCHER_state_24\ : std_logic;
signal \c0.n21372\ : std_logic;
signal \c0.n21346\ : std_logic;
signal \c0.n21364\ : std_logic;
signal \c0.FRAME_MATCHER_state_9\ : std_logic;
signal \c0.n46\ : std_logic;
signal \c0.n20_adj_4482\ : std_logic;
signal \c0.n21_adj_4480_cascade_\ : std_logic;
signal \c0.n19_adj_4481\ : std_logic;
signal \c0.n14789\ : std_logic;
signal \c0.FRAME_MATCHER_state_18\ : std_logic;
signal \c0.FRAME_MATCHER_state_16\ : std_logic;
signal \c0.FRAME_MATCHER_state_17\ : std_logic;
signal \c0.n21682\ : std_logic;
signal \c0.FRAME_MATCHER_state_4\ : std_logic;
signal \c0.n47\ : std_logic;
signal \c0.FRAME_MATCHER_state_25\ : std_logic;
signal \c0.n21374\ : std_logic;
signal \c0.FRAME_MATCHER_state_10\ : std_logic;
signal \c0.n21348\ : std_logic;
signal \c0.FRAME_MATCHER_state_7\ : std_logic;
signal \c0.n21342\ : std_logic;
signal \c0.FRAME_MATCHER_state_11\ : std_logic;
signal \c0.n21350\ : std_logic;
signal encoder1_position_13 : std_logic;
signal data_out_frame_12_5 : std_logic;
signal \c0.n14_adj_4364\ : std_logic;
signal \c0.n13\ : std_logic;
signal \c0.n13_adj_4366_cascade_\ : std_logic;
signal \c0.n14_adj_4365\ : std_logic;
signal \c0.n14_adj_4400\ : std_logic;
signal \c0.n17600_cascade_\ : std_logic;
signal \c0.data_in_frame_10_4\ : std_logic;
signal \c0.n21908\ : std_logic;
signal count_enable_adj_4544 : std_logic;
signal n2185 : std_logic;
signal \c0.n13839\ : std_logic;
signal \c0.n22015\ : std_logic;
signal encoder0_position_29 : std_logic;
signal \c0.data_out_frame_29__7__N_856\ : std_logic;
signal \c0.n22382\ : std_logic;
signal \c0.n6_adj_4311\ : std_logic;
signal \c0.n22427\ : std_logic;
signal encoder0_position_19 : std_logic;
signal \c0.n21885\ : std_logic;
signal \c0.n22200\ : std_logic;
signal \c0.n22200_cascade_\ : std_logic;
signal \c0.n21970\ : std_logic;
signal \c0.n13705\ : std_logic;
signal n2259 : std_logic;
signal n2267 : std_logic;
signal n2261 : std_logic;
signal n2255 : std_logic;
signal encoder0_position_16 : std_logic;
signal \c0.n22408\ : std_logic;
signal encoder0_position_4 : std_logic;
signal \c0.n22227_cascade_\ : std_logic;
signal \c0.n22128\ : std_logic;
signal \c0.n10444\ : std_logic;
signal encoder1_position_20 : std_logic;
signal \c0.n6_adj_4312\ : std_logic;
signal encoder0_position_12 : std_logic;
signal \c0.n22477\ : std_logic;
signal \c0.n22477_cascade_\ : std_logic;
signal \c0.n6_adj_4333\ : std_logic;
signal n2243 : std_logic;
signal encoder0_position_28 : std_logic;
signal encoder0_position_9 : std_logic;
signal \c0.n6_adj_4315_cascade_\ : std_logic;
signal \c0.n20171\ : std_logic;
signal \c0.data_out_frame_29__7__N_847\ : std_logic;
signal \c0.data_out_frame_29__7__N_847_cascade_\ : std_logic;
signal encoder0_position_11 : std_logic;
signal \c0.n10_adj_4332\ : std_logic;
signal encoder0_position_24 : std_logic;
signal \c0.n21931\ : std_logic;
signal \c0.r_SM_Main_2_N_3755_0\ : std_logic;
signal \c0.n14322\ : std_logic;
signal \c0.n14322_cascade_\ : std_logic;
signal \c0.n14871\ : std_logic;
signal \c0.tx_transmit_N_3651\ : std_logic;
signal \c0.n23975\ : std_logic;
signal \c0.n18_adj_4403\ : std_logic;
signal \c0.n20875\ : std_logic;
signal \c0.n17602\ : std_logic;
signal \c0.n17602_cascade_\ : std_logic;
signal \c0.n8_adj_4417\ : std_logic;
signal n2245 : std_logic;
signal encoder0_position_26 : std_logic;
signal n2263 : std_logic;
signal encoder0_position_10 : std_logic;
signal data_out_frame_8_2 : std_logic;
signal n2246 : std_logic;
signal encoder0_position_25 : std_logic;
signal data_out_frame_7_6 : std_logic;
signal \c0.byte_transmit_counter_0\ : std_logic;
signal \c0.n5_adj_4350\ : std_logic;
signal control_mode_2 : std_logic;
signal encoder0_position_23 : std_logic;
signal encoder0_position_8 : std_logic;
signal \c0.n22032\ : std_logic;
signal data_in_3_0 : std_logic;
signal control_mode_5 : std_logic;
signal \c0.n23215_cascade_\ : std_logic;
signal \data_out_frame_29_7_N_1483_2\ : std_logic;
signal \c0.n6_adj_4338\ : std_logic;
signal \c0.data_out_frame_0__7__N_2568_cascade_\ : std_logic;
signal \c0.n1220_cascade_\ : std_logic;
signal \c0.n4_adj_4373\ : std_logic;
signal \c0.n5024_cascade_\ : std_logic;
signal \c0.n21773\ : std_logic;
signal \c0.n21773_cascade_\ : std_logic;
signal \c0.data_out_frame_29_7_N_1483_1\ : std_logic;
signal \c0.n4_adj_4328_cascade_\ : std_logic;
signal \c0.data_out_frame_0__7__N_2568\ : std_logic;
signal \c0.FRAME_MATCHER_state_1\ : std_logic;
signal \c0.n4_adj_4391\ : std_logic;
signal \c0.n38_adj_4390\ : std_logic;
signal \c0.n8107\ : std_logic;
signal \c0.n49\ : std_logic;
signal \c0.n50\ : std_logic;
signal \c0.n54\ : std_logic;
signal \c0.n22665\ : std_logic;
signal \c0.n3239\ : std_logic;
signal \c0.n63_adj_4293_cascade_\ : std_logic;
signal \c0.n13020\ : std_logic;
signal \c0.n4_adj_4345\ : std_logic;
signal \c0.n84_cascade_\ : std_logic;
signal \c0.n12990\ : std_logic;
signal \c0.n7_adj_4344\ : std_logic;
signal \c0.n12967\ : std_logic;
signal \c0.FRAME_MATCHER_state_0\ : std_logic;
signal \c0.n12996\ : std_logic;
signal \c0.n4_adj_4419\ : std_logic;
signal \c0.FRAME_MATCHER_state_30\ : std_logic;
signal \c0.n8_adj_4396\ : std_logic;
signal \c0.n21737_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_state_6\ : std_logic;
signal \c0.n21340\ : std_logic;
signal \c0.FRAME_MATCHER_state_19\ : std_logic;
signal \c0.n8_adj_4398\ : std_logic;
signal \c0.FRAME_MATCHER_state_5\ : std_logic;
signal \c0.n21338\ : std_logic;
signal \c0.n38_adj_4407_cascade_\ : std_logic;
signal \c0.n23836\ : std_logic;
signal \c0.n43_adj_4410_cascade_\ : std_logic;
signal \c0.n22443_cascade_\ : std_logic;
signal \c0.n21986_cascade_\ : std_logic;
signal data_in_frame_6_0 : std_logic;
signal \c0.n6_adj_4393_cascade_\ : std_logic;
signal \c0.n13086_cascade_\ : std_logic;
signal \c0.n25_adj_4408\ : std_logic;
signal \c0.n23648\ : std_logic;
signal \c0.n16_adj_4401\ : std_logic;
signal \c0.n21893\ : std_logic;
signal \c0.n44_adj_4409\ : std_logic;
signal \c0.data_in_frame_20_6\ : std_logic;
signal \n21744_cascade_\ : std_logic;
signal data_in_frame_6_3 : std_logic;
signal n2253 : std_logic;
signal \c0.n21816\ : std_logic;
signal \c0.n21740_cascade_\ : std_logic;
signal encoder0_position_18 : std_logic;
signal encoder0_position_3 : std_logic;
signal encoder0_position_31 : std_logic;
signal \c0.n21813\ : std_logic;
signal data_in_frame_6_5 : std_logic;
signal \c0.tx.n23987\ : std_logic;
signal \c0.tx.r_Clock_Count_6\ : std_logic;
signal n313 : std_logic;
signal \r_SM_Main_2_adj_4549\ : std_logic;
signal n8 : std_logic;
signal \r_Clock_Count_8\ : std_logic;
signal n2249 : std_logic;
signal count_enable : std_logic;
signal encoder0_position_22 : std_logic;
signal data_in_2_4 : std_logic;
signal data_in_1_4 : std_logic;
signal \c0.FRAME_MATCHER_rx_data_ready_prev\ : std_logic;
signal \c0.n17790_cascade_\ : std_logic;
signal \c0.n21775_cascade_\ : std_logic;
signal data_in_3_4 : std_logic;
signal control_mode_1 : std_logic;
signal control_mode_3 : std_logic;
signal control_mode_4 : std_logic;
signal control_mode_7 : std_logic;
signal \n23726_cascade_\ : std_logic;
signal control_mode_6 : std_logic;
signal \c0.n12876\ : std_logic;
signal \c0.n21022\ : std_logic;
signal \c0.n12991\ : std_logic;
signal \c0.n5024\ : std_logic;
signal \c0.n5_adj_4342_cascade_\ : std_logic;
signal \c0.n21686\ : std_logic;
signal \c0.FRAME_MATCHER_state_3\ : std_logic;
signal \c0.n21686_cascade_\ : std_logic;
signal \c0.n21334\ : std_logic;
signal \c0.n44_adj_4336\ : std_logic;
signal \c0.n1_adj_4349\ : std_logic;
signal \c0.n21734\ : std_logic;
signal \c0.n13021\ : std_logic;
signal \c0.n23965\ : std_logic;
signal \c0.n22575\ : std_logic;
signal \c0.n45_adj_4389\ : std_logic;
signal rx_data_ready : std_logic;
signal data_in_3_1 : std_logic;
signal \c0.n1\ : std_logic;
signal \c0.n19783\ : std_logic;
signal \c0.n937\ : std_logic;
signal \c0.FRAME_MATCHER_state_12\ : std_logic;
signal \c0.n21352\ : std_logic;
signal \c0.n20_adj_4327\ : std_logic;
signal \c0.n12992\ : std_logic;
signal \c0.n9668\ : std_logic;
signal \c0.n7_adj_4356\ : std_logic;
signal \c0.FRAME_MATCHER_state_28\ : std_logic;
signal \c0.n21378\ : std_logic;
signal \c0.FRAME_MATCHER_state_31\ : std_logic;
signal \c0.n21332\ : std_logic;
signal \c0.FRAME_MATCHER_state_13\ : std_logic;
signal \c0.n21354\ : std_logic;
signal \c0.FRAME_MATCHER_state_15\ : std_logic;
signal \c0.n21358\ : std_logic;
signal \c0.n21957\ : std_logic;
signal \c0.n21957_cascade_\ : std_logic;
signal \c0.n22287\ : std_logic;
signal \c0.data_in_frame_3_3\ : std_logic;
signal \c0.data_in_frame_5_4\ : std_logic;
signal \c0.n23838\ : std_logic;
signal \c0.n21902_cascade_\ : std_logic;
signal \c0.data_in_frame_3_0\ : std_logic;
signal \c0.n21902\ : std_logic;
signal \c0.data_in_frame_5_2\ : std_logic;
signal \c0.n21879_cascade_\ : std_logic;
signal \c0.data_in_frame_3_4\ : std_logic;
signal \c0.n22290\ : std_logic;
signal \c0.n22258\ : std_logic;
signal \c0.n22258_cascade_\ : std_logic;
signal \c0.n29_adj_4374\ : std_logic;
signal \c0.n27_adj_4377_cascade_\ : std_logic;
signal \c0.n14072_cascade_\ : std_logic;
signal \c0.n14072\ : std_logic;
signal \c0.n6_adj_4385_cascade_\ : std_logic;
signal \c0.n21803\ : std_logic;
signal \c0.n18_adj_4370\ : std_logic;
signal \c0.n22194\ : std_logic;
signal \c0.n21803_cascade_\ : std_logic;
signal \c0.n30_adj_4371\ : std_logic;
signal \c0.data_in_frame_0_1\ : std_logic;
signal \c0.data_in_frame_0_0\ : std_logic;
signal \c0.n13376_cascade_\ : std_logic;
signal \c0.n13376\ : std_logic;
signal data_in_frame_1_6 : std_logic;
signal data_in_frame_6_2 : std_logic;
signal \c0.n13386_cascade_\ : std_logic;
signal \c0.data_in_frame_4_4\ : std_logic;
signal \c0.n22261\ : std_logic;
signal \c0.data_in_frame_2_1\ : std_logic;
signal \c0.n22261_cascade_\ : std_logic;
signal \c0.n22320\ : std_logic;
signal \c0.n28_adj_4372\ : std_logic;
signal \c0.data_in_frame_3_6\ : std_logic;
signal \c0.data_in_frame_4_1\ : std_logic;
signal \c0.n22218\ : std_logic;
signal \c0.n21928_cascade_\ : std_logic;
signal \c0.data_in_frame_2_3\ : std_logic;
signal \c0.n21791\ : std_logic;
signal \c0.n21882_cascade_\ : std_logic;
signal \c0.data_out_frame_0__7__N_2744\ : std_logic;
signal \c0.data_out_frame_0__7__N_2744_cascade_\ : std_logic;
signal \c0.n6_adj_4272_cascade_\ : std_logic;
signal \c0.data_in_frame_3_7\ : std_logic;
signal \c0.data_in_frame_4_7\ : std_logic;
signal \c0.data_in_frame_5_1\ : std_logic;
signal \c0.n21992\ : std_logic;
signal \c0.data_in_frame_2_2\ : std_logic;
signal data_in_frame_1_7 : std_logic;
signal \c0.n39_adj_4406\ : std_logic;
signal data_in_frame_6_7 : std_logic;
signal \c0.n21882\ : std_logic;
signal \c0.n21928\ : std_logic;
signal \c0.n14037_cascade_\ : std_logic;
signal \c0.n6_adj_4369\ : std_logic;
signal \c0.n5_adj_4368\ : std_logic;
signal \c0.data_out_frame_29__7__N_1474\ : std_logic;
signal data_in_frame_6_6 : std_logic;
signal \c0.data_in_frame_0_2\ : std_logic;
signal \c0.data_in_frame_2_4\ : std_logic;
signal \c0.data_in_frame_5_0\ : std_logic;
signal \c0.data_in_frame_2_0\ : std_logic;
signal data_in_frame_6_1 : std_logic;
signal \n4_cascade_\ : std_logic;
signal \c0.data_in_frame_4_6\ : std_logic;
signal n4 : std_logic;
signal \c0.n21758_cascade_\ : std_logic;
signal \c0.n17790\ : std_logic;
signal data_in_frame_1_0 : std_logic;
signal n23726 : std_logic;
signal control_mode_0 : std_logic;
signal \c0.data_in_frame_29_4\ : std_logic;
signal \c0.n10_adj_4286_cascade_\ : std_logic;
signal \c0.data_in_frame_28_2\ : std_logic;
signal \c0.data_in_frame_29_0\ : std_logic;
signal \c0.n17600\ : std_logic;
signal \c0.n19_cascade_\ : std_logic;
signal \c0.n23389\ : std_logic;
signal \c0.n32_adj_4295_cascade_\ : std_logic;
signal \c0.n23523\ : std_logic;
signal \c0.n34\ : std_logic;
signal \c0.data_in_frame_29_2\ : std_logic;
signal \c0.data_in_frame_29_1\ : std_logic;
signal \c0.n23388_cascade_\ : std_logic;
signal \c0.n30_adj_4299\ : std_logic;
signal \c0.n15_adj_4376_cascade_\ : std_logic;
signal \c0.n17_adj_4378\ : std_logic;
signal \c0.n18_adj_4379_cascade_\ : std_logic;
signal \c0.n27_adj_4383\ : std_logic;
signal \c0.n30_adj_4380_cascade_\ : std_logic;
signal \c0.n28_adj_4381\ : std_logic;
signal \c0.n13000\ : std_logic;
signal data_in_frame_22_1 : std_logic;
signal \c0.rx.n22611_cascade_\ : std_logic;
signal \c0.rx.n8_cascade_\ : std_logic;
signal \c0.n29_adj_4382\ : std_logic;
signal \c0.n161\ : std_logic;
signal \bfn_19_1_0_\ : std_logic;
signal \c0.n3\ : std_logic;
signal \c0.n19442\ : std_logic;
signal \c0.n19442_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19442_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19442_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19442_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19442_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19442_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19442_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_2_0_\ : std_logic;
signal \c0.n19443\ : std_logic;
signal \c0.n19443_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19443_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19443_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19443_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19443_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19443_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19443_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_3_0_\ : std_logic;
signal \c0.n19444\ : std_logic;
signal \c0.n19444_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19444_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19444_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19444_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19444_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19444_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19444_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_4_0_\ : std_logic;
signal \c0.n19445\ : std_logic;
signal \c0.n19445_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19445_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19445_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19445_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19445_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19445_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19445_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_4\ : std_logic;
signal \bfn_19_5_0_\ : std_logic;
signal \c0.n3_adj_4470\ : std_logic;
signal \c0.n19446\ : std_logic;
signal \c0.n19446_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19446_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19446_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19446_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19446_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19446_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19446_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_6_0_\ : std_logic;
signal \c0.n3_adj_4468\ : std_logic;
signal \c0.n19447\ : std_logic;
signal \c0.n19447_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19447_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19447_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19447_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19447_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19447_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19447_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_7_0_\ : std_logic;
signal \c0.n3_adj_4467\ : std_logic;
signal \c0.n19448\ : std_logic;
signal \c0.n19448_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19448_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19448_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19448_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19448_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19448_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19448_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_7\ : std_logic;
signal \bfn_19_8_0_\ : std_logic;
signal \c0.n3_adj_4465\ : std_logic;
signal \c0.n19449\ : std_logic;
signal \c0.n19449_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19449_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19449_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19449_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19449_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19449_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19449_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_8\ : std_logic;
signal \bfn_19_9_0_\ : std_logic;
signal \c0.n3_adj_4463\ : std_logic;
signal \c0.n19450\ : std_logic;
signal \c0.n19450_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19450_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19450_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19450_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19450_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19450_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19450_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_9\ : std_logic;
signal \bfn_19_10_0_\ : std_logic;
signal \c0.n3_adj_4462\ : std_logic;
signal \c0.n19451\ : std_logic;
signal \c0.n19451_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19451_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19451_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19451_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19451_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19451_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19451_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_11_0_\ : std_logic;
signal \c0.n19452\ : std_logic;
signal \c0.n19452_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19452_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19452_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19452_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19452_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19452_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19452_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_11\ : std_logic;
signal \bfn_19_12_0_\ : std_logic;
signal \c0.n3_adj_4458\ : std_logic;
signal \c0.n19453\ : std_logic;
signal \c0.n19453_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19453_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19453_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19453_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19453_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19453_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19453_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_12\ : std_logic;
signal \bfn_19_13_0_\ : std_logic;
signal \c0.n3_adj_4456\ : std_logic;
signal \c0.n19454\ : std_logic;
signal \c0.n19454_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19454_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19454_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19454_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19454_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19454_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19454_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_14_0_\ : std_logic;
signal \c0.n19455\ : std_logic;
signal \c0.n19455_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19455_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19455_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19455_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19455_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19455_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19455_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_14\ : std_logic;
signal \bfn_19_15_0_\ : std_logic;
signal \c0.n3_adj_4453\ : std_logic;
signal \c0.n19456\ : std_logic;
signal \c0.n19456_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19456_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19456_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19456_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19456_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19456_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19456_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_16_0_\ : std_logic;
signal \c0.n19457\ : std_logic;
signal \c0.n19457_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19457_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19457_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19457_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19457_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19457_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19457_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_17_0_\ : std_logic;
signal \c0.n3_adj_4450\ : std_logic;
signal \c0.n19458\ : std_logic;
signal \c0.n19458_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19458_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19458_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19458_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19458_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19458_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19458_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_17\ : std_logic;
signal \bfn_19_18_0_\ : std_logic;
signal \c0.n3_adj_4448\ : std_logic;
signal \c0.n19459\ : std_logic;
signal \c0.n19459_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19459_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19459_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19459_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19459_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19459_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19459_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_18\ : std_logic;
signal \bfn_19_19_0_\ : std_logic;
signal \c0.n3_adj_4446\ : std_logic;
signal \c0.n19460\ : std_logic;
signal \c0.n19460_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19460_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19460_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19460_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19460_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19460_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19460_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_19\ : std_logic;
signal \bfn_19_20_0_\ : std_logic;
signal \c0.n3_adj_4444\ : std_logic;
signal \c0.n19461\ : std_logic;
signal \c0.n19461_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19461_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19461_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19461_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19461_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19461_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19461_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_21_0_\ : std_logic;
signal \c0.n19462\ : std_logic;
signal \c0.n19462_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19462_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19462_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19462_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19462_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19462_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19462_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_21\ : std_logic;
signal \bfn_19_22_0_\ : std_logic;
signal \c0.n3_adj_4440\ : std_logic;
signal \c0.n19463\ : std_logic;
signal \c0.n19463_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19463_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19463_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19463_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19463_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19463_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19463_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_22\ : std_logic;
signal \bfn_19_23_0_\ : std_logic;
signal \c0.n3_adj_4438\ : std_logic;
signal \c0.n19464\ : std_logic;
signal \c0.n19464_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19464_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19464_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19464_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19464_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19464_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19464_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_23\ : std_logic;
signal \bfn_19_24_0_\ : std_logic;
signal \c0.n3_adj_4436\ : std_logic;
signal \c0.n19465\ : std_logic;
signal \c0.n19465_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19465_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19465_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19465_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19465_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19465_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19465_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_24\ : std_logic;
signal \bfn_19_25_0_\ : std_logic;
signal \c0.n3_adj_4435\ : std_logic;
signal \c0.n19466\ : std_logic;
signal \c0.n19466_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19466_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19466_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19466_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19466_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19466_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19466_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_25\ : std_logic;
signal \bfn_19_26_0_\ : std_logic;
signal \c0.n3_adj_4434\ : std_logic;
signal \c0.n19467\ : std_logic;
signal \c0.n19467_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19467_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19467_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19467_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19467_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19467_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19467_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_26\ : std_logic;
signal \bfn_19_27_0_\ : std_logic;
signal \c0.n3_adj_4433\ : std_logic;
signal \c0.n19468\ : std_logic;
signal \c0.n19468_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19468_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19468_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19468_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19468_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19468_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19468_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_27\ : std_logic;
signal \bfn_19_28_0_\ : std_logic;
signal \c0.n3_adj_4432\ : std_logic;
signal \c0.n19469\ : std_logic;
signal \c0.n19469_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19469_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19469_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19469_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19469_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19469_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19469_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_29_0_\ : std_logic;
signal \c0.n19470\ : std_logic;
signal \c0.n19470_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19470_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19470_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19470_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19470_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19470_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19470_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_29\ : std_logic;
signal \bfn_19_30_0_\ : std_logic;
signal \c0.n3_adj_4428\ : std_logic;
signal \c0.n19471\ : std_logic;
signal \c0.n19471_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19471_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19471_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19471_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19471_THRU_CRY_4_THRU_CO\ : std_logic;
signal \c0.n19471_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19471_THRU_CRY_6_THRU_CO\ : std_logic;
signal \c0.FRAME_MATCHER_i_30\ : std_logic;
signal \bfn_19_31_0_\ : std_logic;
signal \c0.n3_adj_4426\ : std_logic;
signal \c0.n19472\ : std_logic;
signal \c0.n19472_THRU_CRY_0_THRU_CO\ : std_logic;
signal \c0.n19472_THRU_CRY_1_THRU_CO\ : std_logic;
signal \c0.n19472_THRU_CRY_2_THRU_CO\ : std_logic;
signal \c0.n19472_THRU_CRY_3_THRU_CO\ : std_logic;
signal \c0.n19472_THRU_CRY_4_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \c0.n19472_THRU_CRY_5_THRU_CO\ : std_logic;
signal \c0.n19472_THRU_CRY_6_THRU_CO\ : std_logic;
signal \bfn_19_32_0_\ : std_logic;
signal \c0.FRAME_MATCHER_i_31\ : std_logic;
signal \c0.n3_adj_4421\ : std_logic;
signal \c0.n3_adj_4475\ : std_logic;
signal \c0.FRAME_MATCHER_i_3\ : std_logic;
signal \c0.n3_adj_4472\ : std_logic;
signal \c0.n3_adj_4474\ : std_logic;
signal \c0.FRAME_MATCHER_i_5\ : std_logic;
signal \c0.FRAME_MATCHER_i_6\ : std_logic;
signal \c0.n11_adj_4326\ : std_logic;
signal \c0.n10_adj_4399\ : std_logic;
signal \c0.n13033\ : std_logic;
signal \c0.data_in_frame_2_7\ : std_logic;
signal \c0.data_in_frame_0_7\ : std_logic;
signal \c0.data_in_frame_8_4\ : std_logic;
signal \c0.n21861_cascade_\ : std_logic;
signal \c0.n6_adj_4258\ : std_logic;
signal \c0.data_in_frame_9_5\ : std_logic;
signal \c0.n8_adj_4254_cascade_\ : std_logic;
signal \c0.n4_adj_4255\ : std_logic;
signal \c0.data_in_frame_5_5\ : std_logic;
signal \c0.data_in_frame_3_1\ : std_logic;
signal \c0.data_in_frame_3_2\ : std_logic;
signal \c0.n6_adj_4395\ : std_logic;
signal data_in_frame_1_1 : std_logic;
signal data_in_frame_1_5 : std_logic;
signal \c0.n21986\ : std_logic;
signal \c0.n13848_cascade_\ : std_logic;
signal \c0.n13_adj_4405\ : std_logic;
signal \c0.data_in_frame_2_5\ : std_logic;
signal \c0.data_in_frame_0_3\ : std_logic;
signal \c0.n13398\ : std_logic;
signal data_in_frame_1_3 : std_logic;
signal \c0.data_in_frame_3_5\ : std_logic;
signal \c0.n13398_cascade_\ : std_logic;
signal \c0.n13852\ : std_logic;
signal \c0.n21794\ : std_logic;
signal \c0.data_in_frame_8_2\ : std_logic;
signal \c0.n21794_cascade_\ : std_logic;
signal \c0.data_in_frame_5_7\ : std_logic;
signal \c0.n6_adj_4257_cascade_\ : std_logic;
signal \c0.n21825\ : std_logic;
signal \c0.n13771_cascade_\ : std_logic;
signal \c0.n22239\ : std_logic;
signal \c0.n4_cascade_\ : std_logic;
signal \c0.n37\ : std_logic;
signal \c0.n6_adj_4220\ : std_logic;
signal \c0.data_in_frame_8_3\ : std_logic;
signal \c0.n13652\ : std_logic;
signal \c0.n13771\ : std_logic;
signal \c0.data_in_frame_10_3\ : std_logic;
signal \c0.n21964\ : std_logic;
signal \c0.n22280\ : std_logic;
signal \c0.n21964_cascade_\ : std_logic;
signal \c0.n14113\ : std_logic;
signal \c0.n6_adj_4241\ : std_logic;
signal \c0.n13086\ : std_logic;
signal \c0.data_in_frame_8_5\ : std_logic;
signal \c0.n22415_cascade_\ : std_logic;
signal \c0.data_in_frame_10_5\ : std_logic;
signal \c0.n35\ : std_logic;
signal n21744 : std_logic;
signal \c0.n6_adj_4386\ : std_logic;
signal \c0.data_in_frame_4_3\ : std_logic;
signal data_in_frame_6_4 : std_logic;
signal \c0.data_in_frame_4_2\ : std_logic;
signal \FRAME_MATCHER_state_31_N_2976_2\ : std_logic;
signal n22661 : std_logic;
signal encoder0_position_30 : std_logic;
signal data_out_frame_6_6 : std_logic;
signal \c0.n13697\ : std_logic;
signal \c0.n22440_cascade_\ : std_logic;
signal \c0.data_in_frame_10_7\ : std_logic;
signal \c0.n10_adj_4229_cascade_\ : std_logic;
signal \c0.n5943_cascade_\ : std_logic;
signal \c0.n22081_cascade_\ : std_logic;
signal \c0.n22349_cascade_\ : std_logic;
signal \c0.n21858_cascade_\ : std_logic;
signal \c0.FRAME_MATCHER_i_16\ : std_logic;
signal \c0.n16_adj_4375\ : std_logic;
signal \c0.FRAME_MATCHER_i_13\ : std_logic;
signal \c0.n3_adj_4454\ : std_logic;
signal \c0.FRAME_MATCHER_i_15\ : std_logic;
signal \c0.n3_adj_4452\ : std_logic;
signal \c0.FRAME_MATCHER_i_20\ : std_logic;
signal \c0.n3_adj_4442\ : std_logic;
signal \c0.data_in_frame_28_1\ : std_logic;
signal \c0.n21870_cascade_\ : std_logic;
signal \c0.data_in_frame_21_3\ : std_logic;
signal \c0.data_in_frame_23_5\ : std_logic;
signal \c0.data_in_frame_23_4\ : std_logic;
signal \c0.n10_adj_4287_cascade_\ : std_logic;
signal \c0.n22_adj_4298\ : std_logic;
signal \c0.n13266\ : std_logic;
signal \c0.data_in_frame_29_7\ : std_logic;
signal \c0.n21233_cascade_\ : std_logic;
signal \c0.n23506\ : std_logic;
signal \c0.data_in_frame_27_1\ : std_logic;
signal \c0.FRAME_MATCHER_i_10\ : std_logic;
signal \c0.n3_adj_4460\ : std_logic;
signal n18678 : std_logic;
signal \c0.rx.n18655_cascade_\ : std_logic;
signal \c0.rx.n21704_cascade_\ : std_logic;
signal \c0.rx.n22573_cascade_\ : std_logic;
signal \c0.rx.n12_cascade_\ : std_logic;
signal \bfn_20_24_0_\ : std_logic;
signal \c0.rx.r_Clock_Count_1\ : std_logic;
signal \c0.rx.n19533\ : std_logic;
signal \c0.rx.r_Clock_Count_2\ : std_logic;
signal \c0.rx.n19534\ : std_logic;
signal \c0.rx.r_Clock_Count_3\ : std_logic;
signal \c0.rx.n19535\ : std_logic;
signal \c0.rx.n19536\ : std_logic;
signal \c0.rx.n19537\ : std_logic;
signal \c0.rx.n19538\ : std_logic;
signal \c0.rx.n19539\ : std_logic;
signal \c0.rx.n14391\ : std_logic;
signal \c0.rx.n17411\ : std_logic;
signal \c0.data_out_frame_29_7_N_1483_0\ : std_logic;
signal \c0.n1220\ : std_logic;
signal \c0.FRAME_MATCHER_i_28\ : std_logic;
signal \c0.n31_adj_4271\ : std_logic;
signal \c0.n3_adj_4430\ : std_logic;
signal \c0.data_in_frame_7_4\ : std_logic;
signal \c0.n13555_cascade_\ : std_logic;
signal \c0.n13555\ : std_logic;
signal \c0.n22043_cascade_\ : std_logic;
signal \c0.data_in_frame_2_6\ : std_logic;
signal \c0.data_in_frame_0_4\ : std_logic;
signal \c0.n10_adj_4363\ : std_logic;
signal \c0.n22283\ : std_logic;
signal \c0.n13488_cascade_\ : std_logic;
signal \c0.n13180\ : std_logic;
signal \c0.data_in_frame_0_5\ : std_logic;
signal \c0.data_in_frame_0_6\ : std_logic;
signal \c0.n23827\ : std_logic;
signal \c0.data_in_frame_5_3\ : std_logic;
signal \c0.data_in_frame_7_5\ : std_logic;
signal \c0.n12484\ : std_logic;
signal \c0.n20368_cascade_\ : std_logic;
signal \c0.data_in_frame_10_1\ : std_logic;
signal \c0.n22133_cascade_\ : std_logic;
signal \c0.n21925\ : std_logic;
signal \c0.n20927_cascade_\ : std_logic;
signal \c0.n22133\ : std_logic;
signal \c0.n36\ : std_logic;
signal data_in_frame_1_2 : std_logic;
signal \c0.n22334\ : std_logic;
signal \c0.n22334_cascade_\ : std_logic;
signal \c0.n22051\ : std_logic;
signal \c0.n15_adj_4404\ : std_logic;
signal \c0.data_in_frame_8_0\ : std_logic;
signal \c0.data_in_frame_7_7\ : std_logic;
signal \c0.n6_adj_4259\ : std_logic;
signal \c0.n39_adj_4263\ : std_logic;
signal \c0.n40_adj_4261\ : std_logic;
signal \c0.n22060_cascade_\ : std_logic;
signal \c0.n44_adj_4262\ : std_logic;
signal \c0.n11_adj_4266_cascade_\ : std_logic;
signal \c0.n13425\ : std_logic;
signal \c0.n22842_cascade_\ : std_logic;
signal \c0.data_in_frame_5_6\ : std_logic;
signal \c0.n22245\ : std_logic;
signal \c0.n22379\ : std_logic;
signal \c0.n38_adj_4260\ : std_logic;
signal \c0.n6_adj_4256\ : std_logic;
signal \c0.data_in_frame_7_3\ : std_logic;
signal \c0.n13488\ : std_logic;
signal \c0.n22139_cascade_\ : std_logic;
signal \c0.data_in_frame_9_0\ : std_logic;
signal \c0.n13605\ : std_logic;
signal \c0.n13043\ : std_logic;
signal \c0.data_in_frame_8_6\ : std_logic;
signal \c0.n21822_cascade_\ : std_logic;
signal \c0.n22443\ : std_logic;
signal \c0.n10_adj_4242_cascade_\ : std_logic;
signal \c0.data_in_frame_8_1\ : std_logic;
signal \c0.data_in_frame_16_6\ : std_logic;
signal \c0.n13786_cascade_\ : std_logic;
signal \c0.n21170\ : std_logic;
signal \c0.n13974\ : std_logic;
signal \c0.data_in_frame_10_2\ : std_logic;
signal \c0.n20402_cascade_\ : std_logic;
signal \c0.data_in_frame_9_6\ : std_logic;
signal \c0.data_in_frame_9_4\ : std_logic;
signal \c0.n21873\ : std_logic;
signal \c0.n13287\ : std_logic;
signal \c0.n13190\ : std_logic;
signal \c0.n18_adj_4222_cascade_\ : std_logic;
signal \c0.n22270\ : std_logic;
signal \c0.n6_adj_4221\ : std_logic;
signal \c0.n22308\ : std_logic;
signal \c0.n22003_cascade_\ : std_logic;
signal \c0.n5943\ : std_logic;
signal \c0.n6221_cascade_\ : std_logic;
signal \c0.n22003\ : std_logic;
signal \c0.data_in_frame_20_1\ : std_logic;
signal \c0.n6_adj_4226_cascade_\ : std_logic;
signal \c0.n23615_cascade_\ : std_logic;
signal \c0.n22100_cascade_\ : std_logic;
signal \c0.n22081\ : std_logic;
signal \c0.n6_adj_4224\ : std_logic;
signal \c0.n21737\ : std_logic;
signal \c0.n6_adj_4353\ : std_logic;
signal \c0.n5_adj_4342\ : std_logic;
signal \c0.FRAME_MATCHER_state_20\ : std_logic;
signal \c0.n21366\ : std_logic;
signal \c0.n21855\ : std_logic;
signal encoder0_position_2 : std_logic;
signal \c0.n22248\ : std_logic;
signal \c0.n13379\ : std_logic;
signal \c0.data_in_frame_20_7\ : std_logic;
signal \c0.n28_cascade_\ : std_logic;
signal \c0.n23640_cascade_\ : std_logic;
signal \c0.n22305_cascade_\ : std_logic;
signal \c0.data_in_frame_21_1\ : std_logic;
signal \c0.n23640\ : std_logic;
signal \c0.n22305\ : std_logic;
signal \c0.n6_adj_4219_cascade_\ : std_logic;
signal \c0.data_in_frame_21_2\ : std_logic;
signal \c0.n22197\ : std_logic;
signal \c0.n21949_cascade_\ : std_logic;
signal \c0.n20137\ : std_logic;
signal \c0.n22157_cascade_\ : std_logic;
signal \c0.n20846\ : std_logic;
signal \c0.n20846_cascade_\ : std_logic;
signal \c0.data_in_frame_25_4\ : std_logic;
signal \c0.data_in_frame_25_2\ : std_logic;
signal \c0.data_in_frame_25_3\ : std_logic;
signal \c0.data_in_frame_25_5\ : std_logic;
signal \c0.n22370\ : std_logic;
signal \c0.n12_adj_4491\ : std_logic;
signal \c0.n23009\ : std_logic;
signal \c0.n22370_cascade_\ : std_logic;
signal \c0.n23356\ : std_logic;
signal \c0.n13761\ : std_logic;
signal \c0.n22145\ : std_logic;
signal \c0.n21949\ : std_logic;
signal \c0.n22145_cascade_\ : std_logic;
signal \c0.n10_adj_4297\ : std_logic;
signal \c0.n23335_cascade_\ : std_logic;
signal \c0.n21_adj_4300\ : std_logic;
signal \c0.data_in_frame_29_3\ : std_logic;
signal \c0.data_in_frame_28_0\ : std_logic;
signal \c0.n6404\ : std_logic;
signal \c0.n21834\ : std_logic;
signal \c0.n22040\ : std_logic;
signal \c0.n22040_cascade_\ : std_logic;
signal \c0.n21208\ : std_logic;
signal \c0.n21099\ : std_logic;
signal \c0.n22119\ : std_logic;
signal \c0.n21099_cascade_\ : std_logic;
signal \c0.n21160\ : std_logic;
signal \c0.data_in_frame_29_6\ : std_logic;
signal \c0.n63_adj_4293\ : std_logic;
signal \c0.n22148_cascade_\ : std_logic;
signal \c0.n21233\ : std_logic;
signal \c0.n26_adj_4294\ : std_logic;
signal \c0.rx.n12862_cascade_\ : std_logic;
signal \c0.rx.r_Clock_Count_7\ : std_logic;
signal \c0.rx.r_Clock_Count_5\ : std_logic;
signal \c0.rx.r_Clock_Count_6\ : std_logic;
signal \c0.rx.n80_cascade_\ : std_logic;
signal \r_SM_Main_2_N_3681_2_cascade_\ : std_logic;
signal n14283 : std_logic;
signal \c0.rx.r_Clock_Count_4\ : std_logic;
signal \c0.rx.n18655\ : std_logic;
signal \c0.rx.r_Clock_Count_0\ : std_logic;
signal \c0.rx.n80\ : std_logic;
signal \c0.rx.n21783\ : std_logic;
signal \c0.rx.r_Rx_Data_R\ : std_logic;
signal \c0.data_in_frame_12_6\ : std_logic;
signal \c0.data_in_frame_15_3\ : std_logic;
signal \c0.n20927\ : std_logic;
signal \c0.n22060\ : std_logic;
signal \c0.n6_adj_4244_cascade_\ : std_logic;
signal \c0.n21097\ : std_logic;
signal \c0.n20240_cascade_\ : std_logic;
signal \c0.data_in_frame_15_0\ : std_logic;
signal \c0.n22385_cascade_\ : std_logic;
signal data_in_frame_14_5 : std_logic;
signal data_in_frame_14_3 : std_logic;
signal \c0.data_in_frame_4_0\ : std_logic;
signal data_in_frame_1_4 : std_logic;
signal \c0.n21797\ : std_logic;
signal \c0.n13237\ : std_logic;
signal \c0.data_in_frame_7_6\ : std_logic;
signal \c0.data_in_frame_10_0\ : std_logic;
signal \c0.n10_adj_4245_cascade_\ : std_logic;
signal \c0.n13099\ : std_logic;
signal \c0.data_in_frame_9_1\ : std_logic;
signal \c0.n14037\ : std_logic;
signal \c0.n22233\ : std_logic;
signal \c0.data_in_frame_11_3\ : std_logic;
signal \c0.n10_adj_4274\ : std_logic;
signal \c0.n22108\ : std_logic;
signal \c0.n4_adj_4240_cascade_\ : std_logic;
signal \c0.data_in_frame_7_1\ : std_logic;
signal \c0.n6_adj_4273\ : std_logic;
signal \c0.n22139\ : std_logic;
signal \c0.n6_adj_4243\ : std_logic;
signal \c0.n13861\ : std_logic;
signal \c0.n5813_cascade_\ : std_logic;
signal \c0.n21967\ : std_logic;
signal \c0.n20222_cascade_\ : std_logic;
signal \c0.n13677\ : std_logic;
signal \c0.n28_adj_4232_cascade_\ : std_logic;
signal \c0.n32_cascade_\ : std_logic;
signal \c0.n29_adj_4234\ : std_logic;
signal \c0.n13681\ : std_logic;
signal \c0.n21238_cascade_\ : std_logic;
signal \c0.n21989\ : std_logic;
signal \c0.n21238\ : std_logic;
signal \c0.n22430\ : std_logic;
signal \c0.n5810\ : std_logic;
signal \c0.n13719_cascade_\ : std_logic;
signal \c0.n22221\ : std_logic;
signal \c0.n13786\ : std_logic;
signal data_in_frame_14_6 : std_logic;
signal data_in_frame_14_7 : std_logic;
signal \c0.n5996\ : std_logic;
signal \c0.n7_adj_4235\ : std_logic;
signal \c0.n8_adj_4236\ : std_logic;
signal \c0.n20203_cascade_\ : std_logic;
signal \c0.n21120\ : std_logic;
signal \c0.data_in_frame_15_2\ : std_logic;
signal \c0.n22242\ : std_logic;
signal \c0.n20402\ : std_logic;
signal \c0.n20196\ : std_logic;
signal \c0.n22100\ : std_logic;
signal \c0.n21054_cascade_\ : std_logic;
signal \c0.n21043\ : std_logic;
signal \c0.data_in_frame_17_3\ : std_logic;
signal \c0.data_in_frame_17_4\ : std_logic;
signal \c0.n22480\ : std_logic;
signal \c0.data_in_frame_17_5\ : std_logic;
signal \c0.n13719\ : std_logic;
signal \c0.n18\ : std_logic;
signal \c0.n22349\ : std_logic;
signal \c0.n30\ : std_logic;
signal \c0.n22\ : std_logic;
signal \c0.n22355\ : std_logic;
signal \c0.n23062_cascade_\ : std_logic;
signal \c0.data_in_frame_21_0\ : std_logic;
signal \c0.n23062\ : std_logic;
signal \c0.n8\ : std_logic;
signal \c0.n27\ : std_logic;
signal \c0.n22296\ : std_logic;
signal \c0.n21831\ : std_logic;
signal \c0.data_in_frame_17_0\ : std_logic;
signal \c0.n16_adj_4223_cascade_\ : std_logic;
signal \c0.n17\ : std_logic;
signal \c0.n21187\ : std_logic;
signal \c0.n22211_cascade_\ : std_logic;
signal \c0.n21140\ : std_logic;
signal \c0.n22311\ : std_logic;
signal \c0.n22211\ : std_logic;
signal \c0.n23298\ : std_logic;
signal \c0.n7\ : std_logic;
signal \c0.n23298_cascade_\ : std_logic;
signal \c0.n45_adj_4486\ : std_logic;
signal \c0.data_in_frame_27_4\ : std_logic;
signal \c0.n52_cascade_\ : std_logic;
signal \c0.n13872\ : std_logic;
signal \c0.n12420\ : std_logic;
signal \c0.n23615\ : std_logic;
signal \c0.n44_adj_4490\ : std_logic;
signal \c0.n48_adj_4485_cascade_\ : std_logic;
signal \c0.n12_adj_4290\ : std_logic;
signal \c0.data_in_frame_25_1\ : std_logic;
signal \c0.n49_adj_4488\ : std_logic;
signal \c0.n55\ : std_logic;
signal \c0.n53\ : std_logic;
signal \c0.n23416\ : std_logic;
signal \c0.n23416_cascade_\ : std_logic;
signal \c0.n12_adj_4296\ : std_logic;
signal \c0.data_in_frame_27_2\ : std_logic;
signal \c0.n36_adj_4489\ : std_logic;
signal \c0.data_in_frame_19_2\ : std_logic;
signal \c0.n6221\ : std_logic;
signal \c0.n21037\ : std_logic;
signal \c0.data_in_frame_23_6\ : std_logic;
signal \c0.n21037_cascade_\ : std_logic;
signal \c0.data_in_frame_19_4\ : std_logic;
signal \c0.n13282\ : std_logic;
signal \c0.n20370\ : std_logic;
signal \c0.data_in_frame_29_5\ : std_logic;
signal \c0.n22157\ : std_logic;
signal \c0.data_in_frame_27_3\ : std_logic;
signal \c0.n22719\ : std_logic;
signal \c0.n8_adj_4291_cascade_\ : std_logic;
signal \c0.n22148\ : std_logic;
signal \c0.n23811\ : std_logic;
signal n12977 : std_logic;
signal \c0.rx.n21704\ : std_logic;
signal \n14436_cascade_\ : std_logic;
signal \c0.rx.n12862\ : std_logic;
signal n19619 : std_logic;
signal \r_Bit_Index_2\ : std_logic;
signal \n91_cascade_\ : std_logic;
signal \r_SM_Main_2_N_3681_2\ : std_logic;
signal \r_SM_Main_2\ : std_logic;
signal \r_SM_Main_1\ : std_logic;
signal \c0.rx.n14_cascade_\ : std_logic;
signal \c0.rx.n36\ : std_logic;
signal \r_SM_Main_0\ : std_logic;
signal \n21755_cascade_\ : std_logic;
signal data_in_frame_14_1 : std_logic;
signal \c0.FRAME_MATCHER_i_0\ : std_logic;
signal \c0.FRAME_MATCHER_i_1\ : std_logic;
signal \c0.FRAME_MATCHER_i_2\ : std_logic;
signal \c0.n22043\ : std_logic;
signal \c0.data_in_frame_9_7\ : std_logic;
signal \c0.n22471\ : std_logic;
signal \c0.data_in_frame_16_4\ : std_logic;
signal \c0.n20240\ : std_logic;
signal \c0.n22446\ : std_logic;
signal \c0.n22328\ : std_logic;
signal \c0.n22446_cascade_\ : std_logic;
signal \c0.n22424\ : std_logic;
signal \c0.n30_adj_4233\ : std_logic;
signal data_in_frame_14_2 : std_logic;
signal \c0.n22340\ : std_logic;
signal n21755 : std_logic;
signal data_in_frame_14_4 : std_logic;
signal \c0.n15_adj_4269\ : std_logic;
signal \c0.n22464_cascade_\ : std_logic;
signal \c0.n22415\ : std_logic;
signal \c0.n13728\ : std_logic;
signal \c0.n14053\ : std_logic;
signal \c0.data_in_frame_18_1\ : std_logic;
signal \c0.n14053_cascade_\ : std_logic;
signal \c0.data_in_frame_17_7\ : std_logic;
signal \c0.n23586_cascade_\ : std_logic;
signal \c0.data_in_frame_9_3\ : std_logic;
signal \c0.n13210_cascade_\ : std_logic;
signal \c0.data_in_frame_8_7\ : std_logic;
signal \c0.n21822\ : std_logic;
signal \c0.n7_adj_4277_cascade_\ : std_logic;
signal \c0.data_in_frame_11_5\ : std_logic;
signal \c0.n10_adj_4264_cascade_\ : std_logic;
signal \c0.n16_adj_4265\ : std_logic;
signal \c0.data_in_frame_11_6\ : std_logic;
signal \c0.data_in_frame_11_2\ : std_logic;
signal \c0.n20135\ : std_logic;
signal \c0.n22464\ : std_logic;
signal \c0.n21867\ : std_logic;
signal \c0.n6_adj_4225\ : std_logic;
signal \c0.n21982\ : std_logic;
signal data_in_frame_14_0 : std_logic;
signal \c0.n13865\ : std_logic;
signal \c0.data_in_frame_15_6\ : std_logic;
signal \c0.n4_adj_4240\ : std_logic;
signal \c0.n22352_cascade_\ : std_logic;
signal \c0.n22000_cascade_\ : std_logic;
signal \c0.n31\ : std_logic;
signal \c0.data_in_frame_15_7\ : std_logic;
signal \c0.data_in_frame_18_2\ : std_logic;
signal \c0.n22000\ : std_logic;
signal \c0.n12_cascade_\ : std_logic;
signal \c0.n10_adj_4239\ : std_logic;
signal \c0.data_in_frame_18_0\ : std_logic;
signal \c0.n14_adj_4238\ : std_logic;
signal \c0.n22352\ : std_logic;
signal \c0.data_in_frame_18_4\ : std_logic;
signal \c0.n13598\ : std_logic;
signal \c0.n20374\ : std_logic;
signal \c0.data_in_frame_16_5\ : std_logic;
signal \c0.data_in_frame_16_3\ : std_logic;
signal \c0.data_in_frame_16_2\ : std_logic;
signal \c0.n10_adj_4230\ : std_logic;
signal \c0.data_in_frame_13_4\ : std_logic;
signal \c0.data_in_frame_15_5\ : std_logic;
signal \c0.data_in_frame_26_3\ : std_logic;
signal \c0.n20266\ : std_logic;
signal \c0.n22402_cascade_\ : std_logic;
signal \c0.n33\ : std_logic;
signal \c0.n21054\ : std_logic;
signal \c0.n6_adj_4292_cascade_\ : std_logic;
signal \c0.data_in_frame_28_5\ : std_logic;
signal \c0.n23073\ : std_logic;
signal \c0.data_in_frame_21_4\ : std_logic;
signal \c0.n21905\ : std_logic;
signal \c0.n21905_cascade_\ : std_logic;
signal \c0.n21069\ : std_logic;
signal \c0.n22113\ : std_logic;
signal \c0.data_in_frame_20_3\ : std_logic;
signal \c0.n20203\ : std_logic;
signal \c0.n21870\ : std_logic;
signal \c0.n18_adj_4249_cascade_\ : std_logic;
signal \c0.n24_adj_4248\ : std_logic;
signal \c0.n26_adj_4250\ : std_logic;
signal \c0.data_in_frame_15_4\ : std_logic;
signal \c0.n23072\ : std_logic;
signal \c0.n13457\ : std_logic;
signal \c0.n23072_cascade_\ : std_logic;
signal \c0.n21067\ : std_logic;
signal \c0.n14_adj_4251\ : std_logic;
signal \c0.data_in_frame_19_5\ : std_logic;
signal \c0.data_in_frame_26_1\ : std_logic;
signal \c0.n21039\ : std_logic;
signal \c0.n24_adj_4282_cascade_\ : std_logic;
signal \c0.n22711\ : std_logic;
signal \c0.n22711_cascade_\ : std_logic;
signal \c0.n21200\ : std_logic;
signal \c0.n12596\ : std_logic;
signal \c0.n6707\ : std_logic;
signal \c0.n15_adj_4284_cascade_\ : std_logic;
signal \c0.n14_adj_4283\ : std_logic;
signal \c0.n22437\ : std_logic;
signal \c0.data_in_frame_25_0\ : std_logic;
signal \c0.data_in_frame_25_6\ : std_logic;
signal \c0.n22437_cascade_\ : std_logic;
signal \c0.n50_adj_4487\ : std_logic;
signal \c0.n22323\ : std_logic;
signal \c0.n10_adj_4483\ : std_logic;
signal \c0.n20537_cascade_\ : std_logic;
signal \c0.n14_adj_4484\ : std_logic;
signal \c0.n21890\ : std_logic;
signal \c0.n21087\ : std_logic;
signal \c0.n13320_cascade_\ : std_logic;
signal \c0.n22468\ : std_logic;
signal \c0.n10_cascade_\ : std_logic;
signal \c0.n20537\ : std_logic;
signal \c0.n22314\ : std_logic;
signal \c0.data_in_frame_24_3\ : std_logic;
signal \c0.n22142\ : std_logic;
signal \c0.data_in_frame_24_4\ : std_logic;
signal \c0.n22028\ : std_logic;
signal \c0.n22337_cascade_\ : std_logic;
signal \c0.n22020\ : std_logic;
signal \c0.n21095\ : std_logic;
signal \c0.n6_adj_4418\ : std_logic;
signal \c0.data_in_frame_26_4\ : std_logic;
signal \c0.n22337\ : std_logic;
signal \c0.n10_adj_4285_cascade_\ : std_logic;
signal \c0.n22995\ : std_logic;
signal \c0.data_in_frame_26_6\ : std_logic;
signal \c0.n22054\ : std_logic;
signal \c0.data_in_frame_24_6\ : std_logic;
signal \c0.n22434\ : std_logic;
signal \c0.data_in_frame_20_0\ : std_logic;
signal data_in_frame_22_2 : std_logic;
signal \c0.n12594\ : std_logic;
signal \c0.n20596\ : std_logic;
signal \c0.data_in_frame_11_7\ : std_logic;
signal n21760 : std_logic;
signal \c0.data_in_frame_26_2\ : std_logic;
signal \c0.n13993\ : std_logic;
signal n91 : std_logic;
signal n12973 : std_logic;
signal n14917 : std_logic;
signal n14436 : std_logic;
signal \r_Bit_Index_1\ : std_logic;
signal data_in_frame_22_4 : std_logic;
signal \c0.n22191\ : std_logic;
signal \c0.n25\ : std_logic;
signal \r_Bit_Index_0\ : std_logic;
signal \r_Rx_Data\ : std_logic;
signal n12970 : std_logic;
signal \c0.data_in_frame_12_0\ : std_logic;
signal \c0.data_in_frame_24_7\ : std_logic;
signal \c0.data_in_frame_12_1\ : std_logic;
signal \c0.data_in_frame_12_2\ : std_logic;
signal \c0.data_in_frame_13_2\ : std_logic;
signal \c0.data_in_frame_13_1\ : std_logic;
signal \c0.data_in_frame_11_0\ : std_logic;
signal \c0.n22274\ : std_logic;
signal \c0.data_in_frame_10_6\ : std_logic;
signal \c0.n13999_cascade_\ : std_logic;
signal \c0.n21940\ : std_logic;
signal \c0.n13233\ : std_logic;
signal \c0.data_in_frame_9_2\ : std_logic;
signal \c0.n21845\ : std_logic;
signal \c0.n22781\ : std_logic;
signal \c0.data_in_frame_11_1\ : std_logic;
signal \c0.data_in_frame_23_3\ : std_logic;
signal \c0.n22236\ : std_logic;
signal \c0.n4\ : std_logic;
signal \c0.n5965\ : std_logic;
signal \c0.n8_adj_4275\ : std_logic;
signal \c0.n8_adj_4276\ : std_logic;
signal \c0.data_in_frame_13_0\ : std_logic;
signal \c0.data_in_frame_12_7\ : std_logic;
signal \c0.data_in_frame_23_1\ : std_logic;
signal data_in_frame_22_7 : std_logic;
signal \c0.n21995\ : std_logic;
signal \c0.data_in_frame_21_7\ : std_logic;
signal \c0.n13210\ : std_logic;
signal \c0.n22091\ : std_logic;
signal \c0.n21934\ : std_logic;
signal \c0.data_in_frame_4_5\ : std_logic;
signal \c0.n13421\ : std_logic;
signal \c0.data_in_frame_11_4\ : std_logic;
signal \c0.n13421_cascade_\ : std_logic;
signal \c0.n22069\ : std_logic;
signal \c0.n10_adj_4252\ : std_logic;
signal \c0.data_in_frame_7_2\ : std_logic;
signal \c0.n22343\ : std_logic;
signal \c0.n10_adj_4267\ : std_logic;
signal \c0.data_in_frame_12_5\ : std_logic;
signal \c0.n16_adj_4268\ : std_logic;
signal \c0.n21740\ : std_logic;
signal \c0.data_in_frame_7_0\ : std_logic;
signal \c0.data_in_frame_16_1\ : std_logic;
signal \c0.data_in_frame_12_3\ : std_logic;
signal \c0.n21975\ : std_logic;
signal \c0.data_in_frame_17_2\ : std_logic;
signal \c0.data_in_frame_15_1\ : std_logic;
signal \c0.data_in_frame_12_4\ : std_logic;
signal \c0.data_in_frame_13_3\ : std_logic;
signal \c0.data_in_frame_13_5\ : std_logic;
signal \c0.n14081\ : std_logic;
signal \c0.data_in_frame_16_0\ : std_logic;
signal \c0.data_in_frame_20_4\ : std_logic;
signal data_in_frame_22_6 : std_logic;
signal \c0.n20246\ : std_logic;
signal \c0.data_in_frame_13_6\ : std_logic;
signal \c0.data_in_frame_26_5\ : std_logic;
signal \c0.data_in_frame_21_6\ : std_logic;
signal \c0.n21749\ : std_logic;
signal \c0.n9_adj_4237\ : std_logic;
signal \c0.data_in_frame_13_7\ : std_logic;
signal \c0.n22388\ : std_logic;
signal \c0.data_in_frame_17_6\ : std_logic;
signal \c0.n20_adj_4247\ : std_logic;
signal \c0.data_in_frame_20_2\ : std_logic;
signal \c0.n13544\ : std_logic;
signal data_in_frame_22_3 : std_logic;
signal \c0.n23426\ : std_logic;
signal \c0.n22007\ : std_logic;
signal \c0.data_in_frame_19_6\ : std_logic;
signal \c0.data_in_frame_18_5\ : std_logic;
signal \c0.n22385\ : std_logic;
signal \c0.n21126\ : std_logic;
signal \c0.data_in_frame_19_1\ : std_logic;
signal \c0.n22084\ : std_logic;
signal \c0.n22364\ : std_logic;
signal \c0.data_in_frame_19_7\ : std_logic;
signal \c0.n15\ : std_logic;
signal \c0.data_in_frame_20_5\ : std_logic;
signal \c0.data_in_frame_23_0\ : std_logic;
signal \c0.n26_adj_4281\ : std_logic;
signal rx_data_4 : std_logic;
signal \c0.data_in_frame_18_3\ : std_logic;
signal \c0.n22095\ : std_logic;
signal \c0.n21124\ : std_logic;
signal \c0.n22095_cascade_\ : std_logic;
signal \c0.n14143\ : std_logic;
signal \c0.n29\ : std_logic;
signal data_in_frame_22_0 : std_logic;
signal \c0.n22267\ : std_logic;
signal \c0.n22105\ : std_logic;
signal \c0.n22849\ : std_logic;
signal \c0.n20406\ : std_logic;
signal \c0.n5813\ : std_logic;
signal \c0.n21864\ : std_logic;
signal \c0.n13768\ : std_logic;
signal \c0.n22458\ : std_logic;
signal \c0.n21114\ : std_logic;
signal \c0.n18_adj_4246\ : std_logic;
signal \c0.n21_cascade_\ : std_logic;
signal \c0.n22399\ : std_logic;
signal \c0.n24\ : std_logic;
signal \c0.n20\ : std_logic;
signal \c0.data_in_frame_17_1\ : std_logic;
signal \c0.n16\ : std_logic;
signal \c0.n21979\ : std_logic;
signal \c0.n23287\ : std_logic;
signal \c0.n23287_cascade_\ : std_logic;
signal \c0.data_in_frame_19_3\ : std_logic;
signal \c0.n21921\ : std_logic;
signal rx_data_1 : std_logic;
signal \c0.data_in_frame_24_0\ : std_logic;
signal \c0.data_in_frame_24_5\ : std_logic;
signal \c0.n13320\ : std_logic;
signal data_in_frame_22_5 : std_logic;
signal \c0.n22255\ : std_logic;
signal \c0.data_in_frame_23_7\ : std_logic;
signal \c0.n22396\ : std_logic;
signal \c0.n20288\ : std_logic;
signal \c0.n23\ : std_logic;
signal \c0.data_in_frame_24_2\ : std_logic;
signal \c0.n13443\ : std_logic;
signal \c0.n22358\ : std_logic;
signal \c0.n22099\ : std_logic;
signal \c0.data_in_frame_24_1\ : std_logic;
signal \c0.n22057\ : std_logic;
signal \c0.n22373\ : std_logic;
signal \c0.n8_adj_4288_cascade_\ : std_logic;
signal \c0.n24_adj_4289\ : std_logic;
signal \c0.n22215\ : std_logic;
signal \c0.n22402\ : std_logic;
signal \c0.data_in_frame_28_4\ : std_logic;
signal \c0.n22455\ : std_logic;
signal \c0.n22997\ : std_logic;
signal rx_data_3 : std_logic;
signal \c0.data_in_frame_28_3\ : std_logic;
signal \c0.data_in_frame_28_7\ : std_logic;
signal \c0.n9_adj_4217\ : std_logic;
signal \c0.data_in_frame_28_6\ : std_logic;
signal \c0.data_in_frame_27_7\ : std_logic;
signal \c0.data_in_frame_27_6\ : std_logic;
signal \c0.data_in_frame_27_0\ : std_logic;
signal \c0.n6268\ : std_logic;
signal \c0.n9_adj_4278\ : std_logic;
signal \c0.data_in_frame_16_7\ : std_logic;
signal \c0.data_in_frame_19_0\ : std_logic;
signal rx_data_6 : std_logic;
signal \c0.data_in_frame_18_6\ : std_logic;
signal \c0.data_in_frame_18_7\ : std_logic;
signal \c0.data_in_frame_21_5\ : std_logic;
signal \c0.n22123\ : std_logic;
signal \c0.n9_adj_4302\ : std_logic;
signal \c0.data_in_frame_25_7\ : std_logic;
signal rx_data_0 : std_logic;
signal \c0.data_in_frame_26_0\ : std_logic;
signal \c0.n9_adj_4341\ : std_logic;
signal rx_data_7 : std_logic;
signal \c0.data_in_frame_26_7\ : std_logic;
signal \c0.n17596\ : std_logic;
signal rx_data_2 : std_logic;
signal \c0.n21758\ : std_logic;
signal \c0.data_in_frame_23_2\ : std_logic;
signal \c0.n21775\ : std_logic;
signal \c0.n9\ : std_logic;
signal rx_data_5 : std_logic;
signal \c0.data_in_frame_27_5\ : std_logic;
signal \PIN_9_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \PIN_12_wire\ : std_logic;
signal \PIN_13_wire\ : std_logic;
signal \PIN_1_wire\ : std_logic;
signal \PIN_22_wire\ : std_logic;
signal \PIN_23_wire\ : std_logic;
signal \PIN_24_wire\ : std_logic;
signal \PIN_2_wire\ : std_logic;
signal \PIN_3_wire\ : std_logic;
signal \PIN_7_wire\ : std_logic;
signal \PIN_8_wire\ : std_logic;
signal \PIN_9_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \pll32MHz_inst.pll20MHz_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK_wire\ <= CLK;
    LED <= \LED_wire\;
    \PIN_12_wire\ <= PIN_12;
    \PIN_13_wire\ <= PIN_13;
    PIN_1 <= \PIN_1_wire\;
    PIN_22 <= \PIN_22_wire\;
    PIN_23 <= \PIN_23_wire\;
    PIN_24 <= \PIN_24_wire\;
    PIN_2 <= \PIN_2_wire\;
    PIN_3 <= \PIN_3_wire\;
    \PIN_7_wire\ <= PIN_7;
    \PIN_8_wire\ <= PIN_8;
    PIN_9 <= \PIN_9_wire\;
    USBPU <= \USBPU_wire\;
    \pll32MHz_inst.pll20MHz_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';

    \pll32MHz_inst.pll20MHz_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "SHIFTREG_0deg",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "PHASE_AND_DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            BYPASS => \GNDG0\,
            DYNAMICDELAY => \pll32MHz_inst.pll20MHz_inst_DYNAMICDELAY_wire\,
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            PLLOUTGLOBAL => \PIN_9_c\,
            REFERENCECLK => \N__23719\,
            RESETB => \N__47218\,
            SCLK => '0',
            SDI => '0',
            SDO => OPEN
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__70064\,
            DIN => \N__70063\,
            DOUT => \N__70062\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__70064\,
            PADOUT => \N__70063\,
            PADIN => \N__70062\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__70055\,
            DIN => \N__70054\,
            DOUT => \N__70053\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__70055\,
            PADOUT => \N__70054\,
            PADIN => \N__70053\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__23683\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_12_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__70046\,
            DIN => \N__70045\,
            DOUT => \N__70044\,
            PACKAGEPIN => \PIN_12_wire\
        );

    \PIN_12_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__70046\,
            PADOUT => \N__70045\,
            PADIN => \N__70044\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_12_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_13_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__70037\,
            DIN => \N__70036\,
            DOUT => \N__70035\,
            PACKAGEPIN => \PIN_13_wire\
        );

    \PIN_13_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__70037\,
            PADOUT => \N__70036\,
            PADIN => \N__70035\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_13_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__70028\,
            DIN => \N__70027\,
            DOUT => \N__70026\,
            PACKAGEPIN => \PIN_1_wire\
        );

    \PIN_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__70028\,
            PADOUT => \N__70027\,
            PADIN => \N__70026\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_22_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__70019\,
            DIN => \N__70018\,
            DOUT => \N__70017\,
            PACKAGEPIN => \PIN_22_wire\
        );

    \PIN_22_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__70019\,
            PADOUT => \N__70018\,
            PADIN => \N__70017\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_23_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__70010\,
            DIN => \N__70009\,
            DOUT => \N__70008\,
            PACKAGEPIN => \PIN_23_wire\
        );

    \PIN_23_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__70010\,
            PADOUT => \N__70009\,
            PADIN => \N__70008\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_24_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__70001\,
            DIN => \N__70000\,
            DOUT => \N__69999\,
            PACKAGEPIN => \PIN_24_wire\
        );

    \PIN_24_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__70001\,
            PADOUT => \N__70000\,
            PADIN => \N__69999\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69992\,
            DIN => \N__69991\,
            DOUT => \N__69990\,
            PACKAGEPIN => \PIN_2_wire\
        );

    \PIN_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69992\,
            PADOUT => \N__69991\,
            PADIN => \N__69990\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69983\,
            DIN => \N__69982\,
            DOUT => \N__69981\,
            PACKAGEPIN => \PIN_3_wire\
        );

    \PIN_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69983\,
            PADOUT => \N__69982\,
            PADIN => \N__69981\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69974\,
            DIN => \N__69973\,
            DOUT => \N__69972\,
            PACKAGEPIN => \PIN_7_wire\
        );

    \PIN_7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69974\,
            PADOUT => \N__69973\,
            PADIN => \N__69972\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_7_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_8_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69965\,
            DIN => \N__69964\,
            DOUT => \N__69963\,
            PACKAGEPIN => \PIN_8_wire\
        );

    \PIN_8_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69965\,
            PADOUT => \N__69964\,
            PADIN => \N__69963\,
            CLOCKENABLE => 'H',
            DIN0 => \PIN_8_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \PIN_9_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69956\,
            DIN => \N__69955\,
            DOUT => \N__69954\,
            PACKAGEPIN => \PIN_9_wire\
        );

    \PIN_9_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69956\,
            PADOUT => \N__69955\,
            PADIN => \N__69954\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__23689\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__69947\,
            DIN => \N__69946\,
            DOUT => \N__69945\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69947\,
            PADOUT => \N__69946\,
            PADIN => \N__69945\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall1_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__69938\,
            DIN => \N__69937\,
            DOUT => \N__69936\,
            PACKAGEPIN => PIN_4
        );

    \hall1_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69938\,
            PADOUT => \N__69937\,
            PADIN => \N__69936\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall2_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__69929\,
            DIN => \N__69928\,
            DOUT => \N__69927\,
            PACKAGEPIN => PIN_5
        );

    \hall2_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69929\,
            PADOUT => \N__69928\,
            PADIN => \N__69927\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall3_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__69920\,
            DIN => \N__69919\,
            DOUT => \N__69918\,
            PACKAGEPIN => PIN_6
        );

    \hall3_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69920\,
            PADOUT => \N__69919\,
            PADIN => \N__69918\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rx_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__69911\,
            DIN => \N__69910\,
            DOUT => \N__69909\,
            PACKAGEPIN => PIN_11
        );

    \rx_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69911\,
            PADOUT => \N__69910\,
            PADIN => \N__69909\,
            CLOCKENABLE => 'H',
            DIN0 => rx_i,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \tx_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__69902\,
            DIN => \N__69901\,
            DOUT => \N__69900\,
            PACKAGEPIN => PIN_10
        );

    \tx_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__69902\,
            PADOUT => \N__69901\,
            PADIN => \N__69900\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__26524\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__23695\
        );

    \I__17391\ : InMux
    port map (
            O => \N__69883\,
            I => \N__69873\
        );

    \I__17390\ : CascadeMux
    port map (
            O => \N__69882\,
            I => \N__69868\
        );

    \I__17389\ : CascadeMux
    port map (
            O => \N__69881\,
            I => \N__69861\
        );

    \I__17388\ : InMux
    port map (
            O => \N__69880\,
            I => \N__69857\
        );

    \I__17387\ : InMux
    port map (
            O => \N__69879\,
            I => \N__69854\
        );

    \I__17386\ : CascadeMux
    port map (
            O => \N__69878\,
            I => \N__69851\
        );

    \I__17385\ : CascadeMux
    port map (
            O => \N__69877\,
            I => \N__69848\
        );

    \I__17384\ : CascadeMux
    port map (
            O => \N__69876\,
            I => \N__69841\
        );

    \I__17383\ : LocalMux
    port map (
            O => \N__69873\,
            I => \N__69836\
        );

    \I__17382\ : InMux
    port map (
            O => \N__69872\,
            I => \N__69833\
        );

    \I__17381\ : InMux
    port map (
            O => \N__69871\,
            I => \N__69830\
        );

    \I__17380\ : InMux
    port map (
            O => \N__69868\,
            I => \N__69827\
        );

    \I__17379\ : InMux
    port map (
            O => \N__69867\,
            I => \N__69824\
        );

    \I__17378\ : CascadeMux
    port map (
            O => \N__69866\,
            I => \N__69821\
        );

    \I__17377\ : InMux
    port map (
            O => \N__69865\,
            I => \N__69818\
        );

    \I__17376\ : InMux
    port map (
            O => \N__69864\,
            I => \N__69815\
        );

    \I__17375\ : InMux
    port map (
            O => \N__69861\,
            I => \N__69810\
        );

    \I__17374\ : InMux
    port map (
            O => \N__69860\,
            I => \N__69810\
        );

    \I__17373\ : LocalMux
    port map (
            O => \N__69857\,
            I => \N__69807\
        );

    \I__17372\ : LocalMux
    port map (
            O => \N__69854\,
            I => \N__69803\
        );

    \I__17371\ : InMux
    port map (
            O => \N__69851\,
            I => \N__69798\
        );

    \I__17370\ : InMux
    port map (
            O => \N__69848\,
            I => \N__69795\
        );

    \I__17369\ : InMux
    port map (
            O => \N__69847\,
            I => \N__69791\
        );

    \I__17368\ : InMux
    port map (
            O => \N__69846\,
            I => \N__69784\
        );

    \I__17367\ : InMux
    port map (
            O => \N__69845\,
            I => \N__69784\
        );

    \I__17366\ : InMux
    port map (
            O => \N__69844\,
            I => \N__69784\
        );

    \I__17365\ : InMux
    port map (
            O => \N__69841\,
            I => \N__69781\
        );

    \I__17364\ : InMux
    port map (
            O => \N__69840\,
            I => \N__69778\
        );

    \I__17363\ : InMux
    port map (
            O => \N__69839\,
            I => \N__69774\
        );

    \I__17362\ : Span4Mux_v
    port map (
            O => \N__69836\,
            I => \N__69771\
        );

    \I__17361\ : LocalMux
    port map (
            O => \N__69833\,
            I => \N__69766\
        );

    \I__17360\ : LocalMux
    port map (
            O => \N__69830\,
            I => \N__69766\
        );

    \I__17359\ : LocalMux
    port map (
            O => \N__69827\,
            I => \N__69761\
        );

    \I__17358\ : LocalMux
    port map (
            O => \N__69824\,
            I => \N__69761\
        );

    \I__17357\ : InMux
    port map (
            O => \N__69821\,
            I => \N__69758\
        );

    \I__17356\ : LocalMux
    port map (
            O => \N__69818\,
            I => \N__69751\
        );

    \I__17355\ : LocalMux
    port map (
            O => \N__69815\,
            I => \N__69751\
        );

    \I__17354\ : LocalMux
    port map (
            O => \N__69810\,
            I => \N__69751\
        );

    \I__17353\ : Span4Mux_h
    port map (
            O => \N__69807\,
            I => \N__69747\
        );

    \I__17352\ : InMux
    port map (
            O => \N__69806\,
            I => \N__69744\
        );

    \I__17351\ : Span4Mux_v
    port map (
            O => \N__69803\,
            I => \N__69741\
        );

    \I__17350\ : InMux
    port map (
            O => \N__69802\,
            I => \N__69736\
        );

    \I__17349\ : InMux
    port map (
            O => \N__69801\,
            I => \N__69736\
        );

    \I__17348\ : LocalMux
    port map (
            O => \N__69798\,
            I => \N__69731\
        );

    \I__17347\ : LocalMux
    port map (
            O => \N__69795\,
            I => \N__69731\
        );

    \I__17346\ : CascadeMux
    port map (
            O => \N__69794\,
            I => \N__69727\
        );

    \I__17345\ : LocalMux
    port map (
            O => \N__69791\,
            I => \N__69720\
        );

    \I__17344\ : LocalMux
    port map (
            O => \N__69784\,
            I => \N__69720\
        );

    \I__17343\ : LocalMux
    port map (
            O => \N__69781\,
            I => \N__69720\
        );

    \I__17342\ : LocalMux
    port map (
            O => \N__69778\,
            I => \N__69717\
        );

    \I__17341\ : CascadeMux
    port map (
            O => \N__69777\,
            I => \N__69713\
        );

    \I__17340\ : LocalMux
    port map (
            O => \N__69774\,
            I => \N__69710\
        );

    \I__17339\ : Span4Mux_h
    port map (
            O => \N__69771\,
            I => \N__69703\
        );

    \I__17338\ : Span4Mux_v
    port map (
            O => \N__69766\,
            I => \N__69703\
        );

    \I__17337\ : Span4Mux_v
    port map (
            O => \N__69761\,
            I => \N__69703\
        );

    \I__17336\ : LocalMux
    port map (
            O => \N__69758\,
            I => \N__69698\
        );

    \I__17335\ : Span4Mux_v
    port map (
            O => \N__69751\,
            I => \N__69698\
        );

    \I__17334\ : InMux
    port map (
            O => \N__69750\,
            I => \N__69692\
        );

    \I__17333\ : Span4Mux_h
    port map (
            O => \N__69747\,
            I => \N__69687\
        );

    \I__17332\ : LocalMux
    port map (
            O => \N__69744\,
            I => \N__69687\
        );

    \I__17331\ : Span4Mux_h
    port map (
            O => \N__69741\,
            I => \N__69680\
        );

    \I__17330\ : LocalMux
    port map (
            O => \N__69736\,
            I => \N__69680\
        );

    \I__17329\ : Span4Mux_h
    port map (
            O => \N__69731\,
            I => \N__69680\
        );

    \I__17328\ : InMux
    port map (
            O => \N__69730\,
            I => \N__69677\
        );

    \I__17327\ : InMux
    port map (
            O => \N__69727\,
            I => \N__69674\
        );

    \I__17326\ : Span4Mux_v
    port map (
            O => \N__69720\,
            I => \N__69669\
        );

    \I__17325\ : Span4Mux_v
    port map (
            O => \N__69717\,
            I => \N__69669\
        );

    \I__17324\ : InMux
    port map (
            O => \N__69716\,
            I => \N__69666\
        );

    \I__17323\ : InMux
    port map (
            O => \N__69713\,
            I => \N__69663\
        );

    \I__17322\ : Span4Mux_h
    port map (
            O => \N__69710\,
            I => \N__69656\
        );

    \I__17321\ : Span4Mux_h
    port map (
            O => \N__69703\,
            I => \N__69656\
        );

    \I__17320\ : Span4Mux_v
    port map (
            O => \N__69698\,
            I => \N__69656\
        );

    \I__17319\ : InMux
    port map (
            O => \N__69697\,
            I => \N__69649\
        );

    \I__17318\ : InMux
    port map (
            O => \N__69696\,
            I => \N__69649\
        );

    \I__17317\ : InMux
    port map (
            O => \N__69695\,
            I => \N__69649\
        );

    \I__17316\ : LocalMux
    port map (
            O => \N__69692\,
            I => \N__69646\
        );

    \I__17315\ : Span4Mux_v
    port map (
            O => \N__69687\,
            I => \N__69641\
        );

    \I__17314\ : Span4Mux_v
    port map (
            O => \N__69680\,
            I => \N__69641\
        );

    \I__17313\ : LocalMux
    port map (
            O => \N__69677\,
            I => \N__69638\
        );

    \I__17312\ : LocalMux
    port map (
            O => \N__69674\,
            I => \N__69633\
        );

    \I__17311\ : Span4Mux_v
    port map (
            O => \N__69669\,
            I => \N__69633\
        );

    \I__17310\ : LocalMux
    port map (
            O => \N__69666\,
            I => \N__69630\
        );

    \I__17309\ : LocalMux
    port map (
            O => \N__69663\,
            I => \N__69625\
        );

    \I__17308\ : Span4Mux_v
    port map (
            O => \N__69656\,
            I => \N__69625\
        );

    \I__17307\ : LocalMux
    port map (
            O => \N__69649\,
            I => \N__69616\
        );

    \I__17306\ : Sp12to4
    port map (
            O => \N__69646\,
            I => \N__69616\
        );

    \I__17305\ : Sp12to4
    port map (
            O => \N__69641\,
            I => \N__69616\
        );

    \I__17304\ : Span12Mux_v
    port map (
            O => \N__69638\,
            I => \N__69616\
        );

    \I__17303\ : Span4Mux_v
    port map (
            O => \N__69633\,
            I => \N__69613\
        );

    \I__17302\ : Span4Mux_v
    port map (
            O => \N__69630\,
            I => \N__69608\
        );

    \I__17301\ : Span4Mux_v
    port map (
            O => \N__69625\,
            I => \N__69608\
        );

    \I__17300\ : Span12Mux_v
    port map (
            O => \N__69616\,
            I => \N__69605\
        );

    \I__17299\ : Span4Mux_v
    port map (
            O => \N__69613\,
            I => \N__69602\
        );

    \I__17298\ : Odrv4
    port map (
            O => \N__69608\,
            I => \c0.n9_adj_4302\
        );

    \I__17297\ : Odrv12
    port map (
            O => \N__69605\,
            I => \c0.n9_adj_4302\
        );

    \I__17296\ : Odrv4
    port map (
            O => \N__69602\,
            I => \c0.n9_adj_4302\
        );

    \I__17295\ : InMux
    port map (
            O => \N__69595\,
            I => \N__69591\
        );

    \I__17294\ : CascadeMux
    port map (
            O => \N__69594\,
            I => \N__69588\
        );

    \I__17293\ : LocalMux
    port map (
            O => \N__69591\,
            I => \N__69585\
        );

    \I__17292\ : InMux
    port map (
            O => \N__69588\,
            I => \N__69581\
        );

    \I__17291\ : Span4Mux_v
    port map (
            O => \N__69585\,
            I => \N__69578\
        );

    \I__17290\ : InMux
    port map (
            O => \N__69584\,
            I => \N__69575\
        );

    \I__17289\ : LocalMux
    port map (
            O => \N__69581\,
            I => \c0.data_in_frame_25_7\
        );

    \I__17288\ : Odrv4
    port map (
            O => \N__69578\,
            I => \c0.data_in_frame_25_7\
        );

    \I__17287\ : LocalMux
    port map (
            O => \N__69575\,
            I => \c0.data_in_frame_25_7\
        );

    \I__17286\ : InMux
    port map (
            O => \N__69568\,
            I => \N__69552\
        );

    \I__17285\ : InMux
    port map (
            O => \N__69567\,
            I => \N__69549\
        );

    \I__17284\ : InMux
    port map (
            O => \N__69566\,
            I => \N__69545\
        );

    \I__17283\ : InMux
    port map (
            O => \N__69565\,
            I => \N__69542\
        );

    \I__17282\ : InMux
    port map (
            O => \N__69564\,
            I => \N__69539\
        );

    \I__17281\ : InMux
    port map (
            O => \N__69563\,
            I => \N__69534\
        );

    \I__17280\ : InMux
    port map (
            O => \N__69562\,
            I => \N__69529\
        );

    \I__17279\ : InMux
    port map (
            O => \N__69561\,
            I => \N__69529\
        );

    \I__17278\ : InMux
    port map (
            O => \N__69560\,
            I => \N__69526\
        );

    \I__17277\ : InMux
    port map (
            O => \N__69559\,
            I => \N__69521\
        );

    \I__17276\ : InMux
    port map (
            O => \N__69558\,
            I => \N__69521\
        );

    \I__17275\ : InMux
    port map (
            O => \N__69557\,
            I => \N__69518\
        );

    \I__17274\ : InMux
    port map (
            O => \N__69556\,
            I => \N__69513\
        );

    \I__17273\ : InMux
    port map (
            O => \N__69555\,
            I => \N__69513\
        );

    \I__17272\ : LocalMux
    port map (
            O => \N__69552\,
            I => \N__69510\
        );

    \I__17271\ : LocalMux
    port map (
            O => \N__69549\,
            I => \N__69507\
        );

    \I__17270\ : InMux
    port map (
            O => \N__69548\,
            I => \N__69504\
        );

    \I__17269\ : LocalMux
    port map (
            O => \N__69545\,
            I => \N__69497\
        );

    \I__17268\ : LocalMux
    port map (
            O => \N__69542\,
            I => \N__69497\
        );

    \I__17267\ : LocalMux
    port map (
            O => \N__69539\,
            I => \N__69494\
        );

    \I__17266\ : InMux
    port map (
            O => \N__69538\,
            I => \N__69488\
        );

    \I__17265\ : InMux
    port map (
            O => \N__69537\,
            I => \N__69483\
        );

    \I__17264\ : LocalMux
    port map (
            O => \N__69534\,
            I => \N__69477\
        );

    \I__17263\ : LocalMux
    port map (
            O => \N__69529\,
            I => \N__69474\
        );

    \I__17262\ : LocalMux
    port map (
            O => \N__69526\,
            I => \N__69471\
        );

    \I__17261\ : LocalMux
    port map (
            O => \N__69521\,
            I => \N__69468\
        );

    \I__17260\ : LocalMux
    port map (
            O => \N__69518\,
            I => \N__69465\
        );

    \I__17259\ : LocalMux
    port map (
            O => \N__69513\,
            I => \N__69456\
        );

    \I__17258\ : Span4Mux_h
    port map (
            O => \N__69510\,
            I => \N__69456\
        );

    \I__17257\ : Span4Mux_v
    port map (
            O => \N__69507\,
            I => \N__69456\
        );

    \I__17256\ : LocalMux
    port map (
            O => \N__69504\,
            I => \N__69456\
        );

    \I__17255\ : InMux
    port map (
            O => \N__69503\,
            I => \N__69453\
        );

    \I__17254\ : InMux
    port map (
            O => \N__69502\,
            I => \N__69447\
        );

    \I__17253\ : Span4Mux_v
    port map (
            O => \N__69497\,
            I => \N__69442\
        );

    \I__17252\ : Span4Mux_h
    port map (
            O => \N__69494\,
            I => \N__69442\
        );

    \I__17251\ : InMux
    port map (
            O => \N__69493\,
            I => \N__69439\
        );

    \I__17250\ : InMux
    port map (
            O => \N__69492\,
            I => \N__69436\
        );

    \I__17249\ : InMux
    port map (
            O => \N__69491\,
            I => \N__69433\
        );

    \I__17248\ : LocalMux
    port map (
            O => \N__69488\,
            I => \N__69430\
        );

    \I__17247\ : InMux
    port map (
            O => \N__69487\,
            I => \N__69427\
        );

    \I__17246\ : InMux
    port map (
            O => \N__69486\,
            I => \N__69424\
        );

    \I__17245\ : LocalMux
    port map (
            O => \N__69483\,
            I => \N__69421\
        );

    \I__17244\ : InMux
    port map (
            O => \N__69482\,
            I => \N__69418\
        );

    \I__17243\ : InMux
    port map (
            O => \N__69481\,
            I => \N__69413\
        );

    \I__17242\ : InMux
    port map (
            O => \N__69480\,
            I => \N__69413\
        );

    \I__17241\ : Span4Mux_h
    port map (
            O => \N__69477\,
            I => \N__69410\
        );

    \I__17240\ : Span4Mux_h
    port map (
            O => \N__69474\,
            I => \N__69405\
        );

    \I__17239\ : Span4Mux_v
    port map (
            O => \N__69471\,
            I => \N__69405\
        );

    \I__17238\ : Span4Mux_v
    port map (
            O => \N__69468\,
            I => \N__69400\
        );

    \I__17237\ : Span4Mux_h
    port map (
            O => \N__69465\,
            I => \N__69400\
        );

    \I__17236\ : Span4Mux_h
    port map (
            O => \N__69456\,
            I => \N__69397\
        );

    \I__17235\ : LocalMux
    port map (
            O => \N__69453\,
            I => \N__69394\
        );

    \I__17234\ : InMux
    port map (
            O => \N__69452\,
            I => \N__69391\
        );

    \I__17233\ : InMux
    port map (
            O => \N__69451\,
            I => \N__69388\
        );

    \I__17232\ : InMux
    port map (
            O => \N__69450\,
            I => \N__69385\
        );

    \I__17231\ : LocalMux
    port map (
            O => \N__69447\,
            I => \N__69376\
        );

    \I__17230\ : Span4Mux_h
    port map (
            O => \N__69442\,
            I => \N__69376\
        );

    \I__17229\ : LocalMux
    port map (
            O => \N__69439\,
            I => \N__69376\
        );

    \I__17228\ : LocalMux
    port map (
            O => \N__69436\,
            I => \N__69376\
        );

    \I__17227\ : LocalMux
    port map (
            O => \N__69433\,
            I => \N__69371\
        );

    \I__17226\ : Span4Mux_h
    port map (
            O => \N__69430\,
            I => \N__69368\
        );

    \I__17225\ : LocalMux
    port map (
            O => \N__69427\,
            I => \N__69365\
        );

    \I__17224\ : LocalMux
    port map (
            O => \N__69424\,
            I => \N__69360\
        );

    \I__17223\ : Span4Mux_h
    port map (
            O => \N__69421\,
            I => \N__69360\
        );

    \I__17222\ : LocalMux
    port map (
            O => \N__69418\,
            I => \N__69355\
        );

    \I__17221\ : LocalMux
    port map (
            O => \N__69413\,
            I => \N__69355\
        );

    \I__17220\ : Span4Mux_v
    port map (
            O => \N__69410\,
            I => \N__69352\
        );

    \I__17219\ : Span4Mux_h
    port map (
            O => \N__69405\,
            I => \N__69349\
        );

    \I__17218\ : Span4Mux_h
    port map (
            O => \N__69400\,
            I => \N__69344\
        );

    \I__17217\ : Span4Mux_v
    port map (
            O => \N__69397\,
            I => \N__69344\
        );

    \I__17216\ : Span4Mux_v
    port map (
            O => \N__69394\,
            I => \N__69341\
        );

    \I__17215\ : LocalMux
    port map (
            O => \N__69391\,
            I => \N__69338\
        );

    \I__17214\ : LocalMux
    port map (
            O => \N__69388\,
            I => \N__69335\
        );

    \I__17213\ : LocalMux
    port map (
            O => \N__69385\,
            I => \N__69330\
        );

    \I__17212\ : Sp12to4
    port map (
            O => \N__69376\,
            I => \N__69330\
        );

    \I__17211\ : InMux
    port map (
            O => \N__69375\,
            I => \N__69327\
        );

    \I__17210\ : InMux
    port map (
            O => \N__69374\,
            I => \N__69324\
        );

    \I__17209\ : Span4Mux_h
    port map (
            O => \N__69371\,
            I => \N__69319\
        );

    \I__17208\ : Span4Mux_h
    port map (
            O => \N__69368\,
            I => \N__69319\
        );

    \I__17207\ : Span4Mux_h
    port map (
            O => \N__69365\,
            I => \N__69314\
        );

    \I__17206\ : Span4Mux_h
    port map (
            O => \N__69360\,
            I => \N__69314\
        );

    \I__17205\ : Span12Mux_h
    port map (
            O => \N__69355\,
            I => \N__69309\
        );

    \I__17204\ : Sp12to4
    port map (
            O => \N__69352\,
            I => \N__69309\
        );

    \I__17203\ : Span4Mux_h
    port map (
            O => \N__69349\,
            I => \N__69304\
        );

    \I__17202\ : Span4Mux_v
    port map (
            O => \N__69344\,
            I => \N__69304\
        );

    \I__17201\ : Sp12to4
    port map (
            O => \N__69341\,
            I => \N__69295\
        );

    \I__17200\ : Span12Mux_v
    port map (
            O => \N__69338\,
            I => \N__69295\
        );

    \I__17199\ : Span12Mux_s8_h
    port map (
            O => \N__69335\,
            I => \N__69295\
        );

    \I__17198\ : Span12Mux_v
    port map (
            O => \N__69330\,
            I => \N__69295\
        );

    \I__17197\ : LocalMux
    port map (
            O => \N__69327\,
            I => rx_data_0
        );

    \I__17196\ : LocalMux
    port map (
            O => \N__69324\,
            I => rx_data_0
        );

    \I__17195\ : Odrv4
    port map (
            O => \N__69319\,
            I => rx_data_0
        );

    \I__17194\ : Odrv4
    port map (
            O => \N__69314\,
            I => rx_data_0
        );

    \I__17193\ : Odrv12
    port map (
            O => \N__69309\,
            I => rx_data_0
        );

    \I__17192\ : Odrv4
    port map (
            O => \N__69304\,
            I => rx_data_0
        );

    \I__17191\ : Odrv12
    port map (
            O => \N__69295\,
            I => rx_data_0
        );

    \I__17190\ : InMux
    port map (
            O => \N__69280\,
            I => \N__69276\
        );

    \I__17189\ : CascadeMux
    port map (
            O => \N__69279\,
            I => \N__69273\
        );

    \I__17188\ : LocalMux
    port map (
            O => \N__69276\,
            I => \N__69270\
        );

    \I__17187\ : InMux
    port map (
            O => \N__69273\,
            I => \N__69266\
        );

    \I__17186\ : Span4Mux_h
    port map (
            O => \N__69270\,
            I => \N__69263\
        );

    \I__17185\ : InMux
    port map (
            O => \N__69269\,
            I => \N__69260\
        );

    \I__17184\ : LocalMux
    port map (
            O => \N__69266\,
            I => \c0.data_in_frame_26_0\
        );

    \I__17183\ : Odrv4
    port map (
            O => \N__69263\,
            I => \c0.data_in_frame_26_0\
        );

    \I__17182\ : LocalMux
    port map (
            O => \N__69260\,
            I => \c0.data_in_frame_26_0\
        );

    \I__17181\ : CascadeMux
    port map (
            O => \N__69253\,
            I => \N__69250\
        );

    \I__17180\ : InMux
    port map (
            O => \N__69250\,
            I => \N__69246\
        );

    \I__17179\ : InMux
    port map (
            O => \N__69249\,
            I => \N__69241\
        );

    \I__17178\ : LocalMux
    port map (
            O => \N__69246\,
            I => \N__69238\
        );

    \I__17177\ : CascadeMux
    port map (
            O => \N__69245\,
            I => \N__69235\
        );

    \I__17176\ : CascadeMux
    port map (
            O => \N__69244\,
            I => \N__69228\
        );

    \I__17175\ : LocalMux
    port map (
            O => \N__69241\,
            I => \N__69223\
        );

    \I__17174\ : Span4Mux_h
    port map (
            O => \N__69238\,
            I => \N__69220\
        );

    \I__17173\ : InMux
    port map (
            O => \N__69235\,
            I => \N__69217\
        );

    \I__17172\ : CascadeMux
    port map (
            O => \N__69234\,
            I => \N__69214\
        );

    \I__17171\ : CascadeMux
    port map (
            O => \N__69233\,
            I => \N__69207\
        );

    \I__17170\ : CascadeMux
    port map (
            O => \N__69232\,
            I => \N__69200\
        );

    \I__17169\ : InMux
    port map (
            O => \N__69231\,
            I => \N__69194\
        );

    \I__17168\ : InMux
    port map (
            O => \N__69228\,
            I => \N__69184\
        );

    \I__17167\ : InMux
    port map (
            O => \N__69227\,
            I => \N__69184\
        );

    \I__17166\ : InMux
    port map (
            O => \N__69226\,
            I => \N__69184\
        );

    \I__17165\ : Span4Mux_h
    port map (
            O => \N__69223\,
            I => \N__69177\
        );

    \I__17164\ : Span4Mux_h
    port map (
            O => \N__69220\,
            I => \N__69177\
        );

    \I__17163\ : LocalMux
    port map (
            O => \N__69217\,
            I => \N__69177\
        );

    \I__17162\ : InMux
    port map (
            O => \N__69214\,
            I => \N__69174\
        );

    \I__17161\ : InMux
    port map (
            O => \N__69213\,
            I => \N__69169\
        );

    \I__17160\ : InMux
    port map (
            O => \N__69212\,
            I => \N__69169\
        );

    \I__17159\ : InMux
    port map (
            O => \N__69211\,
            I => \N__69165\
        );

    \I__17158\ : InMux
    port map (
            O => \N__69210\,
            I => \N__69162\
        );

    \I__17157\ : InMux
    port map (
            O => \N__69207\,
            I => \N__69155\
        );

    \I__17156\ : InMux
    port map (
            O => \N__69206\,
            I => \N__69155\
        );

    \I__17155\ : InMux
    port map (
            O => \N__69205\,
            I => \N__69155\
        );

    \I__17154\ : InMux
    port map (
            O => \N__69204\,
            I => \N__69152\
        );

    \I__17153\ : InMux
    port map (
            O => \N__69203\,
            I => \N__69148\
        );

    \I__17152\ : InMux
    port map (
            O => \N__69200\,
            I => \N__69143\
        );

    \I__17151\ : InMux
    port map (
            O => \N__69199\,
            I => \N__69143\
        );

    \I__17150\ : InMux
    port map (
            O => \N__69198\,
            I => \N__69138\
        );

    \I__17149\ : InMux
    port map (
            O => \N__69197\,
            I => \N__69138\
        );

    \I__17148\ : LocalMux
    port map (
            O => \N__69194\,
            I => \N__69135\
        );

    \I__17147\ : CascadeMux
    port map (
            O => \N__69193\,
            I => \N__69132\
        );

    \I__17146\ : CascadeMux
    port map (
            O => \N__69192\,
            I => \N__69129\
        );

    \I__17145\ : CascadeMux
    port map (
            O => \N__69191\,
            I => \N__69126\
        );

    \I__17144\ : LocalMux
    port map (
            O => \N__69184\,
            I => \N__69119\
        );

    \I__17143\ : Span4Mux_v
    port map (
            O => \N__69177\,
            I => \N__69119\
        );

    \I__17142\ : LocalMux
    port map (
            O => \N__69174\,
            I => \N__69116\
        );

    \I__17141\ : LocalMux
    port map (
            O => \N__69169\,
            I => \N__69113\
        );

    \I__17140\ : InMux
    port map (
            O => \N__69168\,
            I => \N__69110\
        );

    \I__17139\ : LocalMux
    port map (
            O => \N__69165\,
            I => \N__69107\
        );

    \I__17138\ : LocalMux
    port map (
            O => \N__69162\,
            I => \N__69100\
        );

    \I__17137\ : LocalMux
    port map (
            O => \N__69155\,
            I => \N__69100\
        );

    \I__17136\ : LocalMux
    port map (
            O => \N__69152\,
            I => \N__69100\
        );

    \I__17135\ : InMux
    port map (
            O => \N__69151\,
            I => \N__69097\
        );

    \I__17134\ : LocalMux
    port map (
            O => \N__69148\,
            I => \N__69094\
        );

    \I__17133\ : LocalMux
    port map (
            O => \N__69143\,
            I => \N__69089\
        );

    \I__17132\ : LocalMux
    port map (
            O => \N__69138\,
            I => \N__69089\
        );

    \I__17131\ : Span4Mux_v
    port map (
            O => \N__69135\,
            I => \N__69086\
        );

    \I__17130\ : InMux
    port map (
            O => \N__69132\,
            I => \N__69081\
        );

    \I__17129\ : InMux
    port map (
            O => \N__69129\,
            I => \N__69081\
        );

    \I__17128\ : InMux
    port map (
            O => \N__69126\,
            I => \N__69078\
        );

    \I__17127\ : InMux
    port map (
            O => \N__69125\,
            I => \N__69075\
        );

    \I__17126\ : InMux
    port map (
            O => \N__69124\,
            I => \N__69072\
        );

    \I__17125\ : Sp12to4
    port map (
            O => \N__69119\,
            I => \N__69069\
        );

    \I__17124\ : Span4Mux_h
    port map (
            O => \N__69116\,
            I => \N__69066\
        );

    \I__17123\ : Span4Mux_h
    port map (
            O => \N__69113\,
            I => \N__69059\
        );

    \I__17122\ : LocalMux
    port map (
            O => \N__69110\,
            I => \N__69056\
        );

    \I__17121\ : Span4Mux_h
    port map (
            O => \N__69107\,
            I => \N__69053\
        );

    \I__17120\ : Span4Mux_v
    port map (
            O => \N__69100\,
            I => \N__69050\
        );

    \I__17119\ : LocalMux
    port map (
            O => \N__69097\,
            I => \N__69043\
        );

    \I__17118\ : Sp12to4
    port map (
            O => \N__69094\,
            I => \N__69043\
        );

    \I__17117\ : Span12Mux_v
    port map (
            O => \N__69089\,
            I => \N__69043\
        );

    \I__17116\ : Span4Mux_h
    port map (
            O => \N__69086\,
            I => \N__69034\
        );

    \I__17115\ : LocalMux
    port map (
            O => \N__69081\,
            I => \N__69034\
        );

    \I__17114\ : LocalMux
    port map (
            O => \N__69078\,
            I => \N__69034\
        );

    \I__17113\ : LocalMux
    port map (
            O => \N__69075\,
            I => \N__69034\
        );

    \I__17112\ : LocalMux
    port map (
            O => \N__69072\,
            I => \N__69027\
        );

    \I__17111\ : Span12Mux_h
    port map (
            O => \N__69069\,
            I => \N__69027\
        );

    \I__17110\ : Sp12to4
    port map (
            O => \N__69066\,
            I => \N__69027\
        );

    \I__17109\ : InMux
    port map (
            O => \N__69065\,
            I => \N__69018\
        );

    \I__17108\ : InMux
    port map (
            O => \N__69064\,
            I => \N__69018\
        );

    \I__17107\ : InMux
    port map (
            O => \N__69063\,
            I => \N__69018\
        );

    \I__17106\ : InMux
    port map (
            O => \N__69062\,
            I => \N__69018\
        );

    \I__17105\ : Span4Mux_v
    port map (
            O => \N__69059\,
            I => \N__69015\
        );

    \I__17104\ : Span4Mux_v
    port map (
            O => \N__69056\,
            I => \N__69008\
        );

    \I__17103\ : Span4Mux_v
    port map (
            O => \N__69053\,
            I => \N__69008\
        );

    \I__17102\ : Span4Mux_v
    port map (
            O => \N__69050\,
            I => \N__69008\
        );

    \I__17101\ : Span12Mux_v
    port map (
            O => \N__69043\,
            I => \N__69005\
        );

    \I__17100\ : Sp12to4
    port map (
            O => \N__69034\,
            I => \N__69000\
        );

    \I__17099\ : Span12Mux_v
    port map (
            O => \N__69027\,
            I => \N__69000\
        );

    \I__17098\ : LocalMux
    port map (
            O => \N__69018\,
            I => \c0.n9_adj_4341\
        );

    \I__17097\ : Odrv4
    port map (
            O => \N__69015\,
            I => \c0.n9_adj_4341\
        );

    \I__17096\ : Odrv4
    port map (
            O => \N__69008\,
            I => \c0.n9_adj_4341\
        );

    \I__17095\ : Odrv12
    port map (
            O => \N__69005\,
            I => \c0.n9_adj_4341\
        );

    \I__17094\ : Odrv12
    port map (
            O => \N__69000\,
            I => \c0.n9_adj_4341\
        );

    \I__17093\ : InMux
    port map (
            O => \N__68989\,
            I => \N__68984\
        );

    \I__17092\ : InMux
    port map (
            O => \N__68988\,
            I => \N__68981\
        );

    \I__17091\ : InMux
    port map (
            O => \N__68987\,
            I => \N__68976\
        );

    \I__17090\ : LocalMux
    port map (
            O => \N__68984\,
            I => \N__68965\
        );

    \I__17089\ : LocalMux
    port map (
            O => \N__68981\,
            I => \N__68965\
        );

    \I__17088\ : InMux
    port map (
            O => \N__68980\,
            I => \N__68962\
        );

    \I__17087\ : InMux
    port map (
            O => \N__68979\,
            I => \N__68959\
        );

    \I__17086\ : LocalMux
    port map (
            O => \N__68976\,
            I => \N__68951\
        );

    \I__17085\ : InMux
    port map (
            O => \N__68975\,
            I => \N__68948\
        );

    \I__17084\ : InMux
    port map (
            O => \N__68974\,
            I => \N__68945\
        );

    \I__17083\ : CascadeMux
    port map (
            O => \N__68973\,
            I => \N__68941\
        );

    \I__17082\ : InMux
    port map (
            O => \N__68972\,
            I => \N__68935\
        );

    \I__17081\ : InMux
    port map (
            O => \N__68971\,
            I => \N__68932\
        );

    \I__17080\ : InMux
    port map (
            O => \N__68970\,
            I => \N__68929\
        );

    \I__17079\ : Span4Mux_v
    port map (
            O => \N__68965\,
            I => \N__68926\
        );

    \I__17078\ : LocalMux
    port map (
            O => \N__68962\,
            I => \N__68921\
        );

    \I__17077\ : LocalMux
    port map (
            O => \N__68959\,
            I => \N__68921\
        );

    \I__17076\ : InMux
    port map (
            O => \N__68958\,
            I => \N__68916\
        );

    \I__17075\ : InMux
    port map (
            O => \N__68957\,
            I => \N__68916\
        );

    \I__17074\ : InMux
    port map (
            O => \N__68956\,
            I => \N__68913\
        );

    \I__17073\ : InMux
    port map (
            O => \N__68955\,
            I => \N__68910\
        );

    \I__17072\ : InMux
    port map (
            O => \N__68954\,
            I => \N__68905\
        );

    \I__17071\ : Span4Mux_v
    port map (
            O => \N__68951\,
            I => \N__68900\
        );

    \I__17070\ : LocalMux
    port map (
            O => \N__68948\,
            I => \N__68900\
        );

    \I__17069\ : LocalMux
    port map (
            O => \N__68945\,
            I => \N__68897\
        );

    \I__17068\ : InMux
    port map (
            O => \N__68944\,
            I => \N__68894\
        );

    \I__17067\ : InMux
    port map (
            O => \N__68941\,
            I => \N__68889\
        );

    \I__17066\ : InMux
    port map (
            O => \N__68940\,
            I => \N__68889\
        );

    \I__17065\ : InMux
    port map (
            O => \N__68939\,
            I => \N__68884\
        );

    \I__17064\ : InMux
    port map (
            O => \N__68938\,
            I => \N__68884\
        );

    \I__17063\ : LocalMux
    port map (
            O => \N__68935\,
            I => \N__68877\
        );

    \I__17062\ : LocalMux
    port map (
            O => \N__68932\,
            I => \N__68873\
        );

    \I__17061\ : LocalMux
    port map (
            O => \N__68929\,
            I => \N__68868\
        );

    \I__17060\ : Span4Mux_h
    port map (
            O => \N__68926\,
            I => \N__68868\
        );

    \I__17059\ : Span4Mux_v
    port map (
            O => \N__68921\,
            I => \N__68862\
        );

    \I__17058\ : LocalMux
    port map (
            O => \N__68916\,
            I => \N__68855\
        );

    \I__17057\ : LocalMux
    port map (
            O => \N__68913\,
            I => \N__68855\
        );

    \I__17056\ : LocalMux
    port map (
            O => \N__68910\,
            I => \N__68855\
        );

    \I__17055\ : InMux
    port map (
            O => \N__68909\,
            I => \N__68852\
        );

    \I__17054\ : InMux
    port map (
            O => \N__68908\,
            I => \N__68849\
        );

    \I__17053\ : LocalMux
    port map (
            O => \N__68905\,
            I => \N__68846\
        );

    \I__17052\ : Span4Mux_h
    port map (
            O => \N__68900\,
            I => \N__68837\
        );

    \I__17051\ : Span4Mux_h
    port map (
            O => \N__68897\,
            I => \N__68837\
        );

    \I__17050\ : LocalMux
    port map (
            O => \N__68894\,
            I => \N__68837\
        );

    \I__17049\ : LocalMux
    port map (
            O => \N__68889\,
            I => \N__68837\
        );

    \I__17048\ : LocalMux
    port map (
            O => \N__68884\,
            I => \N__68834\
        );

    \I__17047\ : InMux
    port map (
            O => \N__68883\,
            I => \N__68831\
        );

    \I__17046\ : InMux
    port map (
            O => \N__68882\,
            I => \N__68826\
        );

    \I__17045\ : InMux
    port map (
            O => \N__68881\,
            I => \N__68826\
        );

    \I__17044\ : InMux
    port map (
            O => \N__68880\,
            I => \N__68823\
        );

    \I__17043\ : Span4Mux_h
    port map (
            O => \N__68877\,
            I => \N__68820\
        );

    \I__17042\ : InMux
    port map (
            O => \N__68876\,
            I => \N__68817\
        );

    \I__17041\ : Span4Mux_v
    port map (
            O => \N__68873\,
            I => \N__68812\
        );

    \I__17040\ : Span4Mux_v
    port map (
            O => \N__68868\,
            I => \N__68812\
        );

    \I__17039\ : InMux
    port map (
            O => \N__68867\,
            I => \N__68809\
        );

    \I__17038\ : InMux
    port map (
            O => \N__68866\,
            I => \N__68806\
        );

    \I__17037\ : InMux
    port map (
            O => \N__68865\,
            I => \N__68803\
        );

    \I__17036\ : Span4Mux_h
    port map (
            O => \N__68862\,
            I => \N__68800\
        );

    \I__17035\ : Span4Mux_v
    port map (
            O => \N__68855\,
            I => \N__68797\
        );

    \I__17034\ : LocalMux
    port map (
            O => \N__68852\,
            I => \N__68792\
        );

    \I__17033\ : LocalMux
    port map (
            O => \N__68849\,
            I => \N__68792\
        );

    \I__17032\ : Span4Mux_h
    port map (
            O => \N__68846\,
            I => \N__68789\
        );

    \I__17031\ : Span4Mux_v
    port map (
            O => \N__68837\,
            I => \N__68786\
        );

    \I__17030\ : Span4Mux_v
    port map (
            O => \N__68834\,
            I => \N__68781\
        );

    \I__17029\ : LocalMux
    port map (
            O => \N__68831\,
            I => \N__68776\
        );

    \I__17028\ : LocalMux
    port map (
            O => \N__68826\,
            I => \N__68776\
        );

    \I__17027\ : LocalMux
    port map (
            O => \N__68823\,
            I => \N__68771\
        );

    \I__17026\ : Span4Mux_v
    port map (
            O => \N__68820\,
            I => \N__68771\
        );

    \I__17025\ : LocalMux
    port map (
            O => \N__68817\,
            I => \N__68766\
        );

    \I__17024\ : Span4Mux_v
    port map (
            O => \N__68812\,
            I => \N__68766\
        );

    \I__17023\ : LocalMux
    port map (
            O => \N__68809\,
            I => \N__68763\
        );

    \I__17022\ : LocalMux
    port map (
            O => \N__68806\,
            I => \N__68756\
        );

    \I__17021\ : LocalMux
    port map (
            O => \N__68803\,
            I => \N__68756\
        );

    \I__17020\ : Sp12to4
    port map (
            O => \N__68800\,
            I => \N__68756\
        );

    \I__17019\ : Sp12to4
    port map (
            O => \N__68797\,
            I => \N__68753\
        );

    \I__17018\ : Span4Mux_h
    port map (
            O => \N__68792\,
            I => \N__68746\
        );

    \I__17017\ : Span4Mux_v
    port map (
            O => \N__68789\,
            I => \N__68746\
        );

    \I__17016\ : Span4Mux_h
    port map (
            O => \N__68786\,
            I => \N__68746\
        );

    \I__17015\ : InMux
    port map (
            O => \N__68785\,
            I => \N__68743\
        );

    \I__17014\ : InMux
    port map (
            O => \N__68784\,
            I => \N__68740\
        );

    \I__17013\ : Span4Mux_h
    port map (
            O => \N__68781\,
            I => \N__68731\
        );

    \I__17012\ : Span4Mux_v
    port map (
            O => \N__68776\,
            I => \N__68731\
        );

    \I__17011\ : Span4Mux_h
    port map (
            O => \N__68771\,
            I => \N__68731\
        );

    \I__17010\ : Span4Mux_v
    port map (
            O => \N__68766\,
            I => \N__68731\
        );

    \I__17009\ : Span12Mux_s11_v
    port map (
            O => \N__68763\,
            I => \N__68722\
        );

    \I__17008\ : Span12Mux_s10_h
    port map (
            O => \N__68756\,
            I => \N__68722\
        );

    \I__17007\ : Span12Mux_h
    port map (
            O => \N__68753\,
            I => \N__68722\
        );

    \I__17006\ : Sp12to4
    port map (
            O => \N__68746\,
            I => \N__68722\
        );

    \I__17005\ : LocalMux
    port map (
            O => \N__68743\,
            I => rx_data_7
        );

    \I__17004\ : LocalMux
    port map (
            O => \N__68740\,
            I => rx_data_7
        );

    \I__17003\ : Odrv4
    port map (
            O => \N__68731\,
            I => rx_data_7
        );

    \I__17002\ : Odrv12
    port map (
            O => \N__68722\,
            I => rx_data_7
        );

    \I__17001\ : CascadeMux
    port map (
            O => \N__68713\,
            I => \N__68709\
        );

    \I__17000\ : InMux
    port map (
            O => \N__68712\,
            I => \N__68706\
        );

    \I__16999\ : InMux
    port map (
            O => \N__68709\,
            I => \N__68702\
        );

    \I__16998\ : LocalMux
    port map (
            O => \N__68706\,
            I => \N__68699\
        );

    \I__16997\ : CascadeMux
    port map (
            O => \N__68705\,
            I => \N__68696\
        );

    \I__16996\ : LocalMux
    port map (
            O => \N__68702\,
            I => \N__68690\
        );

    \I__16995\ : Span4Mux_h
    port map (
            O => \N__68699\,
            I => \N__68690\
        );

    \I__16994\ : InMux
    port map (
            O => \N__68696\,
            I => \N__68685\
        );

    \I__16993\ : InMux
    port map (
            O => \N__68695\,
            I => \N__68685\
        );

    \I__16992\ : Odrv4
    port map (
            O => \N__68690\,
            I => \c0.data_in_frame_26_7\
        );

    \I__16991\ : LocalMux
    port map (
            O => \N__68685\,
            I => \c0.data_in_frame_26_7\
        );

    \I__16990\ : CascadeMux
    port map (
            O => \N__68680\,
            I => \N__68675\
        );

    \I__16989\ : CascadeMux
    port map (
            O => \N__68679\,
            I => \N__68666\
        );

    \I__16988\ : InMux
    port map (
            O => \N__68678\,
            I => \N__68663\
        );

    \I__16987\ : InMux
    port map (
            O => \N__68675\,
            I => \N__68660\
        );

    \I__16986\ : InMux
    port map (
            O => \N__68674\,
            I => \N__68655\
        );

    \I__16985\ : InMux
    port map (
            O => \N__68673\,
            I => \N__68650\
        );

    \I__16984\ : InMux
    port map (
            O => \N__68672\,
            I => \N__68650\
        );

    \I__16983\ : CascadeMux
    port map (
            O => \N__68671\,
            I => \N__68647\
        );

    \I__16982\ : InMux
    port map (
            O => \N__68670\,
            I => \N__68644\
        );

    \I__16981\ : InMux
    port map (
            O => \N__68669\,
            I => \N__68639\
        );

    \I__16980\ : InMux
    port map (
            O => \N__68666\,
            I => \N__68639\
        );

    \I__16979\ : LocalMux
    port map (
            O => \N__68663\,
            I => \N__68633\
        );

    \I__16978\ : LocalMux
    port map (
            O => \N__68660\,
            I => \N__68633\
        );

    \I__16977\ : CascadeMux
    port map (
            O => \N__68659\,
            I => \N__68629\
        );

    \I__16976\ : CascadeMux
    port map (
            O => \N__68658\,
            I => \N__68625\
        );

    \I__16975\ : LocalMux
    port map (
            O => \N__68655\,
            I => \N__68620\
        );

    \I__16974\ : LocalMux
    port map (
            O => \N__68650\,
            I => \N__68620\
        );

    \I__16973\ : InMux
    port map (
            O => \N__68647\,
            I => \N__68617\
        );

    \I__16972\ : LocalMux
    port map (
            O => \N__68644\,
            I => \N__68614\
        );

    \I__16971\ : LocalMux
    port map (
            O => \N__68639\,
            I => \N__68611\
        );

    \I__16970\ : InMux
    port map (
            O => \N__68638\,
            I => \N__68608\
        );

    \I__16969\ : Span4Mux_v
    port map (
            O => \N__68633\,
            I => \N__68605\
        );

    \I__16968\ : InMux
    port map (
            O => \N__68632\,
            I => \N__68602\
        );

    \I__16967\ : InMux
    port map (
            O => \N__68629\,
            I => \N__68595\
        );

    \I__16966\ : InMux
    port map (
            O => \N__68628\,
            I => \N__68595\
        );

    \I__16965\ : InMux
    port map (
            O => \N__68625\,
            I => \N__68592\
        );

    \I__16964\ : Span4Mux_h
    port map (
            O => \N__68620\,
            I => \N__68584\
        );

    \I__16963\ : LocalMux
    port map (
            O => \N__68617\,
            I => \N__68584\
        );

    \I__16962\ : Span4Mux_h
    port map (
            O => \N__68614\,
            I => \N__68579\
        );

    \I__16961\ : Span4Mux_v
    port map (
            O => \N__68611\,
            I => \N__68579\
        );

    \I__16960\ : LocalMux
    port map (
            O => \N__68608\,
            I => \N__68576\
        );

    \I__16959\ : Span4Mux_h
    port map (
            O => \N__68605\,
            I => \N__68571\
        );

    \I__16958\ : LocalMux
    port map (
            O => \N__68602\,
            I => \N__68571\
        );

    \I__16957\ : InMux
    port map (
            O => \N__68601\,
            I => \N__68565\
        );

    \I__16956\ : InMux
    port map (
            O => \N__68600\,
            I => \N__68562\
        );

    \I__16955\ : LocalMux
    port map (
            O => \N__68595\,
            I => \N__68557\
        );

    \I__16954\ : LocalMux
    port map (
            O => \N__68592\,
            I => \N__68557\
        );

    \I__16953\ : InMux
    port map (
            O => \N__68591\,
            I => \N__68554\
        );

    \I__16952\ : CascadeMux
    port map (
            O => \N__68590\,
            I => \N__68549\
        );

    \I__16951\ : InMux
    port map (
            O => \N__68589\,
            I => \N__68546\
        );

    \I__16950\ : Span4Mux_h
    port map (
            O => \N__68584\,
            I => \N__68542\
        );

    \I__16949\ : Span4Mux_h
    port map (
            O => \N__68579\,
            I => \N__68539\
        );

    \I__16948\ : Span4Mux_h
    port map (
            O => \N__68576\,
            I => \N__68536\
        );

    \I__16947\ : Span4Mux_v
    port map (
            O => \N__68571\,
            I => \N__68533\
        );

    \I__16946\ : InMux
    port map (
            O => \N__68570\,
            I => \N__68530\
        );

    \I__16945\ : InMux
    port map (
            O => \N__68569\,
            I => \N__68527\
        );

    \I__16944\ : InMux
    port map (
            O => \N__68568\,
            I => \N__68524\
        );

    \I__16943\ : LocalMux
    port map (
            O => \N__68565\,
            I => \N__68517\
        );

    \I__16942\ : LocalMux
    port map (
            O => \N__68562\,
            I => \N__68517\
        );

    \I__16941\ : Span4Mux_v
    port map (
            O => \N__68557\,
            I => \N__68517\
        );

    \I__16940\ : LocalMux
    port map (
            O => \N__68554\,
            I => \N__68513\
        );

    \I__16939\ : InMux
    port map (
            O => \N__68553\,
            I => \N__68506\
        );

    \I__16938\ : InMux
    port map (
            O => \N__68552\,
            I => \N__68506\
        );

    \I__16937\ : InMux
    port map (
            O => \N__68549\,
            I => \N__68506\
        );

    \I__16936\ : LocalMux
    port map (
            O => \N__68546\,
            I => \N__68503\
        );

    \I__16935\ : InMux
    port map (
            O => \N__68545\,
            I => \N__68500\
        );

    \I__16934\ : Span4Mux_h
    port map (
            O => \N__68542\,
            I => \N__68493\
        );

    \I__16933\ : Span4Mux_h
    port map (
            O => \N__68539\,
            I => \N__68493\
        );

    \I__16932\ : Span4Mux_v
    port map (
            O => \N__68536\,
            I => \N__68493\
        );

    \I__16931\ : Sp12to4
    port map (
            O => \N__68533\,
            I => \N__68488\
        );

    \I__16930\ : LocalMux
    port map (
            O => \N__68530\,
            I => \N__68488\
        );

    \I__16929\ : LocalMux
    port map (
            O => \N__68527\,
            I => \N__68485\
        );

    \I__16928\ : LocalMux
    port map (
            O => \N__68524\,
            I => \N__68480\
        );

    \I__16927\ : Span4Mux_v
    port map (
            O => \N__68517\,
            I => \N__68480\
        );

    \I__16926\ : InMux
    port map (
            O => \N__68516\,
            I => \N__68477\
        );

    \I__16925\ : Sp12to4
    port map (
            O => \N__68513\,
            I => \N__68468\
        );

    \I__16924\ : LocalMux
    port map (
            O => \N__68506\,
            I => \N__68468\
        );

    \I__16923\ : Span12Mux_v
    port map (
            O => \N__68503\,
            I => \N__68468\
        );

    \I__16922\ : LocalMux
    port map (
            O => \N__68500\,
            I => \N__68468\
        );

    \I__16921\ : Sp12to4
    port map (
            O => \N__68493\,
            I => \N__68463\
        );

    \I__16920\ : Span12Mux_h
    port map (
            O => \N__68488\,
            I => \N__68463\
        );

    \I__16919\ : Span4Mux_v
    port map (
            O => \N__68485\,
            I => \N__68460\
        );

    \I__16918\ : Span4Mux_h
    port map (
            O => \N__68480\,
            I => \N__68457\
        );

    \I__16917\ : LocalMux
    port map (
            O => \N__68477\,
            I => \N__68450\
        );

    \I__16916\ : Span12Mux_v
    port map (
            O => \N__68468\,
            I => \N__68450\
        );

    \I__16915\ : Span12Mux_v
    port map (
            O => \N__68463\,
            I => \N__68450\
        );

    \I__16914\ : Odrv4
    port map (
            O => \N__68460\,
            I => \c0.n17596\
        );

    \I__16913\ : Odrv4
    port map (
            O => \N__68457\,
            I => \c0.n17596\
        );

    \I__16912\ : Odrv12
    port map (
            O => \N__68450\,
            I => \c0.n17596\
        );

    \I__16911\ : InMux
    port map (
            O => \N__68443\,
            I => \N__68438\
        );

    \I__16910\ : CascadeMux
    port map (
            O => \N__68442\,
            I => \N__68430\
        );

    \I__16909\ : CascadeMux
    port map (
            O => \N__68441\,
            I => \N__68427\
        );

    \I__16908\ : LocalMux
    port map (
            O => \N__68438\,
            I => \N__68423\
        );

    \I__16907\ : InMux
    port map (
            O => \N__68437\,
            I => \N__68420\
        );

    \I__16906\ : CascadeMux
    port map (
            O => \N__68436\,
            I => \N__68413\
        );

    \I__16905\ : InMux
    port map (
            O => \N__68435\,
            I => \N__68407\
        );

    \I__16904\ : InMux
    port map (
            O => \N__68434\,
            I => \N__68404\
        );

    \I__16903\ : InMux
    port map (
            O => \N__68433\,
            I => \N__68399\
        );

    \I__16902\ : InMux
    port map (
            O => \N__68430\,
            I => \N__68399\
        );

    \I__16901\ : InMux
    port map (
            O => \N__68427\,
            I => \N__68396\
        );

    \I__16900\ : InMux
    port map (
            O => \N__68426\,
            I => \N__68390\
        );

    \I__16899\ : Span4Mux_v
    port map (
            O => \N__68423\,
            I => \N__68385\
        );

    \I__16898\ : LocalMux
    port map (
            O => \N__68420\,
            I => \N__68385\
        );

    \I__16897\ : InMux
    port map (
            O => \N__68419\,
            I => \N__68378\
        );

    \I__16896\ : InMux
    port map (
            O => \N__68418\,
            I => \N__68378\
        );

    \I__16895\ : InMux
    port map (
            O => \N__68417\,
            I => \N__68378\
        );

    \I__16894\ : InMux
    port map (
            O => \N__68416\,
            I => \N__68374\
        );

    \I__16893\ : InMux
    port map (
            O => \N__68413\,
            I => \N__68370\
        );

    \I__16892\ : InMux
    port map (
            O => \N__68412\,
            I => \N__68366\
        );

    \I__16891\ : CascadeMux
    port map (
            O => \N__68411\,
            I => \N__68363\
        );

    \I__16890\ : InMux
    port map (
            O => \N__68410\,
            I => \N__68360\
        );

    \I__16889\ : LocalMux
    port map (
            O => \N__68407\,
            I => \N__68349\
        );

    \I__16888\ : LocalMux
    port map (
            O => \N__68404\,
            I => \N__68346\
        );

    \I__16887\ : LocalMux
    port map (
            O => \N__68399\,
            I => \N__68341\
        );

    \I__16886\ : LocalMux
    port map (
            O => \N__68396\,
            I => \N__68341\
        );

    \I__16885\ : InMux
    port map (
            O => \N__68395\,
            I => \N__68338\
        );

    \I__16884\ : InMux
    port map (
            O => \N__68394\,
            I => \N__68333\
        );

    \I__16883\ : InMux
    port map (
            O => \N__68393\,
            I => \N__68333\
        );

    \I__16882\ : LocalMux
    port map (
            O => \N__68390\,
            I => \N__68330\
        );

    \I__16881\ : Span4Mux_h
    port map (
            O => \N__68385\,
            I => \N__68325\
        );

    \I__16880\ : LocalMux
    port map (
            O => \N__68378\,
            I => \N__68325\
        );

    \I__16879\ : InMux
    port map (
            O => \N__68377\,
            I => \N__68322\
        );

    \I__16878\ : LocalMux
    port map (
            O => \N__68374\,
            I => \N__68319\
        );

    \I__16877\ : InMux
    port map (
            O => \N__68373\,
            I => \N__68316\
        );

    \I__16876\ : LocalMux
    port map (
            O => \N__68370\,
            I => \N__68313\
        );

    \I__16875\ : InMux
    port map (
            O => \N__68369\,
            I => \N__68310\
        );

    \I__16874\ : LocalMux
    port map (
            O => \N__68366\,
            I => \N__68307\
        );

    \I__16873\ : InMux
    port map (
            O => \N__68363\,
            I => \N__68304\
        );

    \I__16872\ : LocalMux
    port map (
            O => \N__68360\,
            I => \N__68301\
        );

    \I__16871\ : InMux
    port map (
            O => \N__68359\,
            I => \N__68296\
        );

    \I__16870\ : InMux
    port map (
            O => \N__68358\,
            I => \N__68296\
        );

    \I__16869\ : InMux
    port map (
            O => \N__68357\,
            I => \N__68293\
        );

    \I__16868\ : InMux
    port map (
            O => \N__68356\,
            I => \N__68290\
        );

    \I__16867\ : InMux
    port map (
            O => \N__68355\,
            I => \N__68285\
        );

    \I__16866\ : InMux
    port map (
            O => \N__68354\,
            I => \N__68280\
        );

    \I__16865\ : InMux
    port map (
            O => \N__68353\,
            I => \N__68280\
        );

    \I__16864\ : InMux
    port map (
            O => \N__68352\,
            I => \N__68277\
        );

    \I__16863\ : Span4Mux_v
    port map (
            O => \N__68349\,
            I => \N__68274\
        );

    \I__16862\ : Span4Mux_h
    port map (
            O => \N__68346\,
            I => \N__68269\
        );

    \I__16861\ : Span4Mux_v
    port map (
            O => \N__68341\,
            I => \N__68269\
        );

    \I__16860\ : LocalMux
    port map (
            O => \N__68338\,
            I => \N__68262\
        );

    \I__16859\ : LocalMux
    port map (
            O => \N__68333\,
            I => \N__68262\
        );

    \I__16858\ : Span4Mux_v
    port map (
            O => \N__68330\,
            I => \N__68262\
        );

    \I__16857\ : Span4Mux_v
    port map (
            O => \N__68325\,
            I => \N__68259\
        );

    \I__16856\ : LocalMux
    port map (
            O => \N__68322\,
            I => \N__68256\
        );

    \I__16855\ : Span4Mux_h
    port map (
            O => \N__68319\,
            I => \N__68251\
        );

    \I__16854\ : LocalMux
    port map (
            O => \N__68316\,
            I => \N__68251\
        );

    \I__16853\ : Span4Mux_v
    port map (
            O => \N__68313\,
            I => \N__68248\
        );

    \I__16852\ : LocalMux
    port map (
            O => \N__68310\,
            I => \N__68243\
        );

    \I__16851\ : Span4Mux_v
    port map (
            O => \N__68307\,
            I => \N__68243\
        );

    \I__16850\ : LocalMux
    port map (
            O => \N__68304\,
            I => \N__68238\
        );

    \I__16849\ : Span4Mux_v
    port map (
            O => \N__68301\,
            I => \N__68238\
        );

    \I__16848\ : LocalMux
    port map (
            O => \N__68296\,
            I => \N__68235\
        );

    \I__16847\ : LocalMux
    port map (
            O => \N__68293\,
            I => \N__68230\
        );

    \I__16846\ : LocalMux
    port map (
            O => \N__68290\,
            I => \N__68230\
        );

    \I__16845\ : InMux
    port map (
            O => \N__68289\,
            I => \N__68227\
        );

    \I__16844\ : InMux
    port map (
            O => \N__68288\,
            I => \N__68224\
        );

    \I__16843\ : LocalMux
    port map (
            O => \N__68285\,
            I => \N__68219\
        );

    \I__16842\ : LocalMux
    port map (
            O => \N__68280\,
            I => \N__68219\
        );

    \I__16841\ : LocalMux
    port map (
            O => \N__68277\,
            I => \N__68216\
        );

    \I__16840\ : Span4Mux_v
    port map (
            O => \N__68274\,
            I => \N__68211\
        );

    \I__16839\ : Span4Mux_v
    port map (
            O => \N__68269\,
            I => \N__68211\
        );

    \I__16838\ : Span4Mux_v
    port map (
            O => \N__68262\,
            I => \N__68208\
        );

    \I__16837\ : Span4Mux_h
    port map (
            O => \N__68259\,
            I => \N__68205\
        );

    \I__16836\ : Span4Mux_v
    port map (
            O => \N__68256\,
            I => \N__68196\
        );

    \I__16835\ : Span4Mux_v
    port map (
            O => \N__68251\,
            I => \N__68196\
        );

    \I__16834\ : Span4Mux_h
    port map (
            O => \N__68248\,
            I => \N__68196\
        );

    \I__16833\ : Span4Mux_v
    port map (
            O => \N__68243\,
            I => \N__68196\
        );

    \I__16832\ : Span4Mux_v
    port map (
            O => \N__68238\,
            I => \N__68189\
        );

    \I__16831\ : Span4Mux_v
    port map (
            O => \N__68235\,
            I => \N__68189\
        );

    \I__16830\ : Span4Mux_h
    port map (
            O => \N__68230\,
            I => \N__68189\
        );

    \I__16829\ : LocalMux
    port map (
            O => \N__68227\,
            I => \N__68178\
        );

    \I__16828\ : LocalMux
    port map (
            O => \N__68224\,
            I => \N__68178\
        );

    \I__16827\ : Span12Mux_v
    port map (
            O => \N__68219\,
            I => \N__68178\
        );

    \I__16826\ : Span12Mux_v
    port map (
            O => \N__68216\,
            I => \N__68178\
        );

    \I__16825\ : Sp12to4
    port map (
            O => \N__68211\,
            I => \N__68178\
        );

    \I__16824\ : Odrv4
    port map (
            O => \N__68208\,
            I => rx_data_2
        );

    \I__16823\ : Odrv4
    port map (
            O => \N__68205\,
            I => rx_data_2
        );

    \I__16822\ : Odrv4
    port map (
            O => \N__68196\,
            I => rx_data_2
        );

    \I__16821\ : Odrv4
    port map (
            O => \N__68189\,
            I => rx_data_2
        );

    \I__16820\ : Odrv12
    port map (
            O => \N__68178\,
            I => rx_data_2
        );

    \I__16819\ : InMux
    port map (
            O => \N__68167\,
            I => \N__68152\
        );

    \I__16818\ : InMux
    port map (
            O => \N__68166\,
            I => \N__68149\
        );

    \I__16817\ : InMux
    port map (
            O => \N__68165\,
            I => \N__68132\
        );

    \I__16816\ : CascadeMux
    port map (
            O => \N__68164\,
            I => \N__68129\
        );

    \I__16815\ : InMux
    port map (
            O => \N__68163\,
            I => \N__68122\
        );

    \I__16814\ : InMux
    port map (
            O => \N__68162\,
            I => \N__68122\
        );

    \I__16813\ : InMux
    port map (
            O => \N__68161\,
            I => \N__68122\
        );

    \I__16812\ : InMux
    port map (
            O => \N__68160\,
            I => \N__68117\
        );

    \I__16811\ : InMux
    port map (
            O => \N__68159\,
            I => \N__68117\
        );

    \I__16810\ : InMux
    port map (
            O => \N__68158\,
            I => \N__68112\
        );

    \I__16809\ : InMux
    port map (
            O => \N__68157\,
            I => \N__68112\
        );

    \I__16808\ : InMux
    port map (
            O => \N__68156\,
            I => \N__68104\
        );

    \I__16807\ : InMux
    port map (
            O => \N__68155\,
            I => \N__68104\
        );

    \I__16806\ : LocalMux
    port map (
            O => \N__68152\,
            I => \N__68101\
        );

    \I__16805\ : LocalMux
    port map (
            O => \N__68149\,
            I => \N__68098\
        );

    \I__16804\ : InMux
    port map (
            O => \N__68148\,
            I => \N__68088\
        );

    \I__16803\ : CascadeMux
    port map (
            O => \N__68147\,
            I => \N__68083\
        );

    \I__16802\ : InMux
    port map (
            O => \N__68146\,
            I => \N__68078\
        );

    \I__16801\ : InMux
    port map (
            O => \N__68145\,
            I => \N__68078\
        );

    \I__16800\ : InMux
    port map (
            O => \N__68144\,
            I => \N__68071\
        );

    \I__16799\ : InMux
    port map (
            O => \N__68143\,
            I => \N__68071\
        );

    \I__16798\ : InMux
    port map (
            O => \N__68142\,
            I => \N__68071\
        );

    \I__16797\ : InMux
    port map (
            O => \N__68141\,
            I => \N__68062\
        );

    \I__16796\ : InMux
    port map (
            O => \N__68140\,
            I => \N__68057\
        );

    \I__16795\ : InMux
    port map (
            O => \N__68139\,
            I => \N__68057\
        );

    \I__16794\ : InMux
    port map (
            O => \N__68138\,
            I => \N__68048\
        );

    \I__16793\ : InMux
    port map (
            O => \N__68137\,
            I => \N__68048\
        );

    \I__16792\ : InMux
    port map (
            O => \N__68136\,
            I => \N__68048\
        );

    \I__16791\ : InMux
    port map (
            O => \N__68135\,
            I => \N__68048\
        );

    \I__16790\ : LocalMux
    port map (
            O => \N__68132\,
            I => \N__68045\
        );

    \I__16789\ : InMux
    port map (
            O => \N__68129\,
            I => \N__68039\
        );

    \I__16788\ : LocalMux
    port map (
            O => \N__68122\,
            I => \N__68036\
        );

    \I__16787\ : LocalMux
    port map (
            O => \N__68117\,
            I => \N__68033\
        );

    \I__16786\ : LocalMux
    port map (
            O => \N__68112\,
            I => \N__68030\
        );

    \I__16785\ : InMux
    port map (
            O => \N__68111\,
            I => \N__68023\
        );

    \I__16784\ : InMux
    port map (
            O => \N__68110\,
            I => \N__68023\
        );

    \I__16783\ : InMux
    port map (
            O => \N__68109\,
            I => \N__68023\
        );

    \I__16782\ : LocalMux
    port map (
            O => \N__68104\,
            I => \N__68020\
        );

    \I__16781\ : Span4Mux_v
    port map (
            O => \N__68101\,
            I => \N__68012\
        );

    \I__16780\ : Span4Mux_h
    port map (
            O => \N__68098\,
            I => \N__68012\
        );

    \I__16779\ : InMux
    port map (
            O => \N__68097\,
            I => \N__68009\
        );

    \I__16778\ : InMux
    port map (
            O => \N__68096\,
            I => \N__68003\
        );

    \I__16777\ : InMux
    port map (
            O => \N__68095\,
            I => \N__68000\
        );

    \I__16776\ : InMux
    port map (
            O => \N__68094\,
            I => \N__67995\
        );

    \I__16775\ : InMux
    port map (
            O => \N__68093\,
            I => \N__67995\
        );

    \I__16774\ : InMux
    port map (
            O => \N__68092\,
            I => \N__67990\
        );

    \I__16773\ : InMux
    port map (
            O => \N__68091\,
            I => \N__67990\
        );

    \I__16772\ : LocalMux
    port map (
            O => \N__68088\,
            I => \N__67987\
        );

    \I__16771\ : InMux
    port map (
            O => \N__68087\,
            I => \N__67984\
        );

    \I__16770\ : InMux
    port map (
            O => \N__68086\,
            I => \N__67979\
        );

    \I__16769\ : InMux
    port map (
            O => \N__68083\,
            I => \N__67979\
        );

    \I__16768\ : LocalMux
    port map (
            O => \N__68078\,
            I => \N__67974\
        );

    \I__16767\ : LocalMux
    port map (
            O => \N__68071\,
            I => \N__67974\
        );

    \I__16766\ : InMux
    port map (
            O => \N__68070\,
            I => \N__67971\
        );

    \I__16765\ : InMux
    port map (
            O => \N__68069\,
            I => \N__67966\
        );

    \I__16764\ : InMux
    port map (
            O => \N__68068\,
            I => \N__67966\
        );

    \I__16763\ : InMux
    port map (
            O => \N__68067\,
            I => \N__67959\
        );

    \I__16762\ : InMux
    port map (
            O => \N__68066\,
            I => \N__67959\
        );

    \I__16761\ : InMux
    port map (
            O => \N__68065\,
            I => \N__67959\
        );

    \I__16760\ : LocalMux
    port map (
            O => \N__68062\,
            I => \N__67954\
        );

    \I__16759\ : LocalMux
    port map (
            O => \N__68057\,
            I => \N__67954\
        );

    \I__16758\ : LocalMux
    port map (
            O => \N__68048\,
            I => \N__67949\
        );

    \I__16757\ : Span4Mux_v
    port map (
            O => \N__68045\,
            I => \N__67949\
        );

    \I__16756\ : CascadeMux
    port map (
            O => \N__68044\,
            I => \N__67946\
        );

    \I__16755\ : InMux
    port map (
            O => \N__68043\,
            I => \N__67941\
        );

    \I__16754\ : InMux
    port map (
            O => \N__68042\,
            I => \N__67941\
        );

    \I__16753\ : LocalMux
    port map (
            O => \N__68039\,
            I => \N__67938\
        );

    \I__16752\ : Span4Mux_v
    port map (
            O => \N__68036\,
            I => \N__67933\
        );

    \I__16751\ : Span4Mux_v
    port map (
            O => \N__68033\,
            I => \N__67933\
        );

    \I__16750\ : Span4Mux_h
    port map (
            O => \N__68030\,
            I => \N__67926\
        );

    \I__16749\ : LocalMux
    port map (
            O => \N__68023\,
            I => \N__67926\
        );

    \I__16748\ : Span4Mux_v
    port map (
            O => \N__68020\,
            I => \N__67926\
        );

    \I__16747\ : InMux
    port map (
            O => \N__68019\,
            I => \N__67919\
        );

    \I__16746\ : InMux
    port map (
            O => \N__68018\,
            I => \N__67919\
        );

    \I__16745\ : InMux
    port map (
            O => \N__68017\,
            I => \N__67919\
        );

    \I__16744\ : Span4Mux_h
    port map (
            O => \N__68012\,
            I => \N__67916\
        );

    \I__16743\ : LocalMux
    port map (
            O => \N__68009\,
            I => \N__67913\
        );

    \I__16742\ : InMux
    port map (
            O => \N__68008\,
            I => \N__67904\
        );

    \I__16741\ : InMux
    port map (
            O => \N__68007\,
            I => \N__67904\
        );

    \I__16740\ : InMux
    port map (
            O => \N__68006\,
            I => \N__67904\
        );

    \I__16739\ : LocalMux
    port map (
            O => \N__68003\,
            I => \N__67901\
        );

    \I__16738\ : LocalMux
    port map (
            O => \N__68000\,
            I => \N__67892\
        );

    \I__16737\ : LocalMux
    port map (
            O => \N__67995\,
            I => \N__67892\
        );

    \I__16736\ : LocalMux
    port map (
            O => \N__67990\,
            I => \N__67892\
        );

    \I__16735\ : Span4Mux_h
    port map (
            O => \N__67987\,
            I => \N__67892\
        );

    \I__16734\ : LocalMux
    port map (
            O => \N__67984\,
            I => \N__67885\
        );

    \I__16733\ : LocalMux
    port map (
            O => \N__67979\,
            I => \N__67885\
        );

    \I__16732\ : Span4Mux_v
    port map (
            O => \N__67974\,
            I => \N__67885\
        );

    \I__16731\ : LocalMux
    port map (
            O => \N__67971\,
            I => \N__67874\
        );

    \I__16730\ : LocalMux
    port map (
            O => \N__67966\,
            I => \N__67874\
        );

    \I__16729\ : LocalMux
    port map (
            O => \N__67959\,
            I => \N__67874\
        );

    \I__16728\ : Span4Mux_v
    port map (
            O => \N__67954\,
            I => \N__67874\
        );

    \I__16727\ : Span4Mux_h
    port map (
            O => \N__67949\,
            I => \N__67874\
        );

    \I__16726\ : InMux
    port map (
            O => \N__67946\,
            I => \N__67871\
        );

    \I__16725\ : LocalMux
    port map (
            O => \N__67941\,
            I => \N__67866\
        );

    \I__16724\ : Span4Mux_v
    port map (
            O => \N__67938\,
            I => \N__67866\
        );

    \I__16723\ : Span4Mux_v
    port map (
            O => \N__67933\,
            I => \N__67861\
        );

    \I__16722\ : Span4Mux_v
    port map (
            O => \N__67926\,
            I => \N__67861\
        );

    \I__16721\ : LocalMux
    port map (
            O => \N__67919\,
            I => \N__67854\
        );

    \I__16720\ : Span4Mux_v
    port map (
            O => \N__67916\,
            I => \N__67854\
        );

    \I__16719\ : Span4Mux_h
    port map (
            O => \N__67913\,
            I => \N__67854\
        );

    \I__16718\ : InMux
    port map (
            O => \N__67912\,
            I => \N__67849\
        );

    \I__16717\ : InMux
    port map (
            O => \N__67911\,
            I => \N__67849\
        );

    \I__16716\ : LocalMux
    port map (
            O => \N__67904\,
            I => \N__67838\
        );

    \I__16715\ : Span4Mux_v
    port map (
            O => \N__67901\,
            I => \N__67838\
        );

    \I__16714\ : Span4Mux_v
    port map (
            O => \N__67892\,
            I => \N__67838\
        );

    \I__16713\ : Span4Mux_h
    port map (
            O => \N__67885\,
            I => \N__67838\
        );

    \I__16712\ : Span4Mux_v
    port map (
            O => \N__67874\,
            I => \N__67838\
        );

    \I__16711\ : LocalMux
    port map (
            O => \N__67871\,
            I => \N__67831\
        );

    \I__16710\ : Span4Mux_h
    port map (
            O => \N__67866\,
            I => \N__67831\
        );

    \I__16709\ : Span4Mux_h
    port map (
            O => \N__67861\,
            I => \N__67831\
        );

    \I__16708\ : Span4Mux_v
    port map (
            O => \N__67854\,
            I => \N__67828\
        );

    \I__16707\ : LocalMux
    port map (
            O => \N__67849\,
            I => \c0.n21758\
        );

    \I__16706\ : Odrv4
    port map (
            O => \N__67838\,
            I => \c0.n21758\
        );

    \I__16705\ : Odrv4
    port map (
            O => \N__67831\,
            I => \c0.n21758\
        );

    \I__16704\ : Odrv4
    port map (
            O => \N__67828\,
            I => \c0.n21758\
        );

    \I__16703\ : CascadeMux
    port map (
            O => \N__67819\,
            I => \N__67815\
        );

    \I__16702\ : InMux
    port map (
            O => \N__67818\,
            I => \N__67812\
        );

    \I__16701\ : InMux
    port map (
            O => \N__67815\,
            I => \N__67808\
        );

    \I__16700\ : LocalMux
    port map (
            O => \N__67812\,
            I => \N__67805\
        );

    \I__16699\ : InMux
    port map (
            O => \N__67811\,
            I => \N__67802\
        );

    \I__16698\ : LocalMux
    port map (
            O => \N__67808\,
            I => \c0.data_in_frame_23_2\
        );

    \I__16697\ : Odrv12
    port map (
            O => \N__67805\,
            I => \c0.data_in_frame_23_2\
        );

    \I__16696\ : LocalMux
    port map (
            O => \N__67802\,
            I => \c0.data_in_frame_23_2\
        );

    \I__16695\ : InMux
    port map (
            O => \N__67795\,
            I => \N__67784\
        );

    \I__16694\ : InMux
    port map (
            O => \N__67794\,
            I => \N__67784\
        );

    \I__16693\ : InMux
    port map (
            O => \N__67793\,
            I => \N__67784\
        );

    \I__16692\ : InMux
    port map (
            O => \N__67792\,
            I => \N__67779\
        );

    \I__16691\ : InMux
    port map (
            O => \N__67791\,
            I => \N__67779\
        );

    \I__16690\ : LocalMux
    port map (
            O => \N__67784\,
            I => \N__67770\
        );

    \I__16689\ : LocalMux
    port map (
            O => \N__67779\,
            I => \N__67770\
        );

    \I__16688\ : InMux
    port map (
            O => \N__67778\,
            I => \N__67765\
        );

    \I__16687\ : InMux
    port map (
            O => \N__67777\,
            I => \N__67765\
        );

    \I__16686\ : InMux
    port map (
            O => \N__67776\,
            I => \N__67753\
        );

    \I__16685\ : InMux
    port map (
            O => \N__67775\,
            I => \N__67745\
        );

    \I__16684\ : Span4Mux_v
    port map (
            O => \N__67770\,
            I => \N__67739\
        );

    \I__16683\ : LocalMux
    port map (
            O => \N__67765\,
            I => \N__67739\
        );

    \I__16682\ : InMux
    port map (
            O => \N__67764\,
            I => \N__67734\
        );

    \I__16681\ : InMux
    port map (
            O => \N__67763\,
            I => \N__67734\
        );

    \I__16680\ : InMux
    port map (
            O => \N__67762\,
            I => \N__67724\
        );

    \I__16679\ : InMux
    port map (
            O => \N__67761\,
            I => \N__67724\
        );

    \I__16678\ : InMux
    port map (
            O => \N__67760\,
            I => \N__67724\
        );

    \I__16677\ : InMux
    port map (
            O => \N__67759\,
            I => \N__67721\
        );

    \I__16676\ : InMux
    port map (
            O => \N__67758\,
            I => \N__67718\
        );

    \I__16675\ : InMux
    port map (
            O => \N__67757\,
            I => \N__67715\
        );

    \I__16674\ : InMux
    port map (
            O => \N__67756\,
            I => \N__67712\
        );

    \I__16673\ : LocalMux
    port map (
            O => \N__67753\,
            I => \N__67709\
        );

    \I__16672\ : InMux
    port map (
            O => \N__67752\,
            I => \N__67702\
        );

    \I__16671\ : InMux
    port map (
            O => \N__67751\,
            I => \N__67699\
        );

    \I__16670\ : InMux
    port map (
            O => \N__67750\,
            I => \N__67692\
        );

    \I__16669\ : InMux
    port map (
            O => \N__67749\,
            I => \N__67692\
        );

    \I__16668\ : InMux
    port map (
            O => \N__67748\,
            I => \N__67692\
        );

    \I__16667\ : LocalMux
    port map (
            O => \N__67745\,
            I => \N__67689\
        );

    \I__16666\ : InMux
    port map (
            O => \N__67744\,
            I => \N__67686\
        );

    \I__16665\ : Span4Mux_v
    port map (
            O => \N__67739\,
            I => \N__67682\
        );

    \I__16664\ : LocalMux
    port map (
            O => \N__67734\,
            I => \N__67679\
        );

    \I__16663\ : InMux
    port map (
            O => \N__67733\,
            I => \N__67665\
        );

    \I__16662\ : InMux
    port map (
            O => \N__67732\,
            I => \N__67665\
        );

    \I__16661\ : InMux
    port map (
            O => \N__67731\,
            I => \N__67665\
        );

    \I__16660\ : LocalMux
    port map (
            O => \N__67724\,
            I => \N__67662\
        );

    \I__16659\ : LocalMux
    port map (
            O => \N__67721\,
            I => \N__67659\
        );

    \I__16658\ : LocalMux
    port map (
            O => \N__67718\,
            I => \N__67656\
        );

    \I__16657\ : LocalMux
    port map (
            O => \N__67715\,
            I => \N__67649\
        );

    \I__16656\ : LocalMux
    port map (
            O => \N__67712\,
            I => \N__67649\
        );

    \I__16655\ : Span4Mux_v
    port map (
            O => \N__67709\,
            I => \N__67649\
        );

    \I__16654\ : InMux
    port map (
            O => \N__67708\,
            I => \N__67646\
        );

    \I__16653\ : InMux
    port map (
            O => \N__67707\,
            I => \N__67643\
        );

    \I__16652\ : InMux
    port map (
            O => \N__67706\,
            I => \N__67638\
        );

    \I__16651\ : InMux
    port map (
            O => \N__67705\,
            I => \N__67638\
        );

    \I__16650\ : LocalMux
    port map (
            O => \N__67702\,
            I => \N__67633\
        );

    \I__16649\ : LocalMux
    port map (
            O => \N__67699\,
            I => \N__67633\
        );

    \I__16648\ : LocalMux
    port map (
            O => \N__67692\,
            I => \N__67630\
        );

    \I__16647\ : Span4Mux_v
    port map (
            O => \N__67689\,
            I => \N__67625\
        );

    \I__16646\ : LocalMux
    port map (
            O => \N__67686\,
            I => \N__67625\
        );

    \I__16645\ : InMux
    port map (
            O => \N__67685\,
            I => \N__67617\
        );

    \I__16644\ : Span4Mux_h
    port map (
            O => \N__67682\,
            I => \N__67612\
        );

    \I__16643\ : Span4Mux_v
    port map (
            O => \N__67679\,
            I => \N__67612\
        );

    \I__16642\ : InMux
    port map (
            O => \N__67678\,
            I => \N__67606\
        );

    \I__16641\ : InMux
    port map (
            O => \N__67677\,
            I => \N__67603\
        );

    \I__16640\ : InMux
    port map (
            O => \N__67676\,
            I => \N__67600\
        );

    \I__16639\ : InMux
    port map (
            O => \N__67675\,
            I => \N__67597\
        );

    \I__16638\ : InMux
    port map (
            O => \N__67674\,
            I => \N__67592\
        );

    \I__16637\ : InMux
    port map (
            O => \N__67673\,
            I => \N__67592\
        );

    \I__16636\ : InMux
    port map (
            O => \N__67672\,
            I => \N__67589\
        );

    \I__16635\ : LocalMux
    port map (
            O => \N__67665\,
            I => \N__67586\
        );

    \I__16634\ : Span4Mux_v
    port map (
            O => \N__67662\,
            I => \N__67583\
        );

    \I__16633\ : Span4Mux_v
    port map (
            O => \N__67659\,
            I => \N__67576\
        );

    \I__16632\ : Span4Mux_v
    port map (
            O => \N__67656\,
            I => \N__67576\
        );

    \I__16631\ : Span4Mux_v
    port map (
            O => \N__67649\,
            I => \N__67576\
        );

    \I__16630\ : LocalMux
    port map (
            O => \N__67646\,
            I => \N__67573\
        );

    \I__16629\ : LocalMux
    port map (
            O => \N__67643\,
            I => \N__67564\
        );

    \I__16628\ : LocalMux
    port map (
            O => \N__67638\,
            I => \N__67564\
        );

    \I__16627\ : Span4Mux_v
    port map (
            O => \N__67633\,
            I => \N__67564\
        );

    \I__16626\ : Span4Mux_h
    port map (
            O => \N__67630\,
            I => \N__67564\
        );

    \I__16625\ : Span4Mux_v
    port map (
            O => \N__67625\,
            I => \N__67561\
        );

    \I__16624\ : InMux
    port map (
            O => \N__67624\,
            I => \N__67556\
        );

    \I__16623\ : InMux
    port map (
            O => \N__67623\,
            I => \N__67556\
        );

    \I__16622\ : InMux
    port map (
            O => \N__67622\,
            I => \N__67553\
        );

    \I__16621\ : InMux
    port map (
            O => \N__67621\,
            I => \N__67548\
        );

    \I__16620\ : InMux
    port map (
            O => \N__67620\,
            I => \N__67548\
        );

    \I__16619\ : LocalMux
    port map (
            O => \N__67617\,
            I => \N__67545\
        );

    \I__16618\ : Span4Mux_h
    port map (
            O => \N__67612\,
            I => \N__67542\
        );

    \I__16617\ : InMux
    port map (
            O => \N__67611\,
            I => \N__67539\
        );

    \I__16616\ : InMux
    port map (
            O => \N__67610\,
            I => \N__67536\
        );

    \I__16615\ : InMux
    port map (
            O => \N__67609\,
            I => \N__67533\
        );

    \I__16614\ : LocalMux
    port map (
            O => \N__67606\,
            I => \N__67522\
        );

    \I__16613\ : LocalMux
    port map (
            O => \N__67603\,
            I => \N__67522\
        );

    \I__16612\ : LocalMux
    port map (
            O => \N__67600\,
            I => \N__67522\
        );

    \I__16611\ : LocalMux
    port map (
            O => \N__67597\,
            I => \N__67522\
        );

    \I__16610\ : LocalMux
    port map (
            O => \N__67592\,
            I => \N__67522\
        );

    \I__16609\ : LocalMux
    port map (
            O => \N__67589\,
            I => \N__67513\
        );

    \I__16608\ : Span4Mux_v
    port map (
            O => \N__67586\,
            I => \N__67513\
        );

    \I__16607\ : Span4Mux_v
    port map (
            O => \N__67583\,
            I => \N__67513\
        );

    \I__16606\ : Span4Mux_h
    port map (
            O => \N__67576\,
            I => \N__67513\
        );

    \I__16605\ : Span4Mux_v
    port map (
            O => \N__67573\,
            I => \N__67506\
        );

    \I__16604\ : Span4Mux_v
    port map (
            O => \N__67564\,
            I => \N__67506\
        );

    \I__16603\ : Span4Mux_h
    port map (
            O => \N__67561\,
            I => \N__67506\
        );

    \I__16602\ : LocalMux
    port map (
            O => \N__67556\,
            I => \N__67495\
        );

    \I__16601\ : LocalMux
    port map (
            O => \N__67553\,
            I => \N__67495\
        );

    \I__16600\ : LocalMux
    port map (
            O => \N__67548\,
            I => \N__67495\
        );

    \I__16599\ : Span4Mux_v
    port map (
            O => \N__67545\,
            I => \N__67495\
        );

    \I__16598\ : Span4Mux_h
    port map (
            O => \N__67542\,
            I => \N__67495\
        );

    \I__16597\ : LocalMux
    port map (
            O => \N__67539\,
            I => \c0.n21775\
        );

    \I__16596\ : LocalMux
    port map (
            O => \N__67536\,
            I => \c0.n21775\
        );

    \I__16595\ : LocalMux
    port map (
            O => \N__67533\,
            I => \c0.n21775\
        );

    \I__16594\ : Odrv12
    port map (
            O => \N__67522\,
            I => \c0.n21775\
        );

    \I__16593\ : Odrv4
    port map (
            O => \N__67513\,
            I => \c0.n21775\
        );

    \I__16592\ : Odrv4
    port map (
            O => \N__67506\,
            I => \c0.n21775\
        );

    \I__16591\ : Odrv4
    port map (
            O => \N__67495\,
            I => \c0.n21775\
        );

    \I__16590\ : CascadeMux
    port map (
            O => \N__67480\,
            I => \N__67472\
        );

    \I__16589\ : CascadeMux
    port map (
            O => \N__67479\,
            I => \N__67466\
        );

    \I__16588\ : CascadeMux
    port map (
            O => \N__67478\,
            I => \N__67463\
        );

    \I__16587\ : InMux
    port map (
            O => \N__67477\,
            I => \N__67454\
        );

    \I__16586\ : InMux
    port map (
            O => \N__67476\,
            I => \N__67446\
        );

    \I__16585\ : InMux
    port map (
            O => \N__67475\,
            I => \N__67446\
        );

    \I__16584\ : InMux
    port map (
            O => \N__67472\,
            I => \N__67440\
        );

    \I__16583\ : InMux
    port map (
            O => \N__67471\,
            I => \N__67440\
        );

    \I__16582\ : InMux
    port map (
            O => \N__67470\,
            I => \N__67437\
        );

    \I__16581\ : InMux
    port map (
            O => \N__67469\,
            I => \N__67434\
        );

    \I__16580\ : InMux
    port map (
            O => \N__67466\,
            I => \N__67425\
        );

    \I__16579\ : InMux
    port map (
            O => \N__67463\,
            I => \N__67425\
        );

    \I__16578\ : InMux
    port map (
            O => \N__67462\,
            I => \N__67425\
        );

    \I__16577\ : InMux
    port map (
            O => \N__67461\,
            I => \N__67425\
        );

    \I__16576\ : InMux
    port map (
            O => \N__67460\,
            I => \N__67418\
        );

    \I__16575\ : InMux
    port map (
            O => \N__67459\,
            I => \N__67418\
        );

    \I__16574\ : InMux
    port map (
            O => \N__67458\,
            I => \N__67418\
        );

    \I__16573\ : InMux
    port map (
            O => \N__67457\,
            I => \N__67415\
        );

    \I__16572\ : LocalMux
    port map (
            O => \N__67454\,
            I => \N__67412\
        );

    \I__16571\ : InMux
    port map (
            O => \N__67453\,
            I => \N__67409\
        );

    \I__16570\ : InMux
    port map (
            O => \N__67452\,
            I => \N__67404\
        );

    \I__16569\ : InMux
    port map (
            O => \N__67451\,
            I => \N__67399\
        );

    \I__16568\ : LocalMux
    port map (
            O => \N__67446\,
            I => \N__67396\
        );

    \I__16567\ : InMux
    port map (
            O => \N__67445\,
            I => \N__67393\
        );

    \I__16566\ : LocalMux
    port map (
            O => \N__67440\,
            I => \N__67386\
        );

    \I__16565\ : LocalMux
    port map (
            O => \N__67437\,
            I => \N__67386\
        );

    \I__16564\ : LocalMux
    port map (
            O => \N__67434\,
            I => \N__67383\
        );

    \I__16563\ : LocalMux
    port map (
            O => \N__67425\,
            I => \N__67380\
        );

    \I__16562\ : LocalMux
    port map (
            O => \N__67418\,
            I => \N__67376\
        );

    \I__16561\ : LocalMux
    port map (
            O => \N__67415\,
            I => \N__67373\
        );

    \I__16560\ : Span4Mux_h
    port map (
            O => \N__67412\,
            I => \N__67368\
        );

    \I__16559\ : LocalMux
    port map (
            O => \N__67409\,
            I => \N__67368\
        );

    \I__16558\ : InMux
    port map (
            O => \N__67408\,
            I => \N__67365\
        );

    \I__16557\ : InMux
    port map (
            O => \N__67407\,
            I => \N__67358\
        );

    \I__16556\ : LocalMux
    port map (
            O => \N__67404\,
            I => \N__67355\
        );

    \I__16555\ : InMux
    port map (
            O => \N__67403\,
            I => \N__67352\
        );

    \I__16554\ : CascadeMux
    port map (
            O => \N__67402\,
            I => \N__67349\
        );

    \I__16553\ : LocalMux
    port map (
            O => \N__67399\,
            I => \N__67345\
        );

    \I__16552\ : Span4Mux_h
    port map (
            O => \N__67396\,
            I => \N__67340\
        );

    \I__16551\ : LocalMux
    port map (
            O => \N__67393\,
            I => \N__67340\
        );

    \I__16550\ : InMux
    port map (
            O => \N__67392\,
            I => \N__67334\
        );

    \I__16549\ : InMux
    port map (
            O => \N__67391\,
            I => \N__67334\
        );

    \I__16548\ : Span4Mux_v
    port map (
            O => \N__67386\,
            I => \N__67331\
        );

    \I__16547\ : Span4Mux_v
    port map (
            O => \N__67383\,
            I => \N__67326\
        );

    \I__16546\ : Span4Mux_v
    port map (
            O => \N__67380\,
            I => \N__67326\
        );

    \I__16545\ : InMux
    port map (
            O => \N__67379\,
            I => \N__67323\
        );

    \I__16544\ : Span4Mux_v
    port map (
            O => \N__67376\,
            I => \N__67320\
        );

    \I__16543\ : Span4Mux_v
    port map (
            O => \N__67373\,
            I => \N__67317\
        );

    \I__16542\ : Span4Mux_v
    port map (
            O => \N__67368\,
            I => \N__67312\
        );

    \I__16541\ : LocalMux
    port map (
            O => \N__67365\,
            I => \N__67312\
        );

    \I__16540\ : InMux
    port map (
            O => \N__67364\,
            I => \N__67307\
        );

    \I__16539\ : InMux
    port map (
            O => \N__67363\,
            I => \N__67307\
        );

    \I__16538\ : InMux
    port map (
            O => \N__67362\,
            I => \N__67304\
        );

    \I__16537\ : InMux
    port map (
            O => \N__67361\,
            I => \N__67301\
        );

    \I__16536\ : LocalMux
    port map (
            O => \N__67358\,
            I => \N__67296\
        );

    \I__16535\ : Span4Mux_v
    port map (
            O => \N__67355\,
            I => \N__67296\
        );

    \I__16534\ : LocalMux
    port map (
            O => \N__67352\,
            I => \N__67293\
        );

    \I__16533\ : InMux
    port map (
            O => \N__67349\,
            I => \N__67290\
        );

    \I__16532\ : InMux
    port map (
            O => \N__67348\,
            I => \N__67287\
        );

    \I__16531\ : Sp12to4
    port map (
            O => \N__67345\,
            I => \N__67282\
        );

    \I__16530\ : Sp12to4
    port map (
            O => \N__67340\,
            I => \N__67282\
        );

    \I__16529\ : InMux
    port map (
            O => \N__67339\,
            I => \N__67279\
        );

    \I__16528\ : LocalMux
    port map (
            O => \N__67334\,
            I => \N__67272\
        );

    \I__16527\ : Span4Mux_h
    port map (
            O => \N__67331\,
            I => \N__67272\
        );

    \I__16526\ : Span4Mux_h
    port map (
            O => \N__67326\,
            I => \N__67272\
        );

    \I__16525\ : LocalMux
    port map (
            O => \N__67323\,
            I => \N__67269\
        );

    \I__16524\ : Span4Mux_h
    port map (
            O => \N__67320\,
            I => \N__67262\
        );

    \I__16523\ : Span4Mux_h
    port map (
            O => \N__67317\,
            I => \N__67262\
        );

    \I__16522\ : Span4Mux_v
    port map (
            O => \N__67312\,
            I => \N__67262\
        );

    \I__16521\ : LocalMux
    port map (
            O => \N__67307\,
            I => \N__67251\
        );

    \I__16520\ : LocalMux
    port map (
            O => \N__67304\,
            I => \N__67251\
        );

    \I__16519\ : LocalMux
    port map (
            O => \N__67301\,
            I => \N__67251\
        );

    \I__16518\ : Sp12to4
    port map (
            O => \N__67296\,
            I => \N__67251\
        );

    \I__16517\ : Span12Mux_v
    port map (
            O => \N__67293\,
            I => \N__67251\
        );

    \I__16516\ : LocalMux
    port map (
            O => \N__67290\,
            I => \N__67240\
        );

    \I__16515\ : LocalMux
    port map (
            O => \N__67287\,
            I => \N__67240\
        );

    \I__16514\ : Span12Mux_h
    port map (
            O => \N__67282\,
            I => \N__67240\
        );

    \I__16513\ : LocalMux
    port map (
            O => \N__67279\,
            I => \N__67240\
        );

    \I__16512\ : Sp12to4
    port map (
            O => \N__67272\,
            I => \N__67240\
        );

    \I__16511\ : Span4Mux_h
    port map (
            O => \N__67269\,
            I => \N__67237\
        );

    \I__16510\ : Span4Mux_h
    port map (
            O => \N__67262\,
            I => \N__67234\
        );

    \I__16509\ : Span12Mux_v
    port map (
            O => \N__67251\,
            I => \N__67231\
        );

    \I__16508\ : Span12Mux_v
    port map (
            O => \N__67240\,
            I => \N__67228\
        );

    \I__16507\ : Odrv4
    port map (
            O => \N__67237\,
            I => \c0.n9\
        );

    \I__16506\ : Odrv4
    port map (
            O => \N__67234\,
            I => \c0.n9\
        );

    \I__16505\ : Odrv12
    port map (
            O => \N__67231\,
            I => \c0.n9\
        );

    \I__16504\ : Odrv12
    port map (
            O => \N__67228\,
            I => \c0.n9\
        );

    \I__16503\ : InMux
    port map (
            O => \N__67219\,
            I => \N__67211\
        );

    \I__16502\ : InMux
    port map (
            O => \N__67218\,
            I => \N__67203\
        );

    \I__16501\ : InMux
    port map (
            O => \N__67217\,
            I => \N__67196\
        );

    \I__16500\ : InMux
    port map (
            O => \N__67216\,
            I => \N__67196\
        );

    \I__16499\ : InMux
    port map (
            O => \N__67215\,
            I => \N__67193\
        );

    \I__16498\ : InMux
    port map (
            O => \N__67214\,
            I => \N__67190\
        );

    \I__16497\ : LocalMux
    port map (
            O => \N__67211\,
            I => \N__67187\
        );

    \I__16496\ : CascadeMux
    port map (
            O => \N__67210\,
            I => \N__67183\
        );

    \I__16495\ : CascadeMux
    port map (
            O => \N__67209\,
            I => \N__67180\
        );

    \I__16494\ : CascadeMux
    port map (
            O => \N__67208\,
            I => \N__67177\
        );

    \I__16493\ : InMux
    port map (
            O => \N__67207\,
            I => \N__67172\
        );

    \I__16492\ : InMux
    port map (
            O => \N__67206\,
            I => \N__67172\
        );

    \I__16491\ : LocalMux
    port map (
            O => \N__67203\,
            I => \N__67167\
        );

    \I__16490\ : InMux
    port map (
            O => \N__67202\,
            I => \N__67164\
        );

    \I__16489\ : InMux
    port map (
            O => \N__67201\,
            I => \N__67158\
        );

    \I__16488\ : LocalMux
    port map (
            O => \N__67196\,
            I => \N__67154\
        );

    \I__16487\ : LocalMux
    port map (
            O => \N__67193\,
            I => \N__67149\
        );

    \I__16486\ : LocalMux
    port map (
            O => \N__67190\,
            I => \N__67149\
        );

    \I__16485\ : Span4Mux_v
    port map (
            O => \N__67187\,
            I => \N__67146\
        );

    \I__16484\ : InMux
    port map (
            O => \N__67186\,
            I => \N__67143\
        );

    \I__16483\ : InMux
    port map (
            O => \N__67183\,
            I => \N__67139\
        );

    \I__16482\ : InMux
    port map (
            O => \N__67180\,
            I => \N__67134\
        );

    \I__16481\ : InMux
    port map (
            O => \N__67177\,
            I => \N__67134\
        );

    \I__16480\ : LocalMux
    port map (
            O => \N__67172\,
            I => \N__67131\
        );

    \I__16479\ : InMux
    port map (
            O => \N__67171\,
            I => \N__67128\
        );

    \I__16478\ : InMux
    port map (
            O => \N__67170\,
            I => \N__67125\
        );

    \I__16477\ : Span4Mux_v
    port map (
            O => \N__67167\,
            I => \N__67117\
        );

    \I__16476\ : LocalMux
    port map (
            O => \N__67164\,
            I => \N__67117\
        );

    \I__16475\ : InMux
    port map (
            O => \N__67163\,
            I => \N__67114\
        );

    \I__16474\ : InMux
    port map (
            O => \N__67162\,
            I => \N__67111\
        );

    \I__16473\ : InMux
    port map (
            O => \N__67161\,
            I => \N__67108\
        );

    \I__16472\ : LocalMux
    port map (
            O => \N__67158\,
            I => \N__67105\
        );

    \I__16471\ : InMux
    port map (
            O => \N__67157\,
            I => \N__67100\
        );

    \I__16470\ : Span4Mux_v
    port map (
            O => \N__67154\,
            I => \N__67097\
        );

    \I__16469\ : Span4Mux_v
    port map (
            O => \N__67149\,
            I => \N__67094\
        );

    \I__16468\ : Span4Mux_h
    port map (
            O => \N__67146\,
            I => \N__67089\
        );

    \I__16467\ : LocalMux
    port map (
            O => \N__67143\,
            I => \N__67089\
        );

    \I__16466\ : InMux
    port map (
            O => \N__67142\,
            I => \N__67086\
        );

    \I__16465\ : LocalMux
    port map (
            O => \N__67139\,
            I => \N__67083\
        );

    \I__16464\ : LocalMux
    port map (
            O => \N__67134\,
            I => \N__67080\
        );

    \I__16463\ : Span4Mux_v
    port map (
            O => \N__67131\,
            I => \N__67076\
        );

    \I__16462\ : LocalMux
    port map (
            O => \N__67128\,
            I => \N__67071\
        );

    \I__16461\ : LocalMux
    port map (
            O => \N__67125\,
            I => \N__67071\
        );

    \I__16460\ : InMux
    port map (
            O => \N__67124\,
            I => \N__67067\
        );

    \I__16459\ : InMux
    port map (
            O => \N__67123\,
            I => \N__67064\
        );

    \I__16458\ : InMux
    port map (
            O => \N__67122\,
            I => \N__67060\
        );

    \I__16457\ : Span4Mux_h
    port map (
            O => \N__67117\,
            I => \N__67057\
        );

    \I__16456\ : LocalMux
    port map (
            O => \N__67114\,
            I => \N__67054\
        );

    \I__16455\ : LocalMux
    port map (
            O => \N__67111\,
            I => \N__67051\
        );

    \I__16454\ : LocalMux
    port map (
            O => \N__67108\,
            I => \N__67046\
        );

    \I__16453\ : Span4Mux_h
    port map (
            O => \N__67105\,
            I => \N__67046\
        );

    \I__16452\ : InMux
    port map (
            O => \N__67104\,
            I => \N__67043\
        );

    \I__16451\ : InMux
    port map (
            O => \N__67103\,
            I => \N__67040\
        );

    \I__16450\ : LocalMux
    port map (
            O => \N__67100\,
            I => \N__67033\
        );

    \I__16449\ : Span4Mux_h
    port map (
            O => \N__67097\,
            I => \N__67033\
        );

    \I__16448\ : Span4Mux_h
    port map (
            O => \N__67094\,
            I => \N__67033\
        );

    \I__16447\ : Span4Mux_h
    port map (
            O => \N__67089\,
            I => \N__67030\
        );

    \I__16446\ : LocalMux
    port map (
            O => \N__67086\,
            I => \N__67027\
        );

    \I__16445\ : Span4Mux_v
    port map (
            O => \N__67083\,
            I => \N__67022\
        );

    \I__16444\ : Span4Mux_v
    port map (
            O => \N__67080\,
            I => \N__67022\
        );

    \I__16443\ : InMux
    port map (
            O => \N__67079\,
            I => \N__67019\
        );

    \I__16442\ : Span4Mux_h
    port map (
            O => \N__67076\,
            I => \N__67014\
        );

    \I__16441\ : Span4Mux_v
    port map (
            O => \N__67071\,
            I => \N__67014\
        );

    \I__16440\ : InMux
    port map (
            O => \N__67070\,
            I => \N__67011\
        );

    \I__16439\ : LocalMux
    port map (
            O => \N__67067\,
            I => \N__67006\
        );

    \I__16438\ : LocalMux
    port map (
            O => \N__67064\,
            I => \N__67006\
        );

    \I__16437\ : InMux
    port map (
            O => \N__67063\,
            I => \N__67002\
        );

    \I__16436\ : LocalMux
    port map (
            O => \N__67060\,
            I => \N__66991\
        );

    \I__16435\ : Span4Mux_v
    port map (
            O => \N__67057\,
            I => \N__66991\
        );

    \I__16434\ : Span4Mux_v
    port map (
            O => \N__67054\,
            I => \N__66991\
        );

    \I__16433\ : Span4Mux_v
    port map (
            O => \N__67051\,
            I => \N__66991\
        );

    \I__16432\ : Span4Mux_h
    port map (
            O => \N__67046\,
            I => \N__66991\
        );

    \I__16431\ : LocalMux
    port map (
            O => \N__67043\,
            I => \N__66982\
        );

    \I__16430\ : LocalMux
    port map (
            O => \N__67040\,
            I => \N__66982\
        );

    \I__16429\ : Span4Mux_h
    port map (
            O => \N__67033\,
            I => \N__66982\
        );

    \I__16428\ : Span4Mux_v
    port map (
            O => \N__67030\,
            I => \N__66982\
        );

    \I__16427\ : Sp12to4
    port map (
            O => \N__67027\,
            I => \N__66979\
        );

    \I__16426\ : Sp12to4
    port map (
            O => \N__67022\,
            I => \N__66976\
        );

    \I__16425\ : LocalMux
    port map (
            O => \N__67019\,
            I => \N__66971\
        );

    \I__16424\ : Sp12to4
    port map (
            O => \N__67014\,
            I => \N__66968\
        );

    \I__16423\ : LocalMux
    port map (
            O => \N__67011\,
            I => \N__66963\
        );

    \I__16422\ : Sp12to4
    port map (
            O => \N__67006\,
            I => \N__66963\
        );

    \I__16421\ : InMux
    port map (
            O => \N__67005\,
            I => \N__66960\
        );

    \I__16420\ : LocalMux
    port map (
            O => \N__67002\,
            I => \N__66953\
        );

    \I__16419\ : Span4Mux_h
    port map (
            O => \N__66991\,
            I => \N__66953\
        );

    \I__16418\ : Span4Mux_v
    port map (
            O => \N__66982\,
            I => \N__66953\
        );

    \I__16417\ : Span12Mux_s10_v
    port map (
            O => \N__66979\,
            I => \N__66948\
        );

    \I__16416\ : Span12Mux_h
    port map (
            O => \N__66976\,
            I => \N__66948\
        );

    \I__16415\ : InMux
    port map (
            O => \N__66975\,
            I => \N__66945\
        );

    \I__16414\ : InMux
    port map (
            O => \N__66974\,
            I => \N__66942\
        );

    \I__16413\ : Span4Mux_v
    port map (
            O => \N__66971\,
            I => \N__66939\
        );

    \I__16412\ : Span12Mux_s9_h
    port map (
            O => \N__66968\,
            I => \N__66934\
        );

    \I__16411\ : Span12Mux_v
    port map (
            O => \N__66963\,
            I => \N__66934\
        );

    \I__16410\ : LocalMux
    port map (
            O => \N__66960\,
            I => \N__66929\
        );

    \I__16409\ : Span4Mux_v
    port map (
            O => \N__66953\,
            I => \N__66929\
        );

    \I__16408\ : Span12Mux_v
    port map (
            O => \N__66948\,
            I => \N__66926\
        );

    \I__16407\ : LocalMux
    port map (
            O => \N__66945\,
            I => rx_data_5
        );

    \I__16406\ : LocalMux
    port map (
            O => \N__66942\,
            I => rx_data_5
        );

    \I__16405\ : Odrv4
    port map (
            O => \N__66939\,
            I => rx_data_5
        );

    \I__16404\ : Odrv12
    port map (
            O => \N__66934\,
            I => rx_data_5
        );

    \I__16403\ : Odrv4
    port map (
            O => \N__66929\,
            I => rx_data_5
        );

    \I__16402\ : Odrv12
    port map (
            O => \N__66926\,
            I => rx_data_5
        );

    \I__16401\ : CascadeMux
    port map (
            O => \N__66913\,
            I => \N__66909\
        );

    \I__16400\ : CascadeMux
    port map (
            O => \N__66912\,
            I => \N__66905\
        );

    \I__16399\ : InMux
    port map (
            O => \N__66909\,
            I => \N__66902\
        );

    \I__16398\ : InMux
    port map (
            O => \N__66908\,
            I => \N__66899\
        );

    \I__16397\ : InMux
    port map (
            O => \N__66905\,
            I => \N__66896\
        );

    \I__16396\ : LocalMux
    port map (
            O => \N__66902\,
            I => \N__66893\
        );

    \I__16395\ : LocalMux
    port map (
            O => \N__66899\,
            I => \N__66890\
        );

    \I__16394\ : LocalMux
    port map (
            O => \N__66896\,
            I => \N__66883\
        );

    \I__16393\ : Span4Mux_h
    port map (
            O => \N__66893\,
            I => \N__66883\
        );

    \I__16392\ : Span4Mux_h
    port map (
            O => \N__66890\,
            I => \N__66883\
        );

    \I__16391\ : Odrv4
    port map (
            O => \N__66883\,
            I => \c0.data_in_frame_27_5\
        );

    \I__16390\ : InMux
    port map (
            O => \N__66880\,
            I => \N__66877\
        );

    \I__16389\ : LocalMux
    port map (
            O => \N__66877\,
            I => \N__66872\
        );

    \I__16388\ : ClkMux
    port map (
            O => \N__66876\,
            I => \N__66139\
        );

    \I__16387\ : ClkMux
    port map (
            O => \N__66875\,
            I => \N__66139\
        );

    \I__16386\ : Glb2LocalMux
    port map (
            O => \N__66872\,
            I => \N__66139\
        );

    \I__16385\ : ClkMux
    port map (
            O => \N__66871\,
            I => \N__66139\
        );

    \I__16384\ : ClkMux
    port map (
            O => \N__66870\,
            I => \N__66139\
        );

    \I__16383\ : ClkMux
    port map (
            O => \N__66869\,
            I => \N__66139\
        );

    \I__16382\ : ClkMux
    port map (
            O => \N__66868\,
            I => \N__66139\
        );

    \I__16381\ : ClkMux
    port map (
            O => \N__66867\,
            I => \N__66139\
        );

    \I__16380\ : ClkMux
    port map (
            O => \N__66866\,
            I => \N__66139\
        );

    \I__16379\ : ClkMux
    port map (
            O => \N__66865\,
            I => \N__66139\
        );

    \I__16378\ : ClkMux
    port map (
            O => \N__66864\,
            I => \N__66139\
        );

    \I__16377\ : ClkMux
    port map (
            O => \N__66863\,
            I => \N__66139\
        );

    \I__16376\ : ClkMux
    port map (
            O => \N__66862\,
            I => \N__66139\
        );

    \I__16375\ : ClkMux
    port map (
            O => \N__66861\,
            I => \N__66139\
        );

    \I__16374\ : ClkMux
    port map (
            O => \N__66860\,
            I => \N__66139\
        );

    \I__16373\ : ClkMux
    port map (
            O => \N__66859\,
            I => \N__66139\
        );

    \I__16372\ : ClkMux
    port map (
            O => \N__66858\,
            I => \N__66139\
        );

    \I__16371\ : ClkMux
    port map (
            O => \N__66857\,
            I => \N__66139\
        );

    \I__16370\ : ClkMux
    port map (
            O => \N__66856\,
            I => \N__66139\
        );

    \I__16369\ : ClkMux
    port map (
            O => \N__66855\,
            I => \N__66139\
        );

    \I__16368\ : ClkMux
    port map (
            O => \N__66854\,
            I => \N__66139\
        );

    \I__16367\ : ClkMux
    port map (
            O => \N__66853\,
            I => \N__66139\
        );

    \I__16366\ : ClkMux
    port map (
            O => \N__66852\,
            I => \N__66139\
        );

    \I__16365\ : ClkMux
    port map (
            O => \N__66851\,
            I => \N__66139\
        );

    \I__16364\ : ClkMux
    port map (
            O => \N__66850\,
            I => \N__66139\
        );

    \I__16363\ : ClkMux
    port map (
            O => \N__66849\,
            I => \N__66139\
        );

    \I__16362\ : ClkMux
    port map (
            O => \N__66848\,
            I => \N__66139\
        );

    \I__16361\ : ClkMux
    port map (
            O => \N__66847\,
            I => \N__66139\
        );

    \I__16360\ : ClkMux
    port map (
            O => \N__66846\,
            I => \N__66139\
        );

    \I__16359\ : ClkMux
    port map (
            O => \N__66845\,
            I => \N__66139\
        );

    \I__16358\ : ClkMux
    port map (
            O => \N__66844\,
            I => \N__66139\
        );

    \I__16357\ : ClkMux
    port map (
            O => \N__66843\,
            I => \N__66139\
        );

    \I__16356\ : ClkMux
    port map (
            O => \N__66842\,
            I => \N__66139\
        );

    \I__16355\ : ClkMux
    port map (
            O => \N__66841\,
            I => \N__66139\
        );

    \I__16354\ : ClkMux
    port map (
            O => \N__66840\,
            I => \N__66139\
        );

    \I__16353\ : ClkMux
    port map (
            O => \N__66839\,
            I => \N__66139\
        );

    \I__16352\ : ClkMux
    port map (
            O => \N__66838\,
            I => \N__66139\
        );

    \I__16351\ : ClkMux
    port map (
            O => \N__66837\,
            I => \N__66139\
        );

    \I__16350\ : ClkMux
    port map (
            O => \N__66836\,
            I => \N__66139\
        );

    \I__16349\ : ClkMux
    port map (
            O => \N__66835\,
            I => \N__66139\
        );

    \I__16348\ : ClkMux
    port map (
            O => \N__66834\,
            I => \N__66139\
        );

    \I__16347\ : ClkMux
    port map (
            O => \N__66833\,
            I => \N__66139\
        );

    \I__16346\ : ClkMux
    port map (
            O => \N__66832\,
            I => \N__66139\
        );

    \I__16345\ : ClkMux
    port map (
            O => \N__66831\,
            I => \N__66139\
        );

    \I__16344\ : ClkMux
    port map (
            O => \N__66830\,
            I => \N__66139\
        );

    \I__16343\ : ClkMux
    port map (
            O => \N__66829\,
            I => \N__66139\
        );

    \I__16342\ : ClkMux
    port map (
            O => \N__66828\,
            I => \N__66139\
        );

    \I__16341\ : ClkMux
    port map (
            O => \N__66827\,
            I => \N__66139\
        );

    \I__16340\ : ClkMux
    port map (
            O => \N__66826\,
            I => \N__66139\
        );

    \I__16339\ : ClkMux
    port map (
            O => \N__66825\,
            I => \N__66139\
        );

    \I__16338\ : ClkMux
    port map (
            O => \N__66824\,
            I => \N__66139\
        );

    \I__16337\ : ClkMux
    port map (
            O => \N__66823\,
            I => \N__66139\
        );

    \I__16336\ : ClkMux
    port map (
            O => \N__66822\,
            I => \N__66139\
        );

    \I__16335\ : ClkMux
    port map (
            O => \N__66821\,
            I => \N__66139\
        );

    \I__16334\ : ClkMux
    port map (
            O => \N__66820\,
            I => \N__66139\
        );

    \I__16333\ : ClkMux
    port map (
            O => \N__66819\,
            I => \N__66139\
        );

    \I__16332\ : ClkMux
    port map (
            O => \N__66818\,
            I => \N__66139\
        );

    \I__16331\ : ClkMux
    port map (
            O => \N__66817\,
            I => \N__66139\
        );

    \I__16330\ : ClkMux
    port map (
            O => \N__66816\,
            I => \N__66139\
        );

    \I__16329\ : ClkMux
    port map (
            O => \N__66815\,
            I => \N__66139\
        );

    \I__16328\ : ClkMux
    port map (
            O => \N__66814\,
            I => \N__66139\
        );

    \I__16327\ : ClkMux
    port map (
            O => \N__66813\,
            I => \N__66139\
        );

    \I__16326\ : ClkMux
    port map (
            O => \N__66812\,
            I => \N__66139\
        );

    \I__16325\ : ClkMux
    port map (
            O => \N__66811\,
            I => \N__66139\
        );

    \I__16324\ : ClkMux
    port map (
            O => \N__66810\,
            I => \N__66139\
        );

    \I__16323\ : ClkMux
    port map (
            O => \N__66809\,
            I => \N__66139\
        );

    \I__16322\ : ClkMux
    port map (
            O => \N__66808\,
            I => \N__66139\
        );

    \I__16321\ : ClkMux
    port map (
            O => \N__66807\,
            I => \N__66139\
        );

    \I__16320\ : ClkMux
    port map (
            O => \N__66806\,
            I => \N__66139\
        );

    \I__16319\ : ClkMux
    port map (
            O => \N__66805\,
            I => \N__66139\
        );

    \I__16318\ : ClkMux
    port map (
            O => \N__66804\,
            I => \N__66139\
        );

    \I__16317\ : ClkMux
    port map (
            O => \N__66803\,
            I => \N__66139\
        );

    \I__16316\ : ClkMux
    port map (
            O => \N__66802\,
            I => \N__66139\
        );

    \I__16315\ : ClkMux
    port map (
            O => \N__66801\,
            I => \N__66139\
        );

    \I__16314\ : ClkMux
    port map (
            O => \N__66800\,
            I => \N__66139\
        );

    \I__16313\ : ClkMux
    port map (
            O => \N__66799\,
            I => \N__66139\
        );

    \I__16312\ : ClkMux
    port map (
            O => \N__66798\,
            I => \N__66139\
        );

    \I__16311\ : ClkMux
    port map (
            O => \N__66797\,
            I => \N__66139\
        );

    \I__16310\ : ClkMux
    port map (
            O => \N__66796\,
            I => \N__66139\
        );

    \I__16309\ : ClkMux
    port map (
            O => \N__66795\,
            I => \N__66139\
        );

    \I__16308\ : ClkMux
    port map (
            O => \N__66794\,
            I => \N__66139\
        );

    \I__16307\ : ClkMux
    port map (
            O => \N__66793\,
            I => \N__66139\
        );

    \I__16306\ : ClkMux
    port map (
            O => \N__66792\,
            I => \N__66139\
        );

    \I__16305\ : ClkMux
    port map (
            O => \N__66791\,
            I => \N__66139\
        );

    \I__16304\ : ClkMux
    port map (
            O => \N__66790\,
            I => \N__66139\
        );

    \I__16303\ : ClkMux
    port map (
            O => \N__66789\,
            I => \N__66139\
        );

    \I__16302\ : ClkMux
    port map (
            O => \N__66788\,
            I => \N__66139\
        );

    \I__16301\ : ClkMux
    port map (
            O => \N__66787\,
            I => \N__66139\
        );

    \I__16300\ : ClkMux
    port map (
            O => \N__66786\,
            I => \N__66139\
        );

    \I__16299\ : ClkMux
    port map (
            O => \N__66785\,
            I => \N__66139\
        );

    \I__16298\ : ClkMux
    port map (
            O => \N__66784\,
            I => \N__66139\
        );

    \I__16297\ : ClkMux
    port map (
            O => \N__66783\,
            I => \N__66139\
        );

    \I__16296\ : ClkMux
    port map (
            O => \N__66782\,
            I => \N__66139\
        );

    \I__16295\ : ClkMux
    port map (
            O => \N__66781\,
            I => \N__66139\
        );

    \I__16294\ : ClkMux
    port map (
            O => \N__66780\,
            I => \N__66139\
        );

    \I__16293\ : ClkMux
    port map (
            O => \N__66779\,
            I => \N__66139\
        );

    \I__16292\ : ClkMux
    port map (
            O => \N__66778\,
            I => \N__66139\
        );

    \I__16291\ : ClkMux
    port map (
            O => \N__66777\,
            I => \N__66139\
        );

    \I__16290\ : ClkMux
    port map (
            O => \N__66776\,
            I => \N__66139\
        );

    \I__16289\ : ClkMux
    port map (
            O => \N__66775\,
            I => \N__66139\
        );

    \I__16288\ : ClkMux
    port map (
            O => \N__66774\,
            I => \N__66139\
        );

    \I__16287\ : ClkMux
    port map (
            O => \N__66773\,
            I => \N__66139\
        );

    \I__16286\ : ClkMux
    port map (
            O => \N__66772\,
            I => \N__66139\
        );

    \I__16285\ : ClkMux
    port map (
            O => \N__66771\,
            I => \N__66139\
        );

    \I__16284\ : ClkMux
    port map (
            O => \N__66770\,
            I => \N__66139\
        );

    \I__16283\ : ClkMux
    port map (
            O => \N__66769\,
            I => \N__66139\
        );

    \I__16282\ : ClkMux
    port map (
            O => \N__66768\,
            I => \N__66139\
        );

    \I__16281\ : ClkMux
    port map (
            O => \N__66767\,
            I => \N__66139\
        );

    \I__16280\ : ClkMux
    port map (
            O => \N__66766\,
            I => \N__66139\
        );

    \I__16279\ : ClkMux
    port map (
            O => \N__66765\,
            I => \N__66139\
        );

    \I__16278\ : ClkMux
    port map (
            O => \N__66764\,
            I => \N__66139\
        );

    \I__16277\ : ClkMux
    port map (
            O => \N__66763\,
            I => \N__66139\
        );

    \I__16276\ : ClkMux
    port map (
            O => \N__66762\,
            I => \N__66139\
        );

    \I__16275\ : ClkMux
    port map (
            O => \N__66761\,
            I => \N__66139\
        );

    \I__16274\ : ClkMux
    port map (
            O => \N__66760\,
            I => \N__66139\
        );

    \I__16273\ : ClkMux
    port map (
            O => \N__66759\,
            I => \N__66139\
        );

    \I__16272\ : ClkMux
    port map (
            O => \N__66758\,
            I => \N__66139\
        );

    \I__16271\ : ClkMux
    port map (
            O => \N__66757\,
            I => \N__66139\
        );

    \I__16270\ : ClkMux
    port map (
            O => \N__66756\,
            I => \N__66139\
        );

    \I__16269\ : ClkMux
    port map (
            O => \N__66755\,
            I => \N__66139\
        );

    \I__16268\ : ClkMux
    port map (
            O => \N__66754\,
            I => \N__66139\
        );

    \I__16267\ : ClkMux
    port map (
            O => \N__66753\,
            I => \N__66139\
        );

    \I__16266\ : ClkMux
    port map (
            O => \N__66752\,
            I => \N__66139\
        );

    \I__16265\ : ClkMux
    port map (
            O => \N__66751\,
            I => \N__66139\
        );

    \I__16264\ : ClkMux
    port map (
            O => \N__66750\,
            I => \N__66139\
        );

    \I__16263\ : ClkMux
    port map (
            O => \N__66749\,
            I => \N__66139\
        );

    \I__16262\ : ClkMux
    port map (
            O => \N__66748\,
            I => \N__66139\
        );

    \I__16261\ : ClkMux
    port map (
            O => \N__66747\,
            I => \N__66139\
        );

    \I__16260\ : ClkMux
    port map (
            O => \N__66746\,
            I => \N__66139\
        );

    \I__16259\ : ClkMux
    port map (
            O => \N__66745\,
            I => \N__66139\
        );

    \I__16258\ : ClkMux
    port map (
            O => \N__66744\,
            I => \N__66139\
        );

    \I__16257\ : ClkMux
    port map (
            O => \N__66743\,
            I => \N__66139\
        );

    \I__16256\ : ClkMux
    port map (
            O => \N__66742\,
            I => \N__66139\
        );

    \I__16255\ : ClkMux
    port map (
            O => \N__66741\,
            I => \N__66139\
        );

    \I__16254\ : ClkMux
    port map (
            O => \N__66740\,
            I => \N__66139\
        );

    \I__16253\ : ClkMux
    port map (
            O => \N__66739\,
            I => \N__66139\
        );

    \I__16252\ : ClkMux
    port map (
            O => \N__66738\,
            I => \N__66139\
        );

    \I__16251\ : ClkMux
    port map (
            O => \N__66737\,
            I => \N__66139\
        );

    \I__16250\ : ClkMux
    port map (
            O => \N__66736\,
            I => \N__66139\
        );

    \I__16249\ : ClkMux
    port map (
            O => \N__66735\,
            I => \N__66139\
        );

    \I__16248\ : ClkMux
    port map (
            O => \N__66734\,
            I => \N__66139\
        );

    \I__16247\ : ClkMux
    port map (
            O => \N__66733\,
            I => \N__66139\
        );

    \I__16246\ : ClkMux
    port map (
            O => \N__66732\,
            I => \N__66139\
        );

    \I__16245\ : ClkMux
    port map (
            O => \N__66731\,
            I => \N__66139\
        );

    \I__16244\ : ClkMux
    port map (
            O => \N__66730\,
            I => \N__66139\
        );

    \I__16243\ : ClkMux
    port map (
            O => \N__66729\,
            I => \N__66139\
        );

    \I__16242\ : ClkMux
    port map (
            O => \N__66728\,
            I => \N__66139\
        );

    \I__16241\ : ClkMux
    port map (
            O => \N__66727\,
            I => \N__66139\
        );

    \I__16240\ : ClkMux
    port map (
            O => \N__66726\,
            I => \N__66139\
        );

    \I__16239\ : ClkMux
    port map (
            O => \N__66725\,
            I => \N__66139\
        );

    \I__16238\ : ClkMux
    port map (
            O => \N__66724\,
            I => \N__66139\
        );

    \I__16237\ : ClkMux
    port map (
            O => \N__66723\,
            I => \N__66139\
        );

    \I__16236\ : ClkMux
    port map (
            O => \N__66722\,
            I => \N__66139\
        );

    \I__16235\ : ClkMux
    port map (
            O => \N__66721\,
            I => \N__66139\
        );

    \I__16234\ : ClkMux
    port map (
            O => \N__66720\,
            I => \N__66139\
        );

    \I__16233\ : ClkMux
    port map (
            O => \N__66719\,
            I => \N__66139\
        );

    \I__16232\ : ClkMux
    port map (
            O => \N__66718\,
            I => \N__66139\
        );

    \I__16231\ : ClkMux
    port map (
            O => \N__66717\,
            I => \N__66139\
        );

    \I__16230\ : ClkMux
    port map (
            O => \N__66716\,
            I => \N__66139\
        );

    \I__16229\ : ClkMux
    port map (
            O => \N__66715\,
            I => \N__66139\
        );

    \I__16228\ : ClkMux
    port map (
            O => \N__66714\,
            I => \N__66139\
        );

    \I__16227\ : ClkMux
    port map (
            O => \N__66713\,
            I => \N__66139\
        );

    \I__16226\ : ClkMux
    port map (
            O => \N__66712\,
            I => \N__66139\
        );

    \I__16225\ : ClkMux
    port map (
            O => \N__66711\,
            I => \N__66139\
        );

    \I__16224\ : ClkMux
    port map (
            O => \N__66710\,
            I => \N__66139\
        );

    \I__16223\ : ClkMux
    port map (
            O => \N__66709\,
            I => \N__66139\
        );

    \I__16222\ : ClkMux
    port map (
            O => \N__66708\,
            I => \N__66139\
        );

    \I__16221\ : ClkMux
    port map (
            O => \N__66707\,
            I => \N__66139\
        );

    \I__16220\ : ClkMux
    port map (
            O => \N__66706\,
            I => \N__66139\
        );

    \I__16219\ : ClkMux
    port map (
            O => \N__66705\,
            I => \N__66139\
        );

    \I__16218\ : ClkMux
    port map (
            O => \N__66704\,
            I => \N__66139\
        );

    \I__16217\ : ClkMux
    port map (
            O => \N__66703\,
            I => \N__66139\
        );

    \I__16216\ : ClkMux
    port map (
            O => \N__66702\,
            I => \N__66139\
        );

    \I__16215\ : ClkMux
    port map (
            O => \N__66701\,
            I => \N__66139\
        );

    \I__16214\ : ClkMux
    port map (
            O => \N__66700\,
            I => \N__66139\
        );

    \I__16213\ : ClkMux
    port map (
            O => \N__66699\,
            I => \N__66139\
        );

    \I__16212\ : ClkMux
    port map (
            O => \N__66698\,
            I => \N__66139\
        );

    \I__16211\ : ClkMux
    port map (
            O => \N__66697\,
            I => \N__66139\
        );

    \I__16210\ : ClkMux
    port map (
            O => \N__66696\,
            I => \N__66139\
        );

    \I__16209\ : ClkMux
    port map (
            O => \N__66695\,
            I => \N__66139\
        );

    \I__16208\ : ClkMux
    port map (
            O => \N__66694\,
            I => \N__66139\
        );

    \I__16207\ : ClkMux
    port map (
            O => \N__66693\,
            I => \N__66139\
        );

    \I__16206\ : ClkMux
    port map (
            O => \N__66692\,
            I => \N__66139\
        );

    \I__16205\ : ClkMux
    port map (
            O => \N__66691\,
            I => \N__66139\
        );

    \I__16204\ : ClkMux
    port map (
            O => \N__66690\,
            I => \N__66139\
        );

    \I__16203\ : ClkMux
    port map (
            O => \N__66689\,
            I => \N__66139\
        );

    \I__16202\ : ClkMux
    port map (
            O => \N__66688\,
            I => \N__66139\
        );

    \I__16201\ : ClkMux
    port map (
            O => \N__66687\,
            I => \N__66139\
        );

    \I__16200\ : ClkMux
    port map (
            O => \N__66686\,
            I => \N__66139\
        );

    \I__16199\ : ClkMux
    port map (
            O => \N__66685\,
            I => \N__66139\
        );

    \I__16198\ : ClkMux
    port map (
            O => \N__66684\,
            I => \N__66139\
        );

    \I__16197\ : ClkMux
    port map (
            O => \N__66683\,
            I => \N__66139\
        );

    \I__16196\ : ClkMux
    port map (
            O => \N__66682\,
            I => \N__66139\
        );

    \I__16195\ : ClkMux
    port map (
            O => \N__66681\,
            I => \N__66139\
        );

    \I__16194\ : ClkMux
    port map (
            O => \N__66680\,
            I => \N__66139\
        );

    \I__16193\ : ClkMux
    port map (
            O => \N__66679\,
            I => \N__66139\
        );

    \I__16192\ : ClkMux
    port map (
            O => \N__66678\,
            I => \N__66139\
        );

    \I__16191\ : ClkMux
    port map (
            O => \N__66677\,
            I => \N__66139\
        );

    \I__16190\ : ClkMux
    port map (
            O => \N__66676\,
            I => \N__66139\
        );

    \I__16189\ : ClkMux
    port map (
            O => \N__66675\,
            I => \N__66139\
        );

    \I__16188\ : ClkMux
    port map (
            O => \N__66674\,
            I => \N__66139\
        );

    \I__16187\ : ClkMux
    port map (
            O => \N__66673\,
            I => \N__66139\
        );

    \I__16186\ : ClkMux
    port map (
            O => \N__66672\,
            I => \N__66139\
        );

    \I__16185\ : ClkMux
    port map (
            O => \N__66671\,
            I => \N__66139\
        );

    \I__16184\ : ClkMux
    port map (
            O => \N__66670\,
            I => \N__66139\
        );

    \I__16183\ : ClkMux
    port map (
            O => \N__66669\,
            I => \N__66139\
        );

    \I__16182\ : ClkMux
    port map (
            O => \N__66668\,
            I => \N__66139\
        );

    \I__16181\ : ClkMux
    port map (
            O => \N__66667\,
            I => \N__66139\
        );

    \I__16180\ : ClkMux
    port map (
            O => \N__66666\,
            I => \N__66139\
        );

    \I__16179\ : ClkMux
    port map (
            O => \N__66665\,
            I => \N__66139\
        );

    \I__16178\ : ClkMux
    port map (
            O => \N__66664\,
            I => \N__66139\
        );

    \I__16177\ : ClkMux
    port map (
            O => \N__66663\,
            I => \N__66139\
        );

    \I__16176\ : ClkMux
    port map (
            O => \N__66662\,
            I => \N__66139\
        );

    \I__16175\ : ClkMux
    port map (
            O => \N__66661\,
            I => \N__66139\
        );

    \I__16174\ : ClkMux
    port map (
            O => \N__66660\,
            I => \N__66139\
        );

    \I__16173\ : ClkMux
    port map (
            O => \N__66659\,
            I => \N__66139\
        );

    \I__16172\ : ClkMux
    port map (
            O => \N__66658\,
            I => \N__66139\
        );

    \I__16171\ : ClkMux
    port map (
            O => \N__66657\,
            I => \N__66139\
        );

    \I__16170\ : ClkMux
    port map (
            O => \N__66656\,
            I => \N__66139\
        );

    \I__16169\ : ClkMux
    port map (
            O => \N__66655\,
            I => \N__66139\
        );

    \I__16168\ : ClkMux
    port map (
            O => \N__66654\,
            I => \N__66139\
        );

    \I__16167\ : ClkMux
    port map (
            O => \N__66653\,
            I => \N__66139\
        );

    \I__16166\ : ClkMux
    port map (
            O => \N__66652\,
            I => \N__66139\
        );

    \I__16165\ : ClkMux
    port map (
            O => \N__66651\,
            I => \N__66139\
        );

    \I__16164\ : ClkMux
    port map (
            O => \N__66650\,
            I => \N__66139\
        );

    \I__16163\ : ClkMux
    port map (
            O => \N__66649\,
            I => \N__66139\
        );

    \I__16162\ : ClkMux
    port map (
            O => \N__66648\,
            I => \N__66139\
        );

    \I__16161\ : ClkMux
    port map (
            O => \N__66647\,
            I => \N__66139\
        );

    \I__16160\ : ClkMux
    port map (
            O => \N__66646\,
            I => \N__66139\
        );

    \I__16159\ : ClkMux
    port map (
            O => \N__66645\,
            I => \N__66139\
        );

    \I__16158\ : ClkMux
    port map (
            O => \N__66644\,
            I => \N__66139\
        );

    \I__16157\ : ClkMux
    port map (
            O => \N__66643\,
            I => \N__66139\
        );

    \I__16156\ : ClkMux
    port map (
            O => \N__66642\,
            I => \N__66139\
        );

    \I__16155\ : ClkMux
    port map (
            O => \N__66641\,
            I => \N__66139\
        );

    \I__16154\ : ClkMux
    port map (
            O => \N__66640\,
            I => \N__66139\
        );

    \I__16153\ : ClkMux
    port map (
            O => \N__66639\,
            I => \N__66139\
        );

    \I__16152\ : ClkMux
    port map (
            O => \N__66638\,
            I => \N__66139\
        );

    \I__16151\ : ClkMux
    port map (
            O => \N__66637\,
            I => \N__66139\
        );

    \I__16150\ : ClkMux
    port map (
            O => \N__66636\,
            I => \N__66139\
        );

    \I__16149\ : ClkMux
    port map (
            O => \N__66635\,
            I => \N__66139\
        );

    \I__16148\ : ClkMux
    port map (
            O => \N__66634\,
            I => \N__66139\
        );

    \I__16147\ : ClkMux
    port map (
            O => \N__66633\,
            I => \N__66139\
        );

    \I__16146\ : ClkMux
    port map (
            O => \N__66632\,
            I => \N__66139\
        );

    \I__16145\ : ClkMux
    port map (
            O => \N__66631\,
            I => \N__66139\
        );

    \I__16144\ : ClkMux
    port map (
            O => \N__66630\,
            I => \N__66139\
        );

    \I__16143\ : GlobalMux
    port map (
            O => \N__66139\,
            I => \PIN_9_c\
        );

    \I__16142\ : InMux
    port map (
            O => \N__66136\,
            I => \N__66132\
        );

    \I__16141\ : InMux
    port map (
            O => \N__66135\,
            I => \N__66129\
        );

    \I__16140\ : LocalMux
    port map (
            O => \N__66132\,
            I => \N__66125\
        );

    \I__16139\ : LocalMux
    port map (
            O => \N__66129\,
            I => \N__66121\
        );

    \I__16138\ : InMux
    port map (
            O => \N__66128\,
            I => \N__66118\
        );

    \I__16137\ : Span4Mux_h
    port map (
            O => \N__66125\,
            I => \N__66115\
        );

    \I__16136\ : InMux
    port map (
            O => \N__66124\,
            I => \N__66112\
        );

    \I__16135\ : Span4Mux_h
    port map (
            O => \N__66121\,
            I => \N__66107\
        );

    \I__16134\ : LocalMux
    port map (
            O => \N__66118\,
            I => \N__66107\
        );

    \I__16133\ : Span4Mux_h
    port map (
            O => \N__66115\,
            I => \N__66104\
        );

    \I__16132\ : LocalMux
    port map (
            O => \N__66112\,
            I => \c0.data_in_frame_27_7\
        );

    \I__16131\ : Odrv4
    port map (
            O => \N__66107\,
            I => \c0.data_in_frame_27_7\
        );

    \I__16130\ : Odrv4
    port map (
            O => \N__66104\,
            I => \c0.data_in_frame_27_7\
        );

    \I__16129\ : InMux
    port map (
            O => \N__66097\,
            I => \N__66092\
        );

    \I__16128\ : CascadeMux
    port map (
            O => \N__66096\,
            I => \N__66089\
        );

    \I__16127\ : CascadeMux
    port map (
            O => \N__66095\,
            I => \N__66086\
        );

    \I__16126\ : LocalMux
    port map (
            O => \N__66092\,
            I => \N__66083\
        );

    \I__16125\ : InMux
    port map (
            O => \N__66089\,
            I => \N__66080\
        );

    \I__16124\ : InMux
    port map (
            O => \N__66086\,
            I => \N__66077\
        );

    \I__16123\ : Span4Mux_h
    port map (
            O => \N__66083\,
            I => \N__66072\
        );

    \I__16122\ : LocalMux
    port map (
            O => \N__66080\,
            I => \N__66072\
        );

    \I__16121\ : LocalMux
    port map (
            O => \N__66077\,
            I => \c0.data_in_frame_27_6\
        );

    \I__16120\ : Odrv4
    port map (
            O => \N__66072\,
            I => \c0.data_in_frame_27_6\
        );

    \I__16119\ : InMux
    port map (
            O => \N__66067\,
            I => \N__66060\
        );

    \I__16118\ : InMux
    port map (
            O => \N__66066\,
            I => \N__66060\
        );

    \I__16117\ : InMux
    port map (
            O => \N__66065\,
            I => \N__66057\
        );

    \I__16116\ : LocalMux
    port map (
            O => \N__66060\,
            I => \N__66054\
        );

    \I__16115\ : LocalMux
    port map (
            O => \N__66057\,
            I => \c0.data_in_frame_27_0\
        );

    \I__16114\ : Odrv4
    port map (
            O => \N__66054\,
            I => \c0.data_in_frame_27_0\
        );

    \I__16113\ : InMux
    port map (
            O => \N__66049\,
            I => \N__66045\
        );

    \I__16112\ : InMux
    port map (
            O => \N__66048\,
            I => \N__66042\
        );

    \I__16111\ : LocalMux
    port map (
            O => \N__66045\,
            I => \N__66039\
        );

    \I__16110\ : LocalMux
    port map (
            O => \N__66042\,
            I => \N__66034\
        );

    \I__16109\ : Span4Mux_h
    port map (
            O => \N__66039\,
            I => \N__66034\
        );

    \I__16108\ : Odrv4
    port map (
            O => \N__66034\,
            I => \c0.n6268\
        );

    \I__16107\ : InMux
    port map (
            O => \N__66031\,
            I => \N__66025\
        );

    \I__16106\ : InMux
    port map (
            O => \N__66030\,
            I => \N__66022\
        );

    \I__16105\ : CascadeMux
    port map (
            O => \N__66029\,
            I => \N__66016\
        );

    \I__16104\ : CascadeMux
    port map (
            O => \N__66028\,
            I => \N__66009\
        );

    \I__16103\ : LocalMux
    port map (
            O => \N__66025\,
            I => \N__66004\
        );

    \I__16102\ : LocalMux
    port map (
            O => \N__66022\,
            I => \N__65998\
        );

    \I__16101\ : InMux
    port map (
            O => \N__66021\,
            I => \N__65993\
        );

    \I__16100\ : InMux
    port map (
            O => \N__66020\,
            I => \N__65993\
        );

    \I__16099\ : CascadeMux
    port map (
            O => \N__66019\,
            I => \N__65988\
        );

    \I__16098\ : InMux
    port map (
            O => \N__66016\,
            I => \N__65985\
        );

    \I__16097\ : CascadeMux
    port map (
            O => \N__66015\,
            I => \N__65982\
        );

    \I__16096\ : InMux
    port map (
            O => \N__66014\,
            I => \N__65977\
        );

    \I__16095\ : InMux
    port map (
            O => \N__66013\,
            I => \N__65977\
        );

    \I__16094\ : CascadeMux
    port map (
            O => \N__66012\,
            I => \N__65974\
        );

    \I__16093\ : InMux
    port map (
            O => \N__66009\,
            I => \N__65964\
        );

    \I__16092\ : InMux
    port map (
            O => \N__66008\,
            I => \N__65964\
        );

    \I__16091\ : InMux
    port map (
            O => \N__66007\,
            I => \N__65961\
        );

    \I__16090\ : Span4Mux_v
    port map (
            O => \N__66004\,
            I => \N__65958\
        );

    \I__16089\ : InMux
    port map (
            O => \N__66003\,
            I => \N__65953\
        );

    \I__16088\ : InMux
    port map (
            O => \N__66002\,
            I => \N__65953\
        );

    \I__16087\ : InMux
    port map (
            O => \N__66001\,
            I => \N__65950\
        );

    \I__16086\ : Span4Mux_h
    port map (
            O => \N__65998\,
            I => \N__65944\
        );

    \I__16085\ : LocalMux
    port map (
            O => \N__65993\,
            I => \N__65944\
        );

    \I__16084\ : InMux
    port map (
            O => \N__65992\,
            I => \N__65941\
        );

    \I__16083\ : CascadeMux
    port map (
            O => \N__65991\,
            I => \N__65933\
        );

    \I__16082\ : InMux
    port map (
            O => \N__65988\,
            I => \N__65929\
        );

    \I__16081\ : LocalMux
    port map (
            O => \N__65985\,
            I => \N__65926\
        );

    \I__16080\ : InMux
    port map (
            O => \N__65982\,
            I => \N__65923\
        );

    \I__16079\ : LocalMux
    port map (
            O => \N__65977\,
            I => \N__65920\
        );

    \I__16078\ : InMux
    port map (
            O => \N__65974\,
            I => \N__65917\
        );

    \I__16077\ : InMux
    port map (
            O => \N__65973\,
            I => \N__65908\
        );

    \I__16076\ : InMux
    port map (
            O => \N__65972\,
            I => \N__65908\
        );

    \I__16075\ : InMux
    port map (
            O => \N__65971\,
            I => \N__65908\
        );

    \I__16074\ : InMux
    port map (
            O => \N__65970\,
            I => \N__65908\
        );

    \I__16073\ : InMux
    port map (
            O => \N__65969\,
            I => \N__65905\
        );

    \I__16072\ : LocalMux
    port map (
            O => \N__65964\,
            I => \N__65900\
        );

    \I__16071\ : LocalMux
    port map (
            O => \N__65961\,
            I => \N__65900\
        );

    \I__16070\ : Span4Mux_h
    port map (
            O => \N__65958\,
            I => \N__65894\
        );

    \I__16069\ : LocalMux
    port map (
            O => \N__65953\,
            I => \N__65894\
        );

    \I__16068\ : LocalMux
    port map (
            O => \N__65950\,
            I => \N__65891\
        );

    \I__16067\ : InMux
    port map (
            O => \N__65949\,
            I => \N__65888\
        );

    \I__16066\ : Span4Mux_h
    port map (
            O => \N__65944\,
            I => \N__65885\
        );

    \I__16065\ : LocalMux
    port map (
            O => \N__65941\,
            I => \N__65882\
        );

    \I__16064\ : InMux
    port map (
            O => \N__65940\,
            I => \N__65879\
        );

    \I__16063\ : InMux
    port map (
            O => \N__65939\,
            I => \N__65876\
        );

    \I__16062\ : InMux
    port map (
            O => \N__65938\,
            I => \N__65869\
        );

    \I__16061\ : InMux
    port map (
            O => \N__65937\,
            I => \N__65869\
        );

    \I__16060\ : InMux
    port map (
            O => \N__65936\,
            I => \N__65869\
        );

    \I__16059\ : InMux
    port map (
            O => \N__65933\,
            I => \N__65866\
        );

    \I__16058\ : InMux
    port map (
            O => \N__65932\,
            I => \N__65862\
        );

    \I__16057\ : LocalMux
    port map (
            O => \N__65929\,
            I => \N__65859\
        );

    \I__16056\ : Span4Mux_h
    port map (
            O => \N__65926\,
            I => \N__65850\
        );

    \I__16055\ : LocalMux
    port map (
            O => \N__65923\,
            I => \N__65850\
        );

    \I__16054\ : Span4Mux_v
    port map (
            O => \N__65920\,
            I => \N__65850\
        );

    \I__16053\ : LocalMux
    port map (
            O => \N__65917\,
            I => \N__65850\
        );

    \I__16052\ : LocalMux
    port map (
            O => \N__65908\,
            I => \N__65847\
        );

    \I__16051\ : LocalMux
    port map (
            O => \N__65905\,
            I => \N__65842\
        );

    \I__16050\ : Span4Mux_h
    port map (
            O => \N__65900\,
            I => \N__65842\
        );

    \I__16049\ : InMux
    port map (
            O => \N__65899\,
            I => \N__65839\
        );

    \I__16048\ : Span4Mux_v
    port map (
            O => \N__65894\,
            I => \N__65834\
        );

    \I__16047\ : Span4Mux_v
    port map (
            O => \N__65891\,
            I => \N__65834\
        );

    \I__16046\ : LocalMux
    port map (
            O => \N__65888\,
            I => \N__65825\
        );

    \I__16045\ : Span4Mux_v
    port map (
            O => \N__65885\,
            I => \N__65825\
        );

    \I__16044\ : Span4Mux_h
    port map (
            O => \N__65882\,
            I => \N__65825\
        );

    \I__16043\ : LocalMux
    port map (
            O => \N__65879\,
            I => \N__65825\
        );

    \I__16042\ : LocalMux
    port map (
            O => \N__65876\,
            I => \N__65822\
        );

    \I__16041\ : LocalMux
    port map (
            O => \N__65869\,
            I => \N__65819\
        );

    \I__16040\ : LocalMux
    port map (
            O => \N__65866\,
            I => \N__65816\
        );

    \I__16039\ : InMux
    port map (
            O => \N__65865\,
            I => \N__65813\
        );

    \I__16038\ : LocalMux
    port map (
            O => \N__65862\,
            I => \N__65806\
        );

    \I__16037\ : Span4Mux_h
    port map (
            O => \N__65859\,
            I => \N__65806\
        );

    \I__16036\ : Span4Mux_v
    port map (
            O => \N__65850\,
            I => \N__65806\
        );

    \I__16035\ : Span4Mux_h
    port map (
            O => \N__65847\,
            I => \N__65801\
        );

    \I__16034\ : Span4Mux_v
    port map (
            O => \N__65842\,
            I => \N__65801\
        );

    \I__16033\ : LocalMux
    port map (
            O => \N__65839\,
            I => \N__65798\
        );

    \I__16032\ : Span4Mux_h
    port map (
            O => \N__65834\,
            I => \N__65793\
        );

    \I__16031\ : Span4Mux_v
    port map (
            O => \N__65825\,
            I => \N__65793\
        );

    \I__16030\ : Span4Mux_v
    port map (
            O => \N__65822\,
            I => \N__65788\
        );

    \I__16029\ : Span4Mux_v
    port map (
            O => \N__65819\,
            I => \N__65788\
        );

    \I__16028\ : Span12Mux_v
    port map (
            O => \N__65816\,
            I => \N__65785\
        );

    \I__16027\ : LocalMux
    port map (
            O => \N__65813\,
            I => \N__65780\
        );

    \I__16026\ : Sp12to4
    port map (
            O => \N__65806\,
            I => \N__65780\
        );

    \I__16025\ : Span4Mux_v
    port map (
            O => \N__65801\,
            I => \N__65777\
        );

    \I__16024\ : Span4Mux_v
    port map (
            O => \N__65798\,
            I => \N__65772\
        );

    \I__16023\ : Span4Mux_h
    port map (
            O => \N__65793\,
            I => \N__65772\
        );

    \I__16022\ : Odrv4
    port map (
            O => \N__65788\,
            I => \c0.n9_adj_4278\
        );

    \I__16021\ : Odrv12
    port map (
            O => \N__65785\,
            I => \c0.n9_adj_4278\
        );

    \I__16020\ : Odrv12
    port map (
            O => \N__65780\,
            I => \c0.n9_adj_4278\
        );

    \I__16019\ : Odrv4
    port map (
            O => \N__65777\,
            I => \c0.n9_adj_4278\
        );

    \I__16018\ : Odrv4
    port map (
            O => \N__65772\,
            I => \c0.n9_adj_4278\
        );

    \I__16017\ : InMux
    port map (
            O => \N__65761\,
            I => \N__65756\
        );

    \I__16016\ : InMux
    port map (
            O => \N__65760\,
            I => \N__65751\
        );

    \I__16015\ : InMux
    port map (
            O => \N__65759\,
            I => \N__65751\
        );

    \I__16014\ : LocalMux
    port map (
            O => \N__65756\,
            I => \N__65747\
        );

    \I__16013\ : LocalMux
    port map (
            O => \N__65751\,
            I => \N__65744\
        );

    \I__16012\ : CascadeMux
    port map (
            O => \N__65750\,
            I => \N__65741\
        );

    \I__16011\ : Span4Mux_h
    port map (
            O => \N__65747\,
            I => \N__65738\
        );

    \I__16010\ : Span4Mux_h
    port map (
            O => \N__65744\,
            I => \N__65735\
        );

    \I__16009\ : InMux
    port map (
            O => \N__65741\,
            I => \N__65732\
        );

    \I__16008\ : Span4Mux_v
    port map (
            O => \N__65738\,
            I => \N__65729\
        );

    \I__16007\ : Span4Mux_v
    port map (
            O => \N__65735\,
            I => \N__65726\
        );

    \I__16006\ : LocalMux
    port map (
            O => \N__65732\,
            I => \c0.data_in_frame_16_7\
        );

    \I__16005\ : Odrv4
    port map (
            O => \N__65729\,
            I => \c0.data_in_frame_16_7\
        );

    \I__16004\ : Odrv4
    port map (
            O => \N__65726\,
            I => \c0.data_in_frame_16_7\
        );

    \I__16003\ : InMux
    port map (
            O => \N__65719\,
            I => \N__65715\
        );

    \I__16002\ : CascadeMux
    port map (
            O => \N__65718\,
            I => \N__65712\
        );

    \I__16001\ : LocalMux
    port map (
            O => \N__65715\,
            I => \N__65709\
        );

    \I__16000\ : InMux
    port map (
            O => \N__65712\,
            I => \N__65706\
        );

    \I__15999\ : Span4Mux_h
    port map (
            O => \N__65709\,
            I => \N__65703\
        );

    \I__15998\ : LocalMux
    port map (
            O => \N__65706\,
            I => \c0.data_in_frame_19_0\
        );

    \I__15997\ : Odrv4
    port map (
            O => \N__65703\,
            I => \c0.data_in_frame_19_0\
        );

    \I__15996\ : InMux
    port map (
            O => \N__65698\,
            I => \N__65693\
        );

    \I__15995\ : InMux
    port map (
            O => \N__65697\,
            I => \N__65690\
        );

    \I__15994\ : CascadeMux
    port map (
            O => \N__65696\,
            I => \N__65686\
        );

    \I__15993\ : LocalMux
    port map (
            O => \N__65693\,
            I => \N__65681\
        );

    \I__15992\ : LocalMux
    port map (
            O => \N__65690\,
            I => \N__65681\
        );

    \I__15991\ : InMux
    port map (
            O => \N__65689\,
            I => \N__65678\
        );

    \I__15990\ : InMux
    port map (
            O => \N__65686\,
            I => \N__65675\
        );

    \I__15989\ : Span4Mux_v
    port map (
            O => \N__65681\,
            I => \N__65667\
        );

    \I__15988\ : LocalMux
    port map (
            O => \N__65678\,
            I => \N__65662\
        );

    \I__15987\ : LocalMux
    port map (
            O => \N__65675\,
            I => \N__65662\
        );

    \I__15986\ : InMux
    port map (
            O => \N__65674\,
            I => \N__65658\
        );

    \I__15985\ : InMux
    port map (
            O => \N__65673\,
            I => \N__65655\
        );

    \I__15984\ : InMux
    port map (
            O => \N__65672\,
            I => \N__65650\
        );

    \I__15983\ : InMux
    port map (
            O => \N__65671\,
            I => \N__65650\
        );

    \I__15982\ : InMux
    port map (
            O => \N__65670\,
            I => \N__65644\
        );

    \I__15981\ : Span4Mux_h
    port map (
            O => \N__65667\,
            I => \N__65639\
        );

    \I__15980\ : Span4Mux_v
    port map (
            O => \N__65662\,
            I => \N__65639\
        );

    \I__15979\ : InMux
    port map (
            O => \N__65661\,
            I => \N__65636\
        );

    \I__15978\ : LocalMux
    port map (
            O => \N__65658\,
            I => \N__65631\
        );

    \I__15977\ : LocalMux
    port map (
            O => \N__65655\,
            I => \N__65631\
        );

    \I__15976\ : LocalMux
    port map (
            O => \N__65650\,
            I => \N__65628\
        );

    \I__15975\ : InMux
    port map (
            O => \N__65649\,
            I => \N__65625\
        );

    \I__15974\ : InMux
    port map (
            O => \N__65648\,
            I => \N__65620\
        );

    \I__15973\ : CascadeMux
    port map (
            O => \N__65647\,
            I => \N__65617\
        );

    \I__15972\ : LocalMux
    port map (
            O => \N__65644\,
            I => \N__65604\
        );

    \I__15971\ : Span4Mux_h
    port map (
            O => \N__65639\,
            I => \N__65604\
        );

    \I__15970\ : LocalMux
    port map (
            O => \N__65636\,
            I => \N__65604\
        );

    \I__15969\ : Span4Mux_v
    port map (
            O => \N__65631\,
            I => \N__65604\
        );

    \I__15968\ : Span4Mux_h
    port map (
            O => \N__65628\,
            I => \N__65604\
        );

    \I__15967\ : LocalMux
    port map (
            O => \N__65625\,
            I => \N__65604\
        );

    \I__15966\ : InMux
    port map (
            O => \N__65624\,
            I => \N__65601\
        );

    \I__15965\ : InMux
    port map (
            O => \N__65623\,
            I => \N__65598\
        );

    \I__15964\ : LocalMux
    port map (
            O => \N__65620\,
            I => \N__65595\
        );

    \I__15963\ : InMux
    port map (
            O => \N__65617\,
            I => \N__65592\
        );

    \I__15962\ : Span4Mux_h
    port map (
            O => \N__65604\,
            I => \N__65588\
        );

    \I__15961\ : LocalMux
    port map (
            O => \N__65601\,
            I => \N__65583\
        );

    \I__15960\ : LocalMux
    port map (
            O => \N__65598\,
            I => \N__65583\
        );

    \I__15959\ : Span4Mux_v
    port map (
            O => \N__65595\,
            I => \N__65577\
        );

    \I__15958\ : LocalMux
    port map (
            O => \N__65592\,
            I => \N__65577\
        );

    \I__15957\ : CascadeMux
    port map (
            O => \N__65591\,
            I => \N__65564\
        );

    \I__15956\ : Span4Mux_v
    port map (
            O => \N__65588\,
            I => \N__65557\
        );

    \I__15955\ : Span4Mux_v
    port map (
            O => \N__65583\,
            I => \N__65557\
        );

    \I__15954\ : InMux
    port map (
            O => \N__65582\,
            I => \N__65554\
        );

    \I__15953\ : Span4Mux_h
    port map (
            O => \N__65577\,
            I => \N__65551\
        );

    \I__15952\ : InMux
    port map (
            O => \N__65576\,
            I => \N__65548\
        );

    \I__15951\ : InMux
    port map (
            O => \N__65575\,
            I => \N__65545\
        );

    \I__15950\ : InMux
    port map (
            O => \N__65574\,
            I => \N__65542\
        );

    \I__15949\ : InMux
    port map (
            O => \N__65573\,
            I => \N__65537\
        );

    \I__15948\ : InMux
    port map (
            O => \N__65572\,
            I => \N__65537\
        );

    \I__15947\ : InMux
    port map (
            O => \N__65571\,
            I => \N__65532\
        );

    \I__15946\ : InMux
    port map (
            O => \N__65570\,
            I => \N__65532\
        );

    \I__15945\ : InMux
    port map (
            O => \N__65569\,
            I => \N__65529\
        );

    \I__15944\ : InMux
    port map (
            O => \N__65568\,
            I => \N__65524\
        );

    \I__15943\ : InMux
    port map (
            O => \N__65567\,
            I => \N__65524\
        );

    \I__15942\ : InMux
    port map (
            O => \N__65564\,
            I => \N__65521\
        );

    \I__15941\ : InMux
    port map (
            O => \N__65563\,
            I => \N__65518\
        );

    \I__15940\ : InMux
    port map (
            O => \N__65562\,
            I => \N__65515\
        );

    \I__15939\ : Sp12to4
    port map (
            O => \N__65557\,
            I => \N__65512\
        );

    \I__15938\ : LocalMux
    port map (
            O => \N__65554\,
            I => \N__65509\
        );

    \I__15937\ : Sp12to4
    port map (
            O => \N__65551\,
            I => \N__65504\
        );

    \I__15936\ : LocalMux
    port map (
            O => \N__65548\,
            I => \N__65504\
        );

    \I__15935\ : LocalMux
    port map (
            O => \N__65545\,
            I => \N__65498\
        );

    \I__15934\ : LocalMux
    port map (
            O => \N__65542\,
            I => \N__65495\
        );

    \I__15933\ : LocalMux
    port map (
            O => \N__65537\,
            I => \N__65492\
        );

    \I__15932\ : LocalMux
    port map (
            O => \N__65532\,
            I => \N__65489\
        );

    \I__15931\ : LocalMux
    port map (
            O => \N__65529\,
            I => \N__65486\
        );

    \I__15930\ : LocalMux
    port map (
            O => \N__65524\,
            I => \N__65481\
        );

    \I__15929\ : LocalMux
    port map (
            O => \N__65521\,
            I => \N__65481\
        );

    \I__15928\ : LocalMux
    port map (
            O => \N__65518\,
            I => \N__65470\
        );

    \I__15927\ : LocalMux
    port map (
            O => \N__65515\,
            I => \N__65470\
        );

    \I__15926\ : Span12Mux_h
    port map (
            O => \N__65512\,
            I => \N__65470\
        );

    \I__15925\ : Span12Mux_h
    port map (
            O => \N__65509\,
            I => \N__65470\
        );

    \I__15924\ : Span12Mux_s9_v
    port map (
            O => \N__65504\,
            I => \N__65470\
        );

    \I__15923\ : InMux
    port map (
            O => \N__65503\,
            I => \N__65465\
        );

    \I__15922\ : InMux
    port map (
            O => \N__65502\,
            I => \N__65465\
        );

    \I__15921\ : InMux
    port map (
            O => \N__65501\,
            I => \N__65462\
        );

    \I__15920\ : Span4Mux_h
    port map (
            O => \N__65498\,
            I => \N__65459\
        );

    \I__15919\ : Span4Mux_v
    port map (
            O => \N__65495\,
            I => \N__65454\
        );

    \I__15918\ : Span4Mux_v
    port map (
            O => \N__65492\,
            I => \N__65454\
        );

    \I__15917\ : Span12Mux_v
    port map (
            O => \N__65489\,
            I => \N__65451\
        );

    \I__15916\ : Span12Mux_v
    port map (
            O => \N__65486\,
            I => \N__65446\
        );

    \I__15915\ : Span12Mux_h
    port map (
            O => \N__65481\,
            I => \N__65446\
        );

    \I__15914\ : Span12Mux_v
    port map (
            O => \N__65470\,
            I => \N__65443\
        );

    \I__15913\ : LocalMux
    port map (
            O => \N__65465\,
            I => rx_data_6
        );

    \I__15912\ : LocalMux
    port map (
            O => \N__65462\,
            I => rx_data_6
        );

    \I__15911\ : Odrv4
    port map (
            O => \N__65459\,
            I => rx_data_6
        );

    \I__15910\ : Odrv4
    port map (
            O => \N__65454\,
            I => rx_data_6
        );

    \I__15909\ : Odrv12
    port map (
            O => \N__65451\,
            I => rx_data_6
        );

    \I__15908\ : Odrv12
    port map (
            O => \N__65446\,
            I => rx_data_6
        );

    \I__15907\ : Odrv12
    port map (
            O => \N__65443\,
            I => rx_data_6
        );

    \I__15906\ : InMux
    port map (
            O => \N__65428\,
            I => \N__65425\
        );

    \I__15905\ : LocalMux
    port map (
            O => \N__65425\,
            I => \N__65421\
        );

    \I__15904\ : CascadeMux
    port map (
            O => \N__65424\,
            I => \N__65418\
        );

    \I__15903\ : Span4Mux_h
    port map (
            O => \N__65421\,
            I => \N__65414\
        );

    \I__15902\ : InMux
    port map (
            O => \N__65418\,
            I => \N__65409\
        );

    \I__15901\ : InMux
    port map (
            O => \N__65417\,
            I => \N__65409\
        );

    \I__15900\ : Odrv4
    port map (
            O => \N__65414\,
            I => \c0.data_in_frame_18_6\
        );

    \I__15899\ : LocalMux
    port map (
            O => \N__65409\,
            I => \c0.data_in_frame_18_6\
        );

    \I__15898\ : CascadeMux
    port map (
            O => \N__65404\,
            I => \N__65401\
        );

    \I__15897\ : InMux
    port map (
            O => \N__65401\,
            I => \N__65397\
        );

    \I__15896\ : CascadeMux
    port map (
            O => \N__65400\,
            I => \N__65394\
        );

    \I__15895\ : LocalMux
    port map (
            O => \N__65397\,
            I => \N__65391\
        );

    \I__15894\ : InMux
    port map (
            O => \N__65394\,
            I => \N__65388\
        );

    \I__15893\ : Span4Mux_h
    port map (
            O => \N__65391\,
            I => \N__65385\
        );

    \I__15892\ : LocalMux
    port map (
            O => \N__65388\,
            I => \N__65380\
        );

    \I__15891\ : Span4Mux_v
    port map (
            O => \N__65385\,
            I => \N__65380\
        );

    \I__15890\ : Span4Mux_v
    port map (
            O => \N__65380\,
            I => \N__65375\
        );

    \I__15889\ : InMux
    port map (
            O => \N__65379\,
            I => \N__65370\
        );

    \I__15888\ : InMux
    port map (
            O => \N__65378\,
            I => \N__65370\
        );

    \I__15887\ : Odrv4
    port map (
            O => \N__65375\,
            I => \c0.data_in_frame_18_7\
        );

    \I__15886\ : LocalMux
    port map (
            O => \N__65370\,
            I => \c0.data_in_frame_18_7\
        );

    \I__15885\ : InMux
    port map (
            O => \N__65365\,
            I => \N__65361\
        );

    \I__15884\ : InMux
    port map (
            O => \N__65364\,
            I => \N__65358\
        );

    \I__15883\ : LocalMux
    port map (
            O => \N__65361\,
            I => \N__65352\
        );

    \I__15882\ : LocalMux
    port map (
            O => \N__65358\,
            I => \N__65349\
        );

    \I__15881\ : InMux
    port map (
            O => \N__65357\,
            I => \N__65344\
        );

    \I__15880\ : InMux
    port map (
            O => \N__65356\,
            I => \N__65344\
        );

    \I__15879\ : InMux
    port map (
            O => \N__65355\,
            I => \N__65341\
        );

    \I__15878\ : Span4Mux_v
    port map (
            O => \N__65352\,
            I => \N__65338\
        );

    \I__15877\ : Span4Mux_h
    port map (
            O => \N__65349\,
            I => \N__65335\
        );

    \I__15876\ : LocalMux
    port map (
            O => \N__65344\,
            I => \c0.data_in_frame_21_5\
        );

    \I__15875\ : LocalMux
    port map (
            O => \N__65341\,
            I => \c0.data_in_frame_21_5\
        );

    \I__15874\ : Odrv4
    port map (
            O => \N__65338\,
            I => \c0.data_in_frame_21_5\
        );

    \I__15873\ : Odrv4
    port map (
            O => \N__65335\,
            I => \c0.data_in_frame_21_5\
        );

    \I__15872\ : InMux
    port map (
            O => \N__65326\,
            I => \N__65323\
        );

    \I__15871\ : LocalMux
    port map (
            O => \N__65323\,
            I => \N__65319\
        );

    \I__15870\ : InMux
    port map (
            O => \N__65322\,
            I => \N__65316\
        );

    \I__15869\ : Span4Mux_h
    port map (
            O => \N__65319\,
            I => \N__65311\
        );

    \I__15868\ : LocalMux
    port map (
            O => \N__65316\,
            I => \N__65311\
        );

    \I__15867\ : Span4Mux_h
    port map (
            O => \N__65311\,
            I => \N__65308\
        );

    \I__15866\ : Odrv4
    port map (
            O => \N__65308\,
            I => \c0.n22123\
        );

    \I__15865\ : InMux
    port map (
            O => \N__65305\,
            I => \N__65301\
        );

    \I__15864\ : InMux
    port map (
            O => \N__65304\,
            I => \N__65298\
        );

    \I__15863\ : LocalMux
    port map (
            O => \N__65301\,
            I => \N__65292\
        );

    \I__15862\ : LocalMux
    port map (
            O => \N__65298\,
            I => \N__65292\
        );

    \I__15861\ : CascadeMux
    port map (
            O => \N__65297\,
            I => \N__65289\
        );

    \I__15860\ : Span4Mux_v
    port map (
            O => \N__65292\,
            I => \N__65286\
        );

    \I__15859\ : InMux
    port map (
            O => \N__65289\,
            I => \N__65283\
        );

    \I__15858\ : Span4Mux_v
    port map (
            O => \N__65286\,
            I => \N__65280\
        );

    \I__15857\ : LocalMux
    port map (
            O => \N__65283\,
            I => \c0.data_in_frame_23_7\
        );

    \I__15856\ : Odrv4
    port map (
            O => \N__65280\,
            I => \c0.data_in_frame_23_7\
        );

    \I__15855\ : CascadeMux
    port map (
            O => \N__65275\,
            I => \N__65272\
        );

    \I__15854\ : InMux
    port map (
            O => \N__65272\,
            I => \N__65269\
        );

    \I__15853\ : LocalMux
    port map (
            O => \N__65269\,
            I => \N__65266\
        );

    \I__15852\ : Span4Mux_h
    port map (
            O => \N__65266\,
            I => \N__65262\
        );

    \I__15851\ : InMux
    port map (
            O => \N__65265\,
            I => \N__65259\
        );

    \I__15850\ : Sp12to4
    port map (
            O => \N__65262\,
            I => \N__65256\
        );

    \I__15849\ : LocalMux
    port map (
            O => \N__65259\,
            I => \N__65253\
        );

    \I__15848\ : Odrv12
    port map (
            O => \N__65256\,
            I => \c0.n22396\
        );

    \I__15847\ : Odrv12
    port map (
            O => \N__65253\,
            I => \c0.n22396\
        );

    \I__15846\ : InMux
    port map (
            O => \N__65248\,
            I => \N__65242\
        );

    \I__15845\ : InMux
    port map (
            O => \N__65247\,
            I => \N__65239\
        );

    \I__15844\ : InMux
    port map (
            O => \N__65246\,
            I => \N__65234\
        );

    \I__15843\ : InMux
    port map (
            O => \N__65245\,
            I => \N__65234\
        );

    \I__15842\ : LocalMux
    port map (
            O => \N__65242\,
            I => \N__65231\
        );

    \I__15841\ : LocalMux
    port map (
            O => \N__65239\,
            I => \N__65227\
        );

    \I__15840\ : LocalMux
    port map (
            O => \N__65234\,
            I => \N__65224\
        );

    \I__15839\ : Span4Mux_h
    port map (
            O => \N__65231\,
            I => \N__65221\
        );

    \I__15838\ : InMux
    port map (
            O => \N__65230\,
            I => \N__65218\
        );

    \I__15837\ : Span4Mux_v
    port map (
            O => \N__65227\,
            I => \N__65213\
        );

    \I__15836\ : Span4Mux_h
    port map (
            O => \N__65224\,
            I => \N__65213\
        );

    \I__15835\ : Odrv4
    port map (
            O => \N__65221\,
            I => \c0.n20288\
        );

    \I__15834\ : LocalMux
    port map (
            O => \N__65218\,
            I => \c0.n20288\
        );

    \I__15833\ : Odrv4
    port map (
            O => \N__65213\,
            I => \c0.n20288\
        );

    \I__15832\ : InMux
    port map (
            O => \N__65206\,
            I => \N__65203\
        );

    \I__15831\ : LocalMux
    port map (
            O => \N__65203\,
            I => \c0.n23\
        );

    \I__15830\ : InMux
    port map (
            O => \N__65200\,
            I => \N__65197\
        );

    \I__15829\ : LocalMux
    port map (
            O => \N__65197\,
            I => \N__65194\
        );

    \I__15828\ : Span4Mux_v
    port map (
            O => \N__65194\,
            I => \N__65189\
        );

    \I__15827\ : InMux
    port map (
            O => \N__65193\,
            I => \N__65186\
        );

    \I__15826\ : CascadeMux
    port map (
            O => \N__65192\,
            I => \N__65183\
        );

    \I__15825\ : Span4Mux_v
    port map (
            O => \N__65189\,
            I => \N__65180\
        );

    \I__15824\ : LocalMux
    port map (
            O => \N__65186\,
            I => \N__65176\
        );

    \I__15823\ : InMux
    port map (
            O => \N__65183\,
            I => \N__65173\
        );

    \I__15822\ : Span4Mux_h
    port map (
            O => \N__65180\,
            I => \N__65170\
        );

    \I__15821\ : InMux
    port map (
            O => \N__65179\,
            I => \N__65167\
        );

    \I__15820\ : Span4Mux_v
    port map (
            O => \N__65176\,
            I => \N__65164\
        );

    \I__15819\ : LocalMux
    port map (
            O => \N__65173\,
            I => \c0.data_in_frame_24_2\
        );

    \I__15818\ : Odrv4
    port map (
            O => \N__65170\,
            I => \c0.data_in_frame_24_2\
        );

    \I__15817\ : LocalMux
    port map (
            O => \N__65167\,
            I => \c0.data_in_frame_24_2\
        );

    \I__15816\ : Odrv4
    port map (
            O => \N__65164\,
            I => \c0.data_in_frame_24_2\
        );

    \I__15815\ : InMux
    port map (
            O => \N__65155\,
            I => \N__65150\
        );

    \I__15814\ : InMux
    port map (
            O => \N__65154\,
            I => \N__65147\
        );

    \I__15813\ : InMux
    port map (
            O => \N__65153\,
            I => \N__65143\
        );

    \I__15812\ : LocalMux
    port map (
            O => \N__65150\,
            I => \N__65140\
        );

    \I__15811\ : LocalMux
    port map (
            O => \N__65147\,
            I => \N__65137\
        );

    \I__15810\ : InMux
    port map (
            O => \N__65146\,
            I => \N__65134\
        );

    \I__15809\ : LocalMux
    port map (
            O => \N__65143\,
            I => \N__65131\
        );

    \I__15808\ : Span4Mux_h
    port map (
            O => \N__65140\,
            I => \N__65128\
        );

    \I__15807\ : Span4Mux_v
    port map (
            O => \N__65137\,
            I => \N__65123\
        );

    \I__15806\ : LocalMux
    port map (
            O => \N__65134\,
            I => \N__65123\
        );

    \I__15805\ : Span4Mux_v
    port map (
            O => \N__65131\,
            I => \N__65120\
        );

    \I__15804\ : Odrv4
    port map (
            O => \N__65128\,
            I => \c0.n13443\
        );

    \I__15803\ : Odrv4
    port map (
            O => \N__65123\,
            I => \c0.n13443\
        );

    \I__15802\ : Odrv4
    port map (
            O => \N__65120\,
            I => \c0.n13443\
        );

    \I__15801\ : CascadeMux
    port map (
            O => \N__65113\,
            I => \N__65110\
        );

    \I__15800\ : InMux
    port map (
            O => \N__65110\,
            I => \N__65107\
        );

    \I__15799\ : LocalMux
    port map (
            O => \N__65107\,
            I => \N__65104\
        );

    \I__15798\ : Span4Mux_v
    port map (
            O => \N__65104\,
            I => \N__65100\
        );

    \I__15797\ : CascadeMux
    port map (
            O => \N__65103\,
            I => \N__65097\
        );

    \I__15796\ : Span4Mux_h
    port map (
            O => \N__65100\,
            I => \N__65094\
        );

    \I__15795\ : InMux
    port map (
            O => \N__65097\,
            I => \N__65091\
        );

    \I__15794\ : Sp12to4
    port map (
            O => \N__65094\,
            I => \N__65086\
        );

    \I__15793\ : LocalMux
    port map (
            O => \N__65091\,
            I => \N__65086\
        );

    \I__15792\ : Span12Mux_v
    port map (
            O => \N__65086\,
            I => \N__65083\
        );

    \I__15791\ : Odrv12
    port map (
            O => \N__65083\,
            I => \c0.n22358\
        );

    \I__15790\ : InMux
    port map (
            O => \N__65080\,
            I => \N__65077\
        );

    \I__15789\ : LocalMux
    port map (
            O => \N__65077\,
            I => \N__65074\
        );

    \I__15788\ : Span4Mux_v
    port map (
            O => \N__65074\,
            I => \N__65070\
        );

    \I__15787\ : InMux
    port map (
            O => \N__65073\,
            I => \N__65067\
        );

    \I__15786\ : Odrv4
    port map (
            O => \N__65070\,
            I => \c0.n22099\
        );

    \I__15785\ : LocalMux
    port map (
            O => \N__65067\,
            I => \c0.n22099\
        );

    \I__15784\ : InMux
    port map (
            O => \N__65062\,
            I => \N__65054\
        );

    \I__15783\ : InMux
    port map (
            O => \N__65061\,
            I => \N__65054\
        );

    \I__15782\ : CascadeMux
    port map (
            O => \N__65060\,
            I => \N__65050\
        );

    \I__15781\ : InMux
    port map (
            O => \N__65059\,
            I => \N__65047\
        );

    \I__15780\ : LocalMux
    port map (
            O => \N__65054\,
            I => \N__65044\
        );

    \I__15779\ : CascadeMux
    port map (
            O => \N__65053\,
            I => \N__65041\
        );

    \I__15778\ : InMux
    port map (
            O => \N__65050\,
            I => \N__65038\
        );

    \I__15777\ : LocalMux
    port map (
            O => \N__65047\,
            I => \N__65035\
        );

    \I__15776\ : Span4Mux_h
    port map (
            O => \N__65044\,
            I => \N__65032\
        );

    \I__15775\ : InMux
    port map (
            O => \N__65041\,
            I => \N__65029\
        );

    \I__15774\ : LocalMux
    port map (
            O => \N__65038\,
            I => \c0.data_in_frame_24_1\
        );

    \I__15773\ : Odrv12
    port map (
            O => \N__65035\,
            I => \c0.data_in_frame_24_1\
        );

    \I__15772\ : Odrv4
    port map (
            O => \N__65032\,
            I => \c0.data_in_frame_24_1\
        );

    \I__15771\ : LocalMux
    port map (
            O => \N__65029\,
            I => \c0.data_in_frame_24_1\
        );

    \I__15770\ : InMux
    port map (
            O => \N__65020\,
            I => \N__65017\
        );

    \I__15769\ : LocalMux
    port map (
            O => \N__65017\,
            I => \N__65013\
        );

    \I__15768\ : InMux
    port map (
            O => \N__65016\,
            I => \N__65010\
        );

    \I__15767\ : Span4Mux_h
    port map (
            O => \N__65013\,
            I => \N__65007\
        );

    \I__15766\ : LocalMux
    port map (
            O => \N__65010\,
            I => \N__65004\
        );

    \I__15765\ : Span4Mux_h
    port map (
            O => \N__65007\,
            I => \N__65001\
        );

    \I__15764\ : Span12Mux_v
    port map (
            O => \N__65004\,
            I => \N__64998\
        );

    \I__15763\ : Span4Mux_v
    port map (
            O => \N__65001\,
            I => \N__64995\
        );

    \I__15762\ : Odrv12
    port map (
            O => \N__64998\,
            I => \c0.n22057\
        );

    \I__15761\ : Odrv4
    port map (
            O => \N__64995\,
            I => \c0.n22057\
        );

    \I__15760\ : InMux
    port map (
            O => \N__64990\,
            I => \N__64986\
        );

    \I__15759\ : InMux
    port map (
            O => \N__64989\,
            I => \N__64983\
        );

    \I__15758\ : LocalMux
    port map (
            O => \N__64986\,
            I => \N__64980\
        );

    \I__15757\ : LocalMux
    port map (
            O => \N__64983\,
            I => \c0.n22373\
        );

    \I__15756\ : Odrv12
    port map (
            O => \N__64980\,
            I => \c0.n22373\
        );

    \I__15755\ : CascadeMux
    port map (
            O => \N__64975\,
            I => \c0.n8_adj_4288_cascade_\
        );

    \I__15754\ : InMux
    port map (
            O => \N__64972\,
            I => \N__64969\
        );

    \I__15753\ : LocalMux
    port map (
            O => \N__64969\,
            I => \N__64966\
        );

    \I__15752\ : Odrv12
    port map (
            O => \N__64966\,
            I => \c0.n24_adj_4289\
        );

    \I__15751\ : InMux
    port map (
            O => \N__64963\,
            I => \N__64957\
        );

    \I__15750\ : InMux
    port map (
            O => \N__64962\,
            I => \N__64957\
        );

    \I__15749\ : LocalMux
    port map (
            O => \N__64957\,
            I => \N__64954\
        );

    \I__15748\ : Odrv4
    port map (
            O => \N__64954\,
            I => \c0.n22215\
        );

    \I__15747\ : InMux
    port map (
            O => \N__64951\,
            I => \N__64948\
        );

    \I__15746\ : LocalMux
    port map (
            O => \N__64948\,
            I => \N__64944\
        );

    \I__15745\ : InMux
    port map (
            O => \N__64947\,
            I => \N__64941\
        );

    \I__15744\ : Span4Mux_v
    port map (
            O => \N__64944\,
            I => \N__64938\
        );

    \I__15743\ : LocalMux
    port map (
            O => \N__64941\,
            I => \c0.n22402\
        );

    \I__15742\ : Odrv4
    port map (
            O => \N__64938\,
            I => \c0.n22402\
        );

    \I__15741\ : CascadeMux
    port map (
            O => \N__64933\,
            I => \N__64929\
        );

    \I__15740\ : CascadeMux
    port map (
            O => \N__64932\,
            I => \N__64926\
        );

    \I__15739\ : InMux
    port map (
            O => \N__64929\,
            I => \N__64923\
        );

    \I__15738\ : InMux
    port map (
            O => \N__64926\,
            I => \N__64920\
        );

    \I__15737\ : LocalMux
    port map (
            O => \N__64923\,
            I => \N__64917\
        );

    \I__15736\ : LocalMux
    port map (
            O => \N__64920\,
            I => \c0.data_in_frame_28_4\
        );

    \I__15735\ : Odrv12
    port map (
            O => \N__64917\,
            I => \c0.data_in_frame_28_4\
        );

    \I__15734\ : InMux
    port map (
            O => \N__64912\,
            I => \N__64908\
        );

    \I__15733\ : InMux
    port map (
            O => \N__64911\,
            I => \N__64905\
        );

    \I__15732\ : LocalMux
    port map (
            O => \N__64908\,
            I => \c0.n22455\
        );

    \I__15731\ : LocalMux
    port map (
            O => \N__64905\,
            I => \c0.n22455\
        );

    \I__15730\ : InMux
    port map (
            O => \N__64900\,
            I => \N__64897\
        );

    \I__15729\ : LocalMux
    port map (
            O => \N__64897\,
            I => \c0.n22997\
        );

    \I__15728\ : InMux
    port map (
            O => \N__64894\,
            I => \N__64889\
        );

    \I__15727\ : CascadeMux
    port map (
            O => \N__64893\,
            I => \N__64880\
        );

    \I__15726\ : CascadeMux
    port map (
            O => \N__64892\,
            I => \N__64876\
        );

    \I__15725\ : LocalMux
    port map (
            O => \N__64889\,
            I => \N__64868\
        );

    \I__15724\ : InMux
    port map (
            O => \N__64888\,
            I => \N__64865\
        );

    \I__15723\ : InMux
    port map (
            O => \N__64887\,
            I => \N__64859\
        );

    \I__15722\ : InMux
    port map (
            O => \N__64886\,
            I => \N__64854\
        );

    \I__15721\ : InMux
    port map (
            O => \N__64885\,
            I => \N__64854\
        );

    \I__15720\ : InMux
    port map (
            O => \N__64884\,
            I => \N__64846\
        );

    \I__15719\ : InMux
    port map (
            O => \N__64883\,
            I => \N__64846\
        );

    \I__15718\ : InMux
    port map (
            O => \N__64880\,
            I => \N__64843\
        );

    \I__15717\ : InMux
    port map (
            O => \N__64879\,
            I => \N__64840\
        );

    \I__15716\ : InMux
    port map (
            O => \N__64876\,
            I => \N__64837\
        );

    \I__15715\ : InMux
    port map (
            O => \N__64875\,
            I => \N__64833\
        );

    \I__15714\ : InMux
    port map (
            O => \N__64874\,
            I => \N__64830\
        );

    \I__15713\ : InMux
    port map (
            O => \N__64873\,
            I => \N__64827\
        );

    \I__15712\ : InMux
    port map (
            O => \N__64872\,
            I => \N__64820\
        );

    \I__15711\ : InMux
    port map (
            O => \N__64871\,
            I => \N__64815\
        );

    \I__15710\ : Span4Mux_v
    port map (
            O => \N__64868\,
            I => \N__64812\
        );

    \I__15709\ : LocalMux
    port map (
            O => \N__64865\,
            I => \N__64809\
        );

    \I__15708\ : InMux
    port map (
            O => \N__64864\,
            I => \N__64806\
        );

    \I__15707\ : InMux
    port map (
            O => \N__64863\,
            I => \N__64803\
        );

    \I__15706\ : InMux
    port map (
            O => \N__64862\,
            I => \N__64800\
        );

    \I__15705\ : LocalMux
    port map (
            O => \N__64859\,
            I => \N__64797\
        );

    \I__15704\ : LocalMux
    port map (
            O => \N__64854\,
            I => \N__64794\
        );

    \I__15703\ : InMux
    port map (
            O => \N__64853\,
            I => \N__64789\
        );

    \I__15702\ : InMux
    port map (
            O => \N__64852\,
            I => \N__64789\
        );

    \I__15701\ : InMux
    port map (
            O => \N__64851\,
            I => \N__64786\
        );

    \I__15700\ : LocalMux
    port map (
            O => \N__64846\,
            I => \N__64781\
        );

    \I__15699\ : LocalMux
    port map (
            O => \N__64843\,
            I => \N__64781\
        );

    \I__15698\ : LocalMux
    port map (
            O => \N__64840\,
            I => \N__64778\
        );

    \I__15697\ : LocalMux
    port map (
            O => \N__64837\,
            I => \N__64775\
        );

    \I__15696\ : InMux
    port map (
            O => \N__64836\,
            I => \N__64772\
        );

    \I__15695\ : LocalMux
    port map (
            O => \N__64833\,
            I => \N__64767\
        );

    \I__15694\ : LocalMux
    port map (
            O => \N__64830\,
            I => \N__64767\
        );

    \I__15693\ : LocalMux
    port map (
            O => \N__64827\,
            I => \N__64764\
        );

    \I__15692\ : InMux
    port map (
            O => \N__64826\,
            I => \N__64761\
        );

    \I__15691\ : InMux
    port map (
            O => \N__64825\,
            I => \N__64758\
        );

    \I__15690\ : InMux
    port map (
            O => \N__64824\,
            I => \N__64755\
        );

    \I__15689\ : InMux
    port map (
            O => \N__64823\,
            I => \N__64752\
        );

    \I__15688\ : LocalMux
    port map (
            O => \N__64820\,
            I => \N__64749\
        );

    \I__15687\ : CascadeMux
    port map (
            O => \N__64819\,
            I => \N__64745\
        );

    \I__15686\ : InMux
    port map (
            O => \N__64818\,
            I => \N__64742\
        );

    \I__15685\ : LocalMux
    port map (
            O => \N__64815\,
            I => \N__64739\
        );

    \I__15684\ : Span4Mux_h
    port map (
            O => \N__64812\,
            I => \N__64734\
        );

    \I__15683\ : Span4Mux_v
    port map (
            O => \N__64809\,
            I => \N__64734\
        );

    \I__15682\ : LocalMux
    port map (
            O => \N__64806\,
            I => \N__64731\
        );

    \I__15681\ : LocalMux
    port map (
            O => \N__64803\,
            I => \N__64726\
        );

    \I__15680\ : LocalMux
    port map (
            O => \N__64800\,
            I => \N__64726\
        );

    \I__15679\ : Span4Mux_h
    port map (
            O => \N__64797\,
            I => \N__64721\
        );

    \I__15678\ : Span4Mux_v
    port map (
            O => \N__64794\,
            I => \N__64721\
        );

    \I__15677\ : LocalMux
    port map (
            O => \N__64789\,
            I => \N__64718\
        );

    \I__15676\ : LocalMux
    port map (
            O => \N__64786\,
            I => \N__64715\
        );

    \I__15675\ : Span4Mux_h
    port map (
            O => \N__64781\,
            I => \N__64706\
        );

    \I__15674\ : Span4Mux_v
    port map (
            O => \N__64778\,
            I => \N__64706\
        );

    \I__15673\ : Span4Mux_h
    port map (
            O => \N__64775\,
            I => \N__64706\
        );

    \I__15672\ : LocalMux
    port map (
            O => \N__64772\,
            I => \N__64706\
        );

    \I__15671\ : Span4Mux_v
    port map (
            O => \N__64767\,
            I => \N__64701\
        );

    \I__15670\ : Span4Mux_h
    port map (
            O => \N__64764\,
            I => \N__64701\
        );

    \I__15669\ : LocalMux
    port map (
            O => \N__64761\,
            I => \N__64695\
        );

    \I__15668\ : LocalMux
    port map (
            O => \N__64758\,
            I => \N__64692\
        );

    \I__15667\ : LocalMux
    port map (
            O => \N__64755\,
            I => \N__64689\
        );

    \I__15666\ : LocalMux
    port map (
            O => \N__64752\,
            I => \N__64686\
        );

    \I__15665\ : Span4Mux_h
    port map (
            O => \N__64749\,
            I => \N__64683\
        );

    \I__15664\ : InMux
    port map (
            O => \N__64748\,
            I => \N__64678\
        );

    \I__15663\ : InMux
    port map (
            O => \N__64745\,
            I => \N__64678\
        );

    \I__15662\ : LocalMux
    port map (
            O => \N__64742\,
            I => \N__64671\
        );

    \I__15661\ : Span4Mux_v
    port map (
            O => \N__64739\,
            I => \N__64671\
        );

    \I__15660\ : Span4Mux_v
    port map (
            O => \N__64734\,
            I => \N__64671\
        );

    \I__15659\ : Span4Mux_v
    port map (
            O => \N__64731\,
            I => \N__64668\
        );

    \I__15658\ : Span4Mux_v
    port map (
            O => \N__64726\,
            I => \N__64665\
        );

    \I__15657\ : Span4Mux_v
    port map (
            O => \N__64721\,
            I => \N__64660\
        );

    \I__15656\ : Span4Mux_h
    port map (
            O => \N__64718\,
            I => \N__64660\
        );

    \I__15655\ : Span4Mux_h
    port map (
            O => \N__64715\,
            I => \N__64653\
        );

    \I__15654\ : Span4Mux_v
    port map (
            O => \N__64706\,
            I => \N__64653\
        );

    \I__15653\ : Span4Mux_h
    port map (
            O => \N__64701\,
            I => \N__64653\
        );

    \I__15652\ : InMux
    port map (
            O => \N__64700\,
            I => \N__64650\
        );

    \I__15651\ : InMux
    port map (
            O => \N__64699\,
            I => \N__64645\
        );

    \I__15650\ : InMux
    port map (
            O => \N__64698\,
            I => \N__64645\
        );

    \I__15649\ : Span4Mux_h
    port map (
            O => \N__64695\,
            I => \N__64642\
        );

    \I__15648\ : Span4Mux_h
    port map (
            O => \N__64692\,
            I => \N__64633\
        );

    \I__15647\ : Span4Mux_v
    port map (
            O => \N__64689\,
            I => \N__64633\
        );

    \I__15646\ : Span4Mux_v
    port map (
            O => \N__64686\,
            I => \N__64633\
        );

    \I__15645\ : Span4Mux_h
    port map (
            O => \N__64683\,
            I => \N__64633\
        );

    \I__15644\ : LocalMux
    port map (
            O => \N__64678\,
            I => \N__64626\
        );

    \I__15643\ : Sp12to4
    port map (
            O => \N__64671\,
            I => \N__64626\
        );

    \I__15642\ : Sp12to4
    port map (
            O => \N__64668\,
            I => \N__64626\
        );

    \I__15641\ : Span4Mux_h
    port map (
            O => \N__64665\,
            I => \N__64621\
        );

    \I__15640\ : Span4Mux_h
    port map (
            O => \N__64660\,
            I => \N__64621\
        );

    \I__15639\ : Span4Mux_v
    port map (
            O => \N__64653\,
            I => \N__64618\
        );

    \I__15638\ : LocalMux
    port map (
            O => \N__64650\,
            I => rx_data_3
        );

    \I__15637\ : LocalMux
    port map (
            O => \N__64645\,
            I => rx_data_3
        );

    \I__15636\ : Odrv4
    port map (
            O => \N__64642\,
            I => rx_data_3
        );

    \I__15635\ : Odrv4
    port map (
            O => \N__64633\,
            I => rx_data_3
        );

    \I__15634\ : Odrv12
    port map (
            O => \N__64626\,
            I => rx_data_3
        );

    \I__15633\ : Odrv4
    port map (
            O => \N__64621\,
            I => rx_data_3
        );

    \I__15632\ : Odrv4
    port map (
            O => \N__64618\,
            I => rx_data_3
        );

    \I__15631\ : CascadeMux
    port map (
            O => \N__64603\,
            I => \N__64600\
        );

    \I__15630\ : InMux
    port map (
            O => \N__64600\,
            I => \N__64596\
        );

    \I__15629\ : InMux
    port map (
            O => \N__64599\,
            I => \N__64593\
        );

    \I__15628\ : LocalMux
    port map (
            O => \N__64596\,
            I => \c0.data_in_frame_28_3\
        );

    \I__15627\ : LocalMux
    port map (
            O => \N__64593\,
            I => \c0.data_in_frame_28_3\
        );

    \I__15626\ : InMux
    port map (
            O => \N__64588\,
            I => \N__64584\
        );

    \I__15625\ : CascadeMux
    port map (
            O => \N__64587\,
            I => \N__64581\
        );

    \I__15624\ : LocalMux
    port map (
            O => \N__64584\,
            I => \N__64578\
        );

    \I__15623\ : InMux
    port map (
            O => \N__64581\,
            I => \N__64575\
        );

    \I__15622\ : Span4Mux_h
    port map (
            O => \N__64578\,
            I => \N__64572\
        );

    \I__15621\ : LocalMux
    port map (
            O => \N__64575\,
            I => \c0.data_in_frame_28_7\
        );

    \I__15620\ : Odrv4
    port map (
            O => \N__64572\,
            I => \c0.data_in_frame_28_7\
        );

    \I__15619\ : CascadeMux
    port map (
            O => \N__64567\,
            I => \N__64562\
        );

    \I__15618\ : InMux
    port map (
            O => \N__64566\,
            I => \N__64557\
        );

    \I__15617\ : InMux
    port map (
            O => \N__64565\,
            I => \N__64553\
        );

    \I__15616\ : InMux
    port map (
            O => \N__64562\,
            I => \N__64546\
        );

    \I__15615\ : InMux
    port map (
            O => \N__64561\,
            I => \N__64543\
        );

    \I__15614\ : InMux
    port map (
            O => \N__64560\,
            I => \N__64540\
        );

    \I__15613\ : LocalMux
    port map (
            O => \N__64557\,
            I => \N__64537\
        );

    \I__15612\ : CascadeMux
    port map (
            O => \N__64556\,
            I => \N__64528\
        );

    \I__15611\ : LocalMux
    port map (
            O => \N__64553\,
            I => \N__64524\
        );

    \I__15610\ : CascadeMux
    port map (
            O => \N__64552\,
            I => \N__64520\
        );

    \I__15609\ : CascadeMux
    port map (
            O => \N__64551\,
            I => \N__64514\
        );

    \I__15608\ : InMux
    port map (
            O => \N__64550\,
            I => \N__64508\
        );

    \I__15607\ : InMux
    port map (
            O => \N__64549\,
            I => \N__64505\
        );

    \I__15606\ : LocalMux
    port map (
            O => \N__64546\,
            I => \N__64502\
        );

    \I__15605\ : LocalMux
    port map (
            O => \N__64543\,
            I => \N__64499\
        );

    \I__15604\ : LocalMux
    port map (
            O => \N__64540\,
            I => \N__64495\
        );

    \I__15603\ : Span4Mux_v
    port map (
            O => \N__64537\,
            I => \N__64492\
        );

    \I__15602\ : InMux
    port map (
            O => \N__64536\,
            I => \N__64487\
        );

    \I__15601\ : InMux
    port map (
            O => \N__64535\,
            I => \N__64487\
        );

    \I__15600\ : InMux
    port map (
            O => \N__64534\,
            I => \N__64482\
        );

    \I__15599\ : InMux
    port map (
            O => \N__64533\,
            I => \N__64482\
        );

    \I__15598\ : InMux
    port map (
            O => \N__64532\,
            I => \N__64478\
        );

    \I__15597\ : InMux
    port map (
            O => \N__64531\,
            I => \N__64473\
        );

    \I__15596\ : InMux
    port map (
            O => \N__64528\,
            I => \N__64473\
        );

    \I__15595\ : InMux
    port map (
            O => \N__64527\,
            I => \N__64470\
        );

    \I__15594\ : Span4Mux_h
    port map (
            O => \N__64524\,
            I => \N__64467\
        );

    \I__15593\ : InMux
    port map (
            O => \N__64523\,
            I => \N__64464\
        );

    \I__15592\ : InMux
    port map (
            O => \N__64520\,
            I => \N__64459\
        );

    \I__15591\ : InMux
    port map (
            O => \N__64519\,
            I => \N__64459\
        );

    \I__15590\ : InMux
    port map (
            O => \N__64518\,
            I => \N__64455\
        );

    \I__15589\ : InMux
    port map (
            O => \N__64517\,
            I => \N__64452\
        );

    \I__15588\ : InMux
    port map (
            O => \N__64514\,
            I => \N__64448\
        );

    \I__15587\ : InMux
    port map (
            O => \N__64513\,
            I => \N__64441\
        );

    \I__15586\ : InMux
    port map (
            O => \N__64512\,
            I => \N__64441\
        );

    \I__15585\ : InMux
    port map (
            O => \N__64511\,
            I => \N__64441\
        );

    \I__15584\ : LocalMux
    port map (
            O => \N__64508\,
            I => \N__64438\
        );

    \I__15583\ : LocalMux
    port map (
            O => \N__64505\,
            I => \N__64435\
        );

    \I__15582\ : Span4Mux_v
    port map (
            O => \N__64502\,
            I => \N__64430\
        );

    \I__15581\ : Span4Mux_h
    port map (
            O => \N__64499\,
            I => \N__64430\
        );

    \I__15580\ : InMux
    port map (
            O => \N__64498\,
            I => \N__64427\
        );

    \I__15579\ : Span4Mux_h
    port map (
            O => \N__64495\,
            I => \N__64420\
        );

    \I__15578\ : Span4Mux_h
    port map (
            O => \N__64492\,
            I => \N__64420\
        );

    \I__15577\ : LocalMux
    port map (
            O => \N__64487\,
            I => \N__64420\
        );

    \I__15576\ : LocalMux
    port map (
            O => \N__64482\,
            I => \N__64417\
        );

    \I__15575\ : InMux
    port map (
            O => \N__64481\,
            I => \N__64414\
        );

    \I__15574\ : LocalMux
    port map (
            O => \N__64478\,
            I => \N__64411\
        );

    \I__15573\ : LocalMux
    port map (
            O => \N__64473\,
            I => \N__64404\
        );

    \I__15572\ : LocalMux
    port map (
            O => \N__64470\,
            I => \N__64404\
        );

    \I__15571\ : Span4Mux_v
    port map (
            O => \N__64467\,
            I => \N__64404\
        );

    \I__15570\ : LocalMux
    port map (
            O => \N__64464\,
            I => \N__64399\
        );

    \I__15569\ : LocalMux
    port map (
            O => \N__64459\,
            I => \N__64399\
        );

    \I__15568\ : CascadeMux
    port map (
            O => \N__64458\,
            I => \N__64396\
        );

    \I__15567\ : LocalMux
    port map (
            O => \N__64455\,
            I => \N__64391\
        );

    \I__15566\ : LocalMux
    port map (
            O => \N__64452\,
            I => \N__64391\
        );

    \I__15565\ : InMux
    port map (
            O => \N__64451\,
            I => \N__64388\
        );

    \I__15564\ : LocalMux
    port map (
            O => \N__64448\,
            I => \N__64385\
        );

    \I__15563\ : LocalMux
    port map (
            O => \N__64441\,
            I => \N__64382\
        );

    \I__15562\ : Span4Mux_h
    port map (
            O => \N__64438\,
            I => \N__64375\
        );

    \I__15561\ : Span4Mux_h
    port map (
            O => \N__64435\,
            I => \N__64375\
        );

    \I__15560\ : Span4Mux_v
    port map (
            O => \N__64430\,
            I => \N__64375\
        );

    \I__15559\ : LocalMux
    port map (
            O => \N__64427\,
            I => \N__64372\
        );

    \I__15558\ : Span4Mux_v
    port map (
            O => \N__64420\,
            I => \N__64365\
        );

    \I__15557\ : Span4Mux_h
    port map (
            O => \N__64417\,
            I => \N__64365\
        );

    \I__15556\ : LocalMux
    port map (
            O => \N__64414\,
            I => \N__64365\
        );

    \I__15555\ : Span4Mux_h
    port map (
            O => \N__64411\,
            I => \N__64358\
        );

    \I__15554\ : Span4Mux_v
    port map (
            O => \N__64404\,
            I => \N__64358\
        );

    \I__15553\ : Span4Mux_h
    port map (
            O => \N__64399\,
            I => \N__64358\
        );

    \I__15552\ : InMux
    port map (
            O => \N__64396\,
            I => \N__64353\
        );

    \I__15551\ : Span4Mux_h
    port map (
            O => \N__64391\,
            I => \N__64350\
        );

    \I__15550\ : LocalMux
    port map (
            O => \N__64388\,
            I => \N__64347\
        );

    \I__15549\ : Span4Mux_v
    port map (
            O => \N__64385\,
            I => \N__64342\
        );

    \I__15548\ : Span12Mux_h
    port map (
            O => \N__64382\,
            I => \N__64339\
        );

    \I__15547\ : Span4Mux_v
    port map (
            O => \N__64375\,
            I => \N__64336\
        );

    \I__15546\ : Span4Mux_v
    port map (
            O => \N__64372\,
            I => \N__64333\
        );

    \I__15545\ : Span4Mux_v
    port map (
            O => \N__64365\,
            I => \N__64328\
        );

    \I__15544\ : Span4Mux_v
    port map (
            O => \N__64358\,
            I => \N__64328\
        );

    \I__15543\ : InMux
    port map (
            O => \N__64357\,
            I => \N__64323\
        );

    \I__15542\ : InMux
    port map (
            O => \N__64356\,
            I => \N__64323\
        );

    \I__15541\ : LocalMux
    port map (
            O => \N__64353\,
            I => \N__64316\
        );

    \I__15540\ : Span4Mux_h
    port map (
            O => \N__64350\,
            I => \N__64316\
        );

    \I__15539\ : Span4Mux_h
    port map (
            O => \N__64347\,
            I => \N__64316\
        );

    \I__15538\ : InMux
    port map (
            O => \N__64346\,
            I => \N__64313\
        );

    \I__15537\ : InMux
    port map (
            O => \N__64345\,
            I => \N__64310\
        );

    \I__15536\ : Sp12to4
    port map (
            O => \N__64342\,
            I => \N__64305\
        );

    \I__15535\ : Span12Mux_v
    port map (
            O => \N__64339\,
            I => \N__64305\
        );

    \I__15534\ : Span4Mux_h
    port map (
            O => \N__64336\,
            I => \N__64302\
        );

    \I__15533\ : Span4Mux_v
    port map (
            O => \N__64333\,
            I => \N__64299\
        );

    \I__15532\ : Span4Mux_h
    port map (
            O => \N__64328\,
            I => \N__64296\
        );

    \I__15531\ : LocalMux
    port map (
            O => \N__64323\,
            I => \N__64291\
        );

    \I__15530\ : Span4Mux_v
    port map (
            O => \N__64316\,
            I => \N__64291\
        );

    \I__15529\ : LocalMux
    port map (
            O => \N__64313\,
            I => \c0.n9_adj_4217\
        );

    \I__15528\ : LocalMux
    port map (
            O => \N__64310\,
            I => \c0.n9_adj_4217\
        );

    \I__15527\ : Odrv12
    port map (
            O => \N__64305\,
            I => \c0.n9_adj_4217\
        );

    \I__15526\ : Odrv4
    port map (
            O => \N__64302\,
            I => \c0.n9_adj_4217\
        );

    \I__15525\ : Odrv4
    port map (
            O => \N__64299\,
            I => \c0.n9_adj_4217\
        );

    \I__15524\ : Odrv4
    port map (
            O => \N__64296\,
            I => \c0.n9_adj_4217\
        );

    \I__15523\ : Odrv4
    port map (
            O => \N__64291\,
            I => \c0.n9_adj_4217\
        );

    \I__15522\ : CascadeMux
    port map (
            O => \N__64276\,
            I => \N__64272\
        );

    \I__15521\ : CascadeMux
    port map (
            O => \N__64275\,
            I => \N__64269\
        );

    \I__15520\ : InMux
    port map (
            O => \N__64272\,
            I => \N__64266\
        );

    \I__15519\ : InMux
    port map (
            O => \N__64269\,
            I => \N__64263\
        );

    \I__15518\ : LocalMux
    port map (
            O => \N__64266\,
            I => \c0.data_in_frame_28_6\
        );

    \I__15517\ : LocalMux
    port map (
            O => \N__64263\,
            I => \c0.data_in_frame_28_6\
        );

    \I__15516\ : InMux
    port map (
            O => \N__64258\,
            I => \N__64254\
        );

    \I__15515\ : InMux
    port map (
            O => \N__64257\,
            I => \N__64251\
        );

    \I__15514\ : LocalMux
    port map (
            O => \N__64254\,
            I => \N__64248\
        );

    \I__15513\ : LocalMux
    port map (
            O => \N__64251\,
            I => \N__64245\
        );

    \I__15512\ : Span4Mux_v
    port map (
            O => \N__64248\,
            I => \N__64239\
        );

    \I__15511\ : Span4Mux_h
    port map (
            O => \N__64245\,
            I => \N__64239\
        );

    \I__15510\ : InMux
    port map (
            O => \N__64244\,
            I => \N__64236\
        );

    \I__15509\ : Sp12to4
    port map (
            O => \N__64239\,
            I => \N__64231\
        );

    \I__15508\ : LocalMux
    port map (
            O => \N__64236\,
            I => \N__64231\
        );

    \I__15507\ : Odrv12
    port map (
            O => \N__64231\,
            I => \c0.n22105\
        );

    \I__15506\ : InMux
    port map (
            O => \N__64228\,
            I => \N__64225\
        );

    \I__15505\ : LocalMux
    port map (
            O => \N__64225\,
            I => \N__64221\
        );

    \I__15504\ : InMux
    port map (
            O => \N__64224\,
            I => \N__64216\
        );

    \I__15503\ : Span4Mux_h
    port map (
            O => \N__64221\,
            I => \N__64213\
        );

    \I__15502\ : InMux
    port map (
            O => \N__64220\,
            I => \N__64208\
        );

    \I__15501\ : InMux
    port map (
            O => \N__64219\,
            I => \N__64208\
        );

    \I__15500\ : LocalMux
    port map (
            O => \N__64216\,
            I => \N__64204\
        );

    \I__15499\ : Span4Mux_v
    port map (
            O => \N__64213\,
            I => \N__64199\
        );

    \I__15498\ : LocalMux
    port map (
            O => \N__64208\,
            I => \N__64199\
        );

    \I__15497\ : InMux
    port map (
            O => \N__64207\,
            I => \N__64196\
        );

    \I__15496\ : Odrv12
    port map (
            O => \N__64204\,
            I => \c0.n22849\
        );

    \I__15495\ : Odrv4
    port map (
            O => \N__64199\,
            I => \c0.n22849\
        );

    \I__15494\ : LocalMux
    port map (
            O => \N__64196\,
            I => \c0.n22849\
        );

    \I__15493\ : InMux
    port map (
            O => \N__64189\,
            I => \N__64186\
        );

    \I__15492\ : LocalMux
    port map (
            O => \N__64186\,
            I => \N__64183\
        );

    \I__15491\ : Span4Mux_h
    port map (
            O => \N__64183\,
            I => \N__64180\
        );

    \I__15490\ : Odrv4
    port map (
            O => \N__64180\,
            I => \c0.n20406\
        );

    \I__15489\ : InMux
    port map (
            O => \N__64177\,
            I => \N__64174\
        );

    \I__15488\ : LocalMux
    port map (
            O => \N__64174\,
            I => \N__64170\
        );

    \I__15487\ : InMux
    port map (
            O => \N__64173\,
            I => \N__64167\
        );

    \I__15486\ : Span12Mux_s10_h
    port map (
            O => \N__64170\,
            I => \N__64164\
        );

    \I__15485\ : LocalMux
    port map (
            O => \N__64167\,
            I => \N__64161\
        );

    \I__15484\ : Odrv12
    port map (
            O => \N__64164\,
            I => \c0.n5813\
        );

    \I__15483\ : Odrv4
    port map (
            O => \N__64161\,
            I => \c0.n5813\
        );

    \I__15482\ : InMux
    port map (
            O => \N__64156\,
            I => \N__64153\
        );

    \I__15481\ : LocalMux
    port map (
            O => \N__64153\,
            I => \N__64149\
        );

    \I__15480\ : InMux
    port map (
            O => \N__64152\,
            I => \N__64146\
        );

    \I__15479\ : Span4Mux_v
    port map (
            O => \N__64149\,
            I => \N__64141\
        );

    \I__15478\ : LocalMux
    port map (
            O => \N__64146\,
            I => \N__64141\
        );

    \I__15477\ : Span4Mux_h
    port map (
            O => \N__64141\,
            I => \N__64138\
        );

    \I__15476\ : Odrv4
    port map (
            O => \N__64138\,
            I => \c0.n21864\
        );

    \I__15475\ : CascadeMux
    port map (
            O => \N__64135\,
            I => \N__64132\
        );

    \I__15474\ : InMux
    port map (
            O => \N__64132\,
            I => \N__64129\
        );

    \I__15473\ : LocalMux
    port map (
            O => \N__64129\,
            I => \N__64126\
        );

    \I__15472\ : Odrv4
    port map (
            O => \N__64126\,
            I => \c0.n13768\
        );

    \I__15471\ : InMux
    port map (
            O => \N__64123\,
            I => \N__64119\
        );

    \I__15470\ : InMux
    port map (
            O => \N__64122\,
            I => \N__64116\
        );

    \I__15469\ : LocalMux
    port map (
            O => \N__64119\,
            I => \c0.n22458\
        );

    \I__15468\ : LocalMux
    port map (
            O => \N__64116\,
            I => \c0.n22458\
        );

    \I__15467\ : InMux
    port map (
            O => \N__64111\,
            I => \N__64106\
        );

    \I__15466\ : InMux
    port map (
            O => \N__64110\,
            I => \N__64101\
        );

    \I__15465\ : InMux
    port map (
            O => \N__64109\,
            I => \N__64101\
        );

    \I__15464\ : LocalMux
    port map (
            O => \N__64106\,
            I => \N__64098\
        );

    \I__15463\ : LocalMux
    port map (
            O => \N__64101\,
            I => \N__64095\
        );

    \I__15462\ : Span4Mux_v
    port map (
            O => \N__64098\,
            I => \N__64092\
        );

    \I__15461\ : Span4Mux_v
    port map (
            O => \N__64095\,
            I => \N__64089\
        );

    \I__15460\ : Odrv4
    port map (
            O => \N__64092\,
            I => \c0.n21114\
        );

    \I__15459\ : Odrv4
    port map (
            O => \N__64089\,
            I => \c0.n21114\
        );

    \I__15458\ : InMux
    port map (
            O => \N__64084\,
            I => \N__64081\
        );

    \I__15457\ : LocalMux
    port map (
            O => \N__64081\,
            I => \N__64078\
        );

    \I__15456\ : Span4Mux_v
    port map (
            O => \N__64078\,
            I => \N__64075\
        );

    \I__15455\ : Odrv4
    port map (
            O => \N__64075\,
            I => \c0.n18_adj_4246\
        );

    \I__15454\ : CascadeMux
    port map (
            O => \N__64072\,
            I => \c0.n21_cascade_\
        );

    \I__15453\ : InMux
    port map (
            O => \N__64069\,
            I => \N__64066\
        );

    \I__15452\ : LocalMux
    port map (
            O => \N__64066\,
            I => \N__64062\
        );

    \I__15451\ : InMux
    port map (
            O => \N__64065\,
            I => \N__64059\
        );

    \I__15450\ : Odrv4
    port map (
            O => \N__64062\,
            I => \c0.n22399\
        );

    \I__15449\ : LocalMux
    port map (
            O => \N__64059\,
            I => \c0.n22399\
        );

    \I__15448\ : InMux
    port map (
            O => \N__64054\,
            I => \N__64051\
        );

    \I__15447\ : LocalMux
    port map (
            O => \N__64051\,
            I => \c0.n24\
        );

    \I__15446\ : InMux
    port map (
            O => \N__64048\,
            I => \N__64045\
        );

    \I__15445\ : LocalMux
    port map (
            O => \N__64045\,
            I => \N__64042\
        );

    \I__15444\ : Span12Mux_s11_h
    port map (
            O => \N__64042\,
            I => \N__64039\
        );

    \I__15443\ : Odrv12
    port map (
            O => \N__64039\,
            I => \c0.n20\
        );

    \I__15442\ : InMux
    port map (
            O => \N__64036\,
            I => \N__64031\
        );

    \I__15441\ : CascadeMux
    port map (
            O => \N__64035\,
            I => \N__64027\
        );

    \I__15440\ : CascadeMux
    port map (
            O => \N__64034\,
            I => \N__64024\
        );

    \I__15439\ : LocalMux
    port map (
            O => \N__64031\,
            I => \N__64021\
        );

    \I__15438\ : CascadeMux
    port map (
            O => \N__64030\,
            I => \N__64018\
        );

    \I__15437\ : InMux
    port map (
            O => \N__64027\,
            I => \N__64014\
        );

    \I__15436\ : InMux
    port map (
            O => \N__64024\,
            I => \N__64011\
        );

    \I__15435\ : Span4Mux_h
    port map (
            O => \N__64021\,
            I => \N__64008\
        );

    \I__15434\ : InMux
    port map (
            O => \N__64018\,
            I => \N__64003\
        );

    \I__15433\ : InMux
    port map (
            O => \N__64017\,
            I => \N__64003\
        );

    \I__15432\ : LocalMux
    port map (
            O => \N__64014\,
            I => \c0.data_in_frame_17_1\
        );

    \I__15431\ : LocalMux
    port map (
            O => \N__64011\,
            I => \c0.data_in_frame_17_1\
        );

    \I__15430\ : Odrv4
    port map (
            O => \N__64008\,
            I => \c0.data_in_frame_17_1\
        );

    \I__15429\ : LocalMux
    port map (
            O => \N__64003\,
            I => \c0.data_in_frame_17_1\
        );

    \I__15428\ : CascadeMux
    port map (
            O => \N__63994\,
            I => \N__63991\
        );

    \I__15427\ : InMux
    port map (
            O => \N__63991\,
            I => \N__63988\
        );

    \I__15426\ : LocalMux
    port map (
            O => \N__63988\,
            I => \N__63985\
        );

    \I__15425\ : Span4Mux_v
    port map (
            O => \N__63985\,
            I => \N__63982\
        );

    \I__15424\ : Odrv4
    port map (
            O => \N__63982\,
            I => \c0.n16\
        );

    \I__15423\ : InMux
    port map (
            O => \N__63979\,
            I => \N__63976\
        );

    \I__15422\ : LocalMux
    port map (
            O => \N__63976\,
            I => \N__63973\
        );

    \I__15421\ : Span4Mux_v
    port map (
            O => \N__63973\,
            I => \N__63970\
        );

    \I__15420\ : Span4Mux_h
    port map (
            O => \N__63970\,
            I => \N__63966\
        );

    \I__15419\ : InMux
    port map (
            O => \N__63969\,
            I => \N__63963\
        );

    \I__15418\ : Odrv4
    port map (
            O => \N__63966\,
            I => \c0.n21979\
        );

    \I__15417\ : LocalMux
    port map (
            O => \N__63963\,
            I => \c0.n21979\
        );

    \I__15416\ : InMux
    port map (
            O => \N__63958\,
            I => \N__63953\
        );

    \I__15415\ : CascadeMux
    port map (
            O => \N__63957\,
            I => \N__63950\
        );

    \I__15414\ : InMux
    port map (
            O => \N__63956\,
            I => \N__63947\
        );

    \I__15413\ : LocalMux
    port map (
            O => \N__63953\,
            I => \N__63944\
        );

    \I__15412\ : InMux
    port map (
            O => \N__63950\,
            I => \N__63941\
        );

    \I__15411\ : LocalMux
    port map (
            O => \N__63947\,
            I => \N__63938\
        );

    \I__15410\ : Span4Mux_v
    port map (
            O => \N__63944\,
            I => \N__63935\
        );

    \I__15409\ : LocalMux
    port map (
            O => \N__63941\,
            I => \N__63932\
        );

    \I__15408\ : Span4Mux_h
    port map (
            O => \N__63938\,
            I => \N__63929\
        );

    \I__15407\ : Odrv4
    port map (
            O => \N__63935\,
            I => \c0.n23287\
        );

    \I__15406\ : Odrv12
    port map (
            O => \N__63932\,
            I => \c0.n23287\
        );

    \I__15405\ : Odrv4
    port map (
            O => \N__63929\,
            I => \c0.n23287\
        );

    \I__15404\ : CascadeMux
    port map (
            O => \N__63922\,
            I => \c0.n23287_cascade_\
        );

    \I__15403\ : InMux
    port map (
            O => \N__63919\,
            I => \N__63914\
        );

    \I__15402\ : InMux
    port map (
            O => \N__63918\,
            I => \N__63911\
        );

    \I__15401\ : CascadeMux
    port map (
            O => \N__63917\,
            I => \N__63908\
        );

    \I__15400\ : LocalMux
    port map (
            O => \N__63914\,
            I => \N__63905\
        );

    \I__15399\ : LocalMux
    port map (
            O => \N__63911\,
            I => \N__63902\
        );

    \I__15398\ : InMux
    port map (
            O => \N__63908\,
            I => \N__63897\
        );

    \I__15397\ : Span4Mux_v
    port map (
            O => \N__63905\,
            I => \N__63894\
        );

    \I__15396\ : Sp12to4
    port map (
            O => \N__63902\,
            I => \N__63891\
        );

    \I__15395\ : InMux
    port map (
            O => \N__63901\,
            I => \N__63886\
        );

    \I__15394\ : InMux
    port map (
            O => \N__63900\,
            I => \N__63886\
        );

    \I__15393\ : LocalMux
    port map (
            O => \N__63897\,
            I => \c0.data_in_frame_19_3\
        );

    \I__15392\ : Odrv4
    port map (
            O => \N__63894\,
            I => \c0.data_in_frame_19_3\
        );

    \I__15391\ : Odrv12
    port map (
            O => \N__63891\,
            I => \c0.data_in_frame_19_3\
        );

    \I__15390\ : LocalMux
    port map (
            O => \N__63886\,
            I => \c0.data_in_frame_19_3\
        );

    \I__15389\ : InMux
    port map (
            O => \N__63877\,
            I => \N__63873\
        );

    \I__15388\ : InMux
    port map (
            O => \N__63876\,
            I => \N__63870\
        );

    \I__15387\ : LocalMux
    port map (
            O => \N__63873\,
            I => \c0.n21921\
        );

    \I__15386\ : LocalMux
    port map (
            O => \N__63870\,
            I => \c0.n21921\
        );

    \I__15385\ : InMux
    port map (
            O => \N__63865\,
            I => \N__63856\
        );

    \I__15384\ : InMux
    port map (
            O => \N__63864\,
            I => \N__63846\
        );

    \I__15383\ : InMux
    port map (
            O => \N__63863\,
            I => \N__63843\
        );

    \I__15382\ : InMux
    port map (
            O => \N__63862\,
            I => \N__63840\
        );

    \I__15381\ : InMux
    port map (
            O => \N__63861\,
            I => \N__63835\
        );

    \I__15380\ : InMux
    port map (
            O => \N__63860\,
            I => \N__63835\
        );

    \I__15379\ : InMux
    port map (
            O => \N__63859\,
            I => \N__63832\
        );

    \I__15378\ : LocalMux
    port map (
            O => \N__63856\,
            I => \N__63827\
        );

    \I__15377\ : InMux
    port map (
            O => \N__63855\,
            I => \N__63820\
        );

    \I__15376\ : InMux
    port map (
            O => \N__63854\,
            I => \N__63820\
        );

    \I__15375\ : InMux
    port map (
            O => \N__63853\,
            I => \N__63817\
        );

    \I__15374\ : InMux
    port map (
            O => \N__63852\,
            I => \N__63810\
        );

    \I__15373\ : InMux
    port map (
            O => \N__63851\,
            I => \N__63807\
        );

    \I__15372\ : InMux
    port map (
            O => \N__63850\,
            I => \N__63804\
        );

    \I__15371\ : InMux
    port map (
            O => \N__63849\,
            I => \N__63801\
        );

    \I__15370\ : LocalMux
    port map (
            O => \N__63846\,
            I => \N__63797\
        );

    \I__15369\ : LocalMux
    port map (
            O => \N__63843\,
            I => \N__63794\
        );

    \I__15368\ : LocalMux
    port map (
            O => \N__63840\,
            I => \N__63790\
        );

    \I__15367\ : LocalMux
    port map (
            O => \N__63835\,
            I => \N__63785\
        );

    \I__15366\ : LocalMux
    port map (
            O => \N__63832\,
            I => \N__63785\
        );

    \I__15365\ : InMux
    port map (
            O => \N__63831\,
            I => \N__63782\
        );

    \I__15364\ : InMux
    port map (
            O => \N__63830\,
            I => \N__63776\
        );

    \I__15363\ : Span4Mux_h
    port map (
            O => \N__63827\,
            I => \N__63773\
        );

    \I__15362\ : InMux
    port map (
            O => \N__63826\,
            I => \N__63770\
        );

    \I__15361\ : InMux
    port map (
            O => \N__63825\,
            I => \N__63765\
        );

    \I__15360\ : LocalMux
    port map (
            O => \N__63820\,
            I => \N__63761\
        );

    \I__15359\ : LocalMux
    port map (
            O => \N__63817\,
            I => \N__63758\
        );

    \I__15358\ : InMux
    port map (
            O => \N__63816\,
            I => \N__63753\
        );

    \I__15357\ : InMux
    port map (
            O => \N__63815\,
            I => \N__63753\
        );

    \I__15356\ : InMux
    port map (
            O => \N__63814\,
            I => \N__63750\
        );

    \I__15355\ : InMux
    port map (
            O => \N__63813\,
            I => \N__63747\
        );

    \I__15354\ : LocalMux
    port map (
            O => \N__63810\,
            I => \N__63744\
        );

    \I__15353\ : LocalMux
    port map (
            O => \N__63807\,
            I => \N__63741\
        );

    \I__15352\ : LocalMux
    port map (
            O => \N__63804\,
            I => \N__63738\
        );

    \I__15351\ : LocalMux
    port map (
            O => \N__63801\,
            I => \N__63735\
        );

    \I__15350\ : InMux
    port map (
            O => \N__63800\,
            I => \N__63732\
        );

    \I__15349\ : Span4Mux_h
    port map (
            O => \N__63797\,
            I => \N__63727\
        );

    \I__15348\ : Span4Mux_v
    port map (
            O => \N__63794\,
            I => \N__63727\
        );

    \I__15347\ : InMux
    port map (
            O => \N__63793\,
            I => \N__63724\
        );

    \I__15346\ : Span4Mux_v
    port map (
            O => \N__63790\,
            I => \N__63717\
        );

    \I__15345\ : Span4Mux_v
    port map (
            O => \N__63785\,
            I => \N__63717\
        );

    \I__15344\ : LocalMux
    port map (
            O => \N__63782\,
            I => \N__63717\
        );

    \I__15343\ : InMux
    port map (
            O => \N__63781\,
            I => \N__63713\
        );

    \I__15342\ : InMux
    port map (
            O => \N__63780\,
            I => \N__63710\
        );

    \I__15341\ : InMux
    port map (
            O => \N__63779\,
            I => \N__63707\
        );

    \I__15340\ : LocalMux
    port map (
            O => \N__63776\,
            I => \N__63700\
        );

    \I__15339\ : Span4Mux_h
    port map (
            O => \N__63773\,
            I => \N__63700\
        );

    \I__15338\ : LocalMux
    port map (
            O => \N__63770\,
            I => \N__63700\
        );

    \I__15337\ : InMux
    port map (
            O => \N__63769\,
            I => \N__63695\
        );

    \I__15336\ : InMux
    port map (
            O => \N__63768\,
            I => \N__63695\
        );

    \I__15335\ : LocalMux
    port map (
            O => \N__63765\,
            I => \N__63692\
        );

    \I__15334\ : InMux
    port map (
            O => \N__63764\,
            I => \N__63689\
        );

    \I__15333\ : Span4Mux_v
    port map (
            O => \N__63761\,
            I => \N__63686\
        );

    \I__15332\ : Span4Mux_h
    port map (
            O => \N__63758\,
            I => \N__63679\
        );

    \I__15331\ : LocalMux
    port map (
            O => \N__63753\,
            I => \N__63679\
        );

    \I__15330\ : LocalMux
    port map (
            O => \N__63750\,
            I => \N__63679\
        );

    \I__15329\ : LocalMux
    port map (
            O => \N__63747\,
            I => \N__63672\
        );

    \I__15328\ : Span4Mux_v
    port map (
            O => \N__63744\,
            I => \N__63672\
        );

    \I__15327\ : Span4Mux_v
    port map (
            O => \N__63741\,
            I => \N__63672\
        );

    \I__15326\ : Span4Mux_h
    port map (
            O => \N__63738\,
            I => \N__63665\
        );

    \I__15325\ : Span4Mux_v
    port map (
            O => \N__63735\,
            I => \N__63665\
        );

    \I__15324\ : LocalMux
    port map (
            O => \N__63732\,
            I => \N__63665\
        );

    \I__15323\ : Sp12to4
    port map (
            O => \N__63727\,
            I => \N__63660\
        );

    \I__15322\ : LocalMux
    port map (
            O => \N__63724\,
            I => \N__63660\
        );

    \I__15321\ : Span4Mux_h
    port map (
            O => \N__63717\,
            I => \N__63657\
        );

    \I__15320\ : InMux
    port map (
            O => \N__63716\,
            I => \N__63654\
        );

    \I__15319\ : LocalMux
    port map (
            O => \N__63713\,
            I => \N__63651\
        );

    \I__15318\ : LocalMux
    port map (
            O => \N__63710\,
            I => \N__63644\
        );

    \I__15317\ : LocalMux
    port map (
            O => \N__63707\,
            I => \N__63644\
        );

    \I__15316\ : Span4Mux_h
    port map (
            O => \N__63700\,
            I => \N__63644\
        );

    \I__15315\ : LocalMux
    port map (
            O => \N__63695\,
            I => \N__63638\
        );

    \I__15314\ : Span4Mux_v
    port map (
            O => \N__63692\,
            I => \N__63638\
        );

    \I__15313\ : LocalMux
    port map (
            O => \N__63689\,
            I => \N__63633\
        );

    \I__15312\ : Span4Mux_h
    port map (
            O => \N__63686\,
            I => \N__63633\
        );

    \I__15311\ : Span4Mux_h
    port map (
            O => \N__63679\,
            I => \N__63626\
        );

    \I__15310\ : Span4Mux_h
    port map (
            O => \N__63672\,
            I => \N__63626\
        );

    \I__15309\ : Span4Mux_v
    port map (
            O => \N__63665\,
            I => \N__63626\
        );

    \I__15308\ : Span12Mux_h
    port map (
            O => \N__63660\,
            I => \N__63623\
        );

    \I__15307\ : Sp12to4
    port map (
            O => \N__63657\,
            I => \N__63620\
        );

    \I__15306\ : LocalMux
    port map (
            O => \N__63654\,
            I => \N__63617\
        );

    \I__15305\ : Span4Mux_h
    port map (
            O => \N__63651\,
            I => \N__63612\
        );

    \I__15304\ : Span4Mux_v
    port map (
            O => \N__63644\,
            I => \N__63612\
        );

    \I__15303\ : InMux
    port map (
            O => \N__63643\,
            I => \N__63609\
        );

    \I__15302\ : Span4Mux_v
    port map (
            O => \N__63638\,
            I => \N__63606\
        );

    \I__15301\ : Span4Mux_v
    port map (
            O => \N__63633\,
            I => \N__63603\
        );

    \I__15300\ : Span4Mux_v
    port map (
            O => \N__63626\,
            I => \N__63600\
        );

    \I__15299\ : Span12Mux_v
    port map (
            O => \N__63623\,
            I => \N__63597\
        );

    \I__15298\ : Span12Mux_s10_v
    port map (
            O => \N__63620\,
            I => \N__63592\
        );

    \I__15297\ : Span12Mux_h
    port map (
            O => \N__63617\,
            I => \N__63592\
        );

    \I__15296\ : Span4Mux_v
    port map (
            O => \N__63612\,
            I => \N__63589\
        );

    \I__15295\ : LocalMux
    port map (
            O => \N__63609\,
            I => rx_data_1
        );

    \I__15294\ : Odrv4
    port map (
            O => \N__63606\,
            I => rx_data_1
        );

    \I__15293\ : Odrv4
    port map (
            O => \N__63603\,
            I => rx_data_1
        );

    \I__15292\ : Odrv4
    port map (
            O => \N__63600\,
            I => rx_data_1
        );

    \I__15291\ : Odrv12
    port map (
            O => \N__63597\,
            I => rx_data_1
        );

    \I__15290\ : Odrv12
    port map (
            O => \N__63592\,
            I => rx_data_1
        );

    \I__15289\ : Odrv4
    port map (
            O => \N__63589\,
            I => rx_data_1
        );

    \I__15288\ : CascadeMux
    port map (
            O => \N__63574\,
            I => \N__63570\
        );

    \I__15287\ : InMux
    port map (
            O => \N__63573\,
            I => \N__63567\
        );

    \I__15286\ : InMux
    port map (
            O => \N__63570\,
            I => \N__63564\
        );

    \I__15285\ : LocalMux
    port map (
            O => \N__63567\,
            I => \N__63561\
        );

    \I__15284\ : LocalMux
    port map (
            O => \N__63564\,
            I => \N__63555\
        );

    \I__15283\ : Span4Mux_v
    port map (
            O => \N__63561\,
            I => \N__63555\
        );

    \I__15282\ : InMux
    port map (
            O => \N__63560\,
            I => \N__63552\
        );

    \I__15281\ : Odrv4
    port map (
            O => \N__63555\,
            I => \c0.data_in_frame_24_0\
        );

    \I__15280\ : LocalMux
    port map (
            O => \N__63552\,
            I => \c0.data_in_frame_24_0\
        );

    \I__15279\ : InMux
    port map (
            O => \N__63547\,
            I => \N__63543\
        );

    \I__15278\ : CascadeMux
    port map (
            O => \N__63546\,
            I => \N__63540\
        );

    \I__15277\ : LocalMux
    port map (
            O => \N__63543\,
            I => \N__63535\
        );

    \I__15276\ : InMux
    port map (
            O => \N__63540\,
            I => \N__63532\
        );

    \I__15275\ : CascadeMux
    port map (
            O => \N__63539\,
            I => \N__63529\
        );

    \I__15274\ : InMux
    port map (
            O => \N__63538\,
            I => \N__63526\
        );

    \I__15273\ : Span4Mux_h
    port map (
            O => \N__63535\,
            I => \N__63523\
        );

    \I__15272\ : LocalMux
    port map (
            O => \N__63532\,
            I => \N__63520\
        );

    \I__15271\ : InMux
    port map (
            O => \N__63529\,
            I => \N__63517\
        );

    \I__15270\ : LocalMux
    port map (
            O => \N__63526\,
            I => \N__63510\
        );

    \I__15269\ : Span4Mux_h
    port map (
            O => \N__63523\,
            I => \N__63510\
        );

    \I__15268\ : Span4Mux_h
    port map (
            O => \N__63520\,
            I => \N__63510\
        );

    \I__15267\ : LocalMux
    port map (
            O => \N__63517\,
            I => \c0.data_in_frame_24_5\
        );

    \I__15266\ : Odrv4
    port map (
            O => \N__63510\,
            I => \c0.data_in_frame_24_5\
        );

    \I__15265\ : CascadeMux
    port map (
            O => \N__63505\,
            I => \N__63502\
        );

    \I__15264\ : InMux
    port map (
            O => \N__63502\,
            I => \N__63498\
        );

    \I__15263\ : InMux
    port map (
            O => \N__63501\,
            I => \N__63495\
        );

    \I__15262\ : LocalMux
    port map (
            O => \N__63498\,
            I => \c0.n13320\
        );

    \I__15261\ : LocalMux
    port map (
            O => \N__63495\,
            I => \c0.n13320\
        );

    \I__15260\ : InMux
    port map (
            O => \N__63490\,
            I => \N__63487\
        );

    \I__15259\ : LocalMux
    port map (
            O => \N__63487\,
            I => \N__63482\
        );

    \I__15258\ : InMux
    port map (
            O => \N__63486\,
            I => \N__63479\
        );

    \I__15257\ : InMux
    port map (
            O => \N__63485\,
            I => \N__63476\
        );

    \I__15256\ : Span4Mux_h
    port map (
            O => \N__63482\,
            I => \N__63470\
        );

    \I__15255\ : LocalMux
    port map (
            O => \N__63479\,
            I => \N__63470\
        );

    \I__15254\ : LocalMux
    port map (
            O => \N__63476\,
            I => \N__63467\
        );

    \I__15253\ : CascadeMux
    port map (
            O => \N__63475\,
            I => \N__63464\
        );

    \I__15252\ : Span4Mux_v
    port map (
            O => \N__63470\,
            I => \N__63459\
        );

    \I__15251\ : Span4Mux_v
    port map (
            O => \N__63467\,
            I => \N__63459\
        );

    \I__15250\ : InMux
    port map (
            O => \N__63464\,
            I => \N__63456\
        );

    \I__15249\ : Sp12to4
    port map (
            O => \N__63459\,
            I => \N__63450\
        );

    \I__15248\ : LocalMux
    port map (
            O => \N__63456\,
            I => \N__63450\
        );

    \I__15247\ : InMux
    port map (
            O => \N__63455\,
            I => \N__63447\
        );

    \I__15246\ : Span12Mux_h
    port map (
            O => \N__63450\,
            I => \N__63444\
        );

    \I__15245\ : LocalMux
    port map (
            O => \N__63447\,
            I => data_in_frame_22_5
        );

    \I__15244\ : Odrv12
    port map (
            O => \N__63444\,
            I => data_in_frame_22_5
        );

    \I__15243\ : InMux
    port map (
            O => \N__63439\,
            I => \N__63436\
        );

    \I__15242\ : LocalMux
    port map (
            O => \N__63436\,
            I => \N__63433\
        );

    \I__15241\ : Span4Mux_h
    port map (
            O => \N__63433\,
            I => \N__63429\
        );

    \I__15240\ : InMux
    port map (
            O => \N__63432\,
            I => \N__63426\
        );

    \I__15239\ : Odrv4
    port map (
            O => \N__63429\,
            I => \c0.n22255\
        );

    \I__15238\ : LocalMux
    port map (
            O => \N__63426\,
            I => \c0.n22255\
        );

    \I__15237\ : CascadeMux
    port map (
            O => \N__63421\,
            I => \N__63418\
        );

    \I__15236\ : InMux
    port map (
            O => \N__63418\,
            I => \N__63413\
        );

    \I__15235\ : CascadeMux
    port map (
            O => \N__63417\,
            I => \N__63410\
        );

    \I__15234\ : CascadeMux
    port map (
            O => \N__63416\,
            I => \N__63407\
        );

    \I__15233\ : LocalMux
    port map (
            O => \N__63413\,
            I => \N__63404\
        );

    \I__15232\ : InMux
    port map (
            O => \N__63410\,
            I => \N__63401\
        );

    \I__15231\ : InMux
    port map (
            O => \N__63407\,
            I => \N__63398\
        );

    \I__15230\ : Span4Mux_h
    port map (
            O => \N__63404\,
            I => \N__63395\
        );

    \I__15229\ : LocalMux
    port map (
            O => \N__63401\,
            I => \c0.data_in_frame_19_1\
        );

    \I__15228\ : LocalMux
    port map (
            O => \N__63398\,
            I => \c0.data_in_frame_19_1\
        );

    \I__15227\ : Odrv4
    port map (
            O => \N__63395\,
            I => \c0.data_in_frame_19_1\
        );

    \I__15226\ : InMux
    port map (
            O => \N__63388\,
            I => \N__63384\
        );

    \I__15225\ : InMux
    port map (
            O => \N__63387\,
            I => \N__63381\
        );

    \I__15224\ : LocalMux
    port map (
            O => \N__63384\,
            I => \N__63378\
        );

    \I__15223\ : LocalMux
    port map (
            O => \N__63381\,
            I => \N__63375\
        );

    \I__15222\ : Span4Mux_h
    port map (
            O => \N__63378\,
            I => \N__63372\
        );

    \I__15221\ : Span4Mux_h
    port map (
            O => \N__63375\,
            I => \N__63369\
        );

    \I__15220\ : Odrv4
    port map (
            O => \N__63372\,
            I => \c0.n22084\
        );

    \I__15219\ : Odrv4
    port map (
            O => \N__63369\,
            I => \c0.n22084\
        );

    \I__15218\ : InMux
    port map (
            O => \N__63364\,
            I => \N__63361\
        );

    \I__15217\ : LocalMux
    port map (
            O => \N__63361\,
            I => \c0.n22364\
        );

    \I__15216\ : CascadeMux
    port map (
            O => \N__63358\,
            I => \N__63352\
        );

    \I__15215\ : InMux
    port map (
            O => \N__63357\,
            I => \N__63348\
        );

    \I__15214\ : InMux
    port map (
            O => \N__63356\,
            I => \N__63345\
        );

    \I__15213\ : CascadeMux
    port map (
            O => \N__63355\,
            I => \N__63342\
        );

    \I__15212\ : InMux
    port map (
            O => \N__63352\,
            I => \N__63339\
        );

    \I__15211\ : InMux
    port map (
            O => \N__63351\,
            I => \N__63336\
        );

    \I__15210\ : LocalMux
    port map (
            O => \N__63348\,
            I => \N__63331\
        );

    \I__15209\ : LocalMux
    port map (
            O => \N__63345\,
            I => \N__63331\
        );

    \I__15208\ : InMux
    port map (
            O => \N__63342\,
            I => \N__63328\
        );

    \I__15207\ : LocalMux
    port map (
            O => \N__63339\,
            I => \N__63321\
        );

    \I__15206\ : LocalMux
    port map (
            O => \N__63336\,
            I => \N__63321\
        );

    \I__15205\ : Span4Mux_h
    port map (
            O => \N__63331\,
            I => \N__63321\
        );

    \I__15204\ : LocalMux
    port map (
            O => \N__63328\,
            I => \c0.data_in_frame_19_7\
        );

    \I__15203\ : Odrv4
    port map (
            O => \N__63321\,
            I => \c0.data_in_frame_19_7\
        );

    \I__15202\ : InMux
    port map (
            O => \N__63316\,
            I => \N__63313\
        );

    \I__15201\ : LocalMux
    port map (
            O => \N__63313\,
            I => \c0.n15\
        );

    \I__15200\ : CascadeMux
    port map (
            O => \N__63310\,
            I => \N__63305\
        );

    \I__15199\ : CascadeMux
    port map (
            O => \N__63309\,
            I => \N__63301\
        );

    \I__15198\ : InMux
    port map (
            O => \N__63308\,
            I => \N__63296\
        );

    \I__15197\ : InMux
    port map (
            O => \N__63305\,
            I => \N__63296\
        );

    \I__15196\ : InMux
    port map (
            O => \N__63304\,
            I => \N__63292\
        );

    \I__15195\ : InMux
    port map (
            O => \N__63301\,
            I => \N__63289\
        );

    \I__15194\ : LocalMux
    port map (
            O => \N__63296\,
            I => \N__63286\
        );

    \I__15193\ : InMux
    port map (
            O => \N__63295\,
            I => \N__63283\
        );

    \I__15192\ : LocalMux
    port map (
            O => \N__63292\,
            I => \N__63280\
        );

    \I__15191\ : LocalMux
    port map (
            O => \N__63289\,
            I => \N__63275\
        );

    \I__15190\ : Span4Mux_v
    port map (
            O => \N__63286\,
            I => \N__63275\
        );

    \I__15189\ : LocalMux
    port map (
            O => \N__63283\,
            I => \c0.data_in_frame_20_5\
        );

    \I__15188\ : Odrv12
    port map (
            O => \N__63280\,
            I => \c0.data_in_frame_20_5\
        );

    \I__15187\ : Odrv4
    port map (
            O => \N__63275\,
            I => \c0.data_in_frame_20_5\
        );

    \I__15186\ : CascadeMux
    port map (
            O => \N__63268\,
            I => \N__63264\
        );

    \I__15185\ : InMux
    port map (
            O => \N__63267\,
            I => \N__63261\
        );

    \I__15184\ : InMux
    port map (
            O => \N__63264\,
            I => \N__63258\
        );

    \I__15183\ : LocalMux
    port map (
            O => \N__63261\,
            I => \N__63254\
        );

    \I__15182\ : LocalMux
    port map (
            O => \N__63258\,
            I => \N__63251\
        );

    \I__15181\ : InMux
    port map (
            O => \N__63257\,
            I => \N__63248\
        );

    \I__15180\ : Span4Mux_h
    port map (
            O => \N__63254\,
            I => \N__63245\
        );

    \I__15179\ : Odrv4
    port map (
            O => \N__63251\,
            I => \c0.data_in_frame_23_0\
        );

    \I__15178\ : LocalMux
    port map (
            O => \N__63248\,
            I => \c0.data_in_frame_23_0\
        );

    \I__15177\ : Odrv4
    port map (
            O => \N__63245\,
            I => \c0.data_in_frame_23_0\
        );

    \I__15176\ : InMux
    port map (
            O => \N__63238\,
            I => \N__63235\
        );

    \I__15175\ : LocalMux
    port map (
            O => \N__63235\,
            I => \N__63232\
        );

    \I__15174\ : Span4Mux_h
    port map (
            O => \N__63232\,
            I => \N__63229\
        );

    \I__15173\ : Odrv4
    port map (
            O => \N__63229\,
            I => \c0.n26_adj_4281\
        );

    \I__15172\ : InMux
    port map (
            O => \N__63226\,
            I => \N__63222\
        );

    \I__15171\ : InMux
    port map (
            O => \N__63225\,
            I => \N__63219\
        );

    \I__15170\ : LocalMux
    port map (
            O => \N__63222\,
            I => \N__63213\
        );

    \I__15169\ : LocalMux
    port map (
            O => \N__63219\,
            I => \N__63210\
        );

    \I__15168\ : InMux
    port map (
            O => \N__63218\,
            I => \N__63207\
        );

    \I__15167\ : CascadeMux
    port map (
            O => \N__63217\,
            I => \N__63201\
        );

    \I__15166\ : CascadeMux
    port map (
            O => \N__63216\,
            I => \N__63198\
        );

    \I__15165\ : Span4Mux_v
    port map (
            O => \N__63213\,
            I => \N__63195\
        );

    \I__15164\ : Span4Mux_h
    port map (
            O => \N__63210\,
            I => \N__63192\
        );

    \I__15163\ : LocalMux
    port map (
            O => \N__63207\,
            I => \N__63189\
        );

    \I__15162\ : InMux
    port map (
            O => \N__63206\,
            I => \N__63185\
        );

    \I__15161\ : InMux
    port map (
            O => \N__63205\,
            I => \N__63182\
        );

    \I__15160\ : InMux
    port map (
            O => \N__63204\,
            I => \N__63179\
        );

    \I__15159\ : InMux
    port map (
            O => \N__63201\,
            I => \N__63165\
        );

    \I__15158\ : InMux
    port map (
            O => \N__63198\,
            I => \N__63165\
        );

    \I__15157\ : Span4Mux_h
    port map (
            O => \N__63195\,
            I => \N__63162\
        );

    \I__15156\ : Span4Mux_v
    port map (
            O => \N__63192\,
            I => \N__63156\
        );

    \I__15155\ : Span4Mux_h
    port map (
            O => \N__63189\,
            I => \N__63156\
        );

    \I__15154\ : InMux
    port map (
            O => \N__63188\,
            I => \N__63153\
        );

    \I__15153\ : LocalMux
    port map (
            O => \N__63185\,
            I => \N__63150\
        );

    \I__15152\ : LocalMux
    port map (
            O => \N__63182\,
            I => \N__63147\
        );

    \I__15151\ : LocalMux
    port map (
            O => \N__63179\,
            I => \N__63140\
        );

    \I__15150\ : InMux
    port map (
            O => \N__63178\,
            I => \N__63136\
        );

    \I__15149\ : InMux
    port map (
            O => \N__63177\,
            I => \N__63133\
        );

    \I__15148\ : InMux
    port map (
            O => \N__63176\,
            I => \N__63130\
        );

    \I__15147\ : InMux
    port map (
            O => \N__63175\,
            I => \N__63125\
        );

    \I__15146\ : InMux
    port map (
            O => \N__63174\,
            I => \N__63125\
        );

    \I__15145\ : InMux
    port map (
            O => \N__63173\,
            I => \N__63120\
        );

    \I__15144\ : CascadeMux
    port map (
            O => \N__63172\,
            I => \N__63117\
        );

    \I__15143\ : InMux
    port map (
            O => \N__63171\,
            I => \N__63114\
        );

    \I__15142\ : InMux
    port map (
            O => \N__63170\,
            I => \N__63111\
        );

    \I__15141\ : LocalMux
    port map (
            O => \N__63165\,
            I => \N__63108\
        );

    \I__15140\ : Span4Mux_h
    port map (
            O => \N__63162\,
            I => \N__63103\
        );

    \I__15139\ : InMux
    port map (
            O => \N__63161\,
            I => \N__63100\
        );

    \I__15138\ : Span4Mux_h
    port map (
            O => \N__63156\,
            I => \N__63093\
        );

    \I__15137\ : LocalMux
    port map (
            O => \N__63153\,
            I => \N__63093\
        );

    \I__15136\ : Span4Mux_v
    port map (
            O => \N__63150\,
            I => \N__63093\
        );

    \I__15135\ : Span4Mux_v
    port map (
            O => \N__63147\,
            I => \N__63089\
        );

    \I__15134\ : InMux
    port map (
            O => \N__63146\,
            I => \N__63086\
        );

    \I__15133\ : InMux
    port map (
            O => \N__63145\,
            I => \N__63083\
        );

    \I__15132\ : InMux
    port map (
            O => \N__63144\,
            I => \N__63078\
        );

    \I__15131\ : InMux
    port map (
            O => \N__63143\,
            I => \N__63078\
        );

    \I__15130\ : Span4Mux_v
    port map (
            O => \N__63140\,
            I => \N__63075\
        );

    \I__15129\ : InMux
    port map (
            O => \N__63139\,
            I => \N__63072\
        );

    \I__15128\ : LocalMux
    port map (
            O => \N__63136\,
            I => \N__63069\
        );

    \I__15127\ : LocalMux
    port map (
            O => \N__63133\,
            I => \N__63062\
        );

    \I__15126\ : LocalMux
    port map (
            O => \N__63130\,
            I => \N__63062\
        );

    \I__15125\ : LocalMux
    port map (
            O => \N__63125\,
            I => \N__63062\
        );

    \I__15124\ : InMux
    port map (
            O => \N__63124\,
            I => \N__63059\
        );

    \I__15123\ : InMux
    port map (
            O => \N__63123\,
            I => \N__63055\
        );

    \I__15122\ : LocalMux
    port map (
            O => \N__63120\,
            I => \N__63052\
        );

    \I__15121\ : InMux
    port map (
            O => \N__63117\,
            I => \N__63049\
        );

    \I__15120\ : LocalMux
    port map (
            O => \N__63114\,
            I => \N__63046\
        );

    \I__15119\ : LocalMux
    port map (
            O => \N__63111\,
            I => \N__63041\
        );

    \I__15118\ : Span4Mux_v
    port map (
            O => \N__63108\,
            I => \N__63041\
        );

    \I__15117\ : InMux
    port map (
            O => \N__63107\,
            I => \N__63038\
        );

    \I__15116\ : InMux
    port map (
            O => \N__63106\,
            I => \N__63035\
        );

    \I__15115\ : Span4Mux_v
    port map (
            O => \N__63103\,
            I => \N__63030\
        );

    \I__15114\ : LocalMux
    port map (
            O => \N__63100\,
            I => \N__63030\
        );

    \I__15113\ : Span4Mux_v
    port map (
            O => \N__63093\,
            I => \N__63027\
        );

    \I__15112\ : InMux
    port map (
            O => \N__63092\,
            I => \N__63024\
        );

    \I__15111\ : Span4Mux_v
    port map (
            O => \N__63089\,
            I => \N__63021\
        );

    \I__15110\ : LocalMux
    port map (
            O => \N__63086\,
            I => \N__63018\
        );

    \I__15109\ : LocalMux
    port map (
            O => \N__63083\,
            I => \N__63015\
        );

    \I__15108\ : LocalMux
    port map (
            O => \N__63078\,
            I => \N__63010\
        );

    \I__15107\ : Span4Mux_v
    port map (
            O => \N__63075\,
            I => \N__63010\
        );

    \I__15106\ : LocalMux
    port map (
            O => \N__63072\,
            I => \N__63001\
        );

    \I__15105\ : Span4Mux_v
    port map (
            O => \N__63069\,
            I => \N__63001\
        );

    \I__15104\ : Span4Mux_v
    port map (
            O => \N__63062\,
            I => \N__63001\
        );

    \I__15103\ : LocalMux
    port map (
            O => \N__63059\,
            I => \N__63001\
        );

    \I__15102\ : InMux
    port map (
            O => \N__63058\,
            I => \N__62997\
        );

    \I__15101\ : LocalMux
    port map (
            O => \N__63055\,
            I => \N__62990\
        );

    \I__15100\ : Span4Mux_h
    port map (
            O => \N__63052\,
            I => \N__62990\
        );

    \I__15099\ : LocalMux
    port map (
            O => \N__63049\,
            I => \N__62990\
        );

    \I__15098\ : Span4Mux_h
    port map (
            O => \N__63046\,
            I => \N__62985\
        );

    \I__15097\ : Span4Mux_h
    port map (
            O => \N__63041\,
            I => \N__62985\
        );

    \I__15096\ : LocalMux
    port map (
            O => \N__63038\,
            I => \N__62982\
        );

    \I__15095\ : LocalMux
    port map (
            O => \N__63035\,
            I => \N__62979\
        );

    \I__15094\ : Span4Mux_v
    port map (
            O => \N__63030\,
            I => \N__62976\
        );

    \I__15093\ : Sp12to4
    port map (
            O => \N__63027\,
            I => \N__62972\
        );

    \I__15092\ : LocalMux
    port map (
            O => \N__63024\,
            I => \N__62967\
        );

    \I__15091\ : Span4Mux_v
    port map (
            O => \N__63021\,
            I => \N__62967\
        );

    \I__15090\ : Span4Mux_v
    port map (
            O => \N__63018\,
            I => \N__62964\
        );

    \I__15089\ : Span4Mux_v
    port map (
            O => \N__63015\,
            I => \N__62961\
        );

    \I__15088\ : Span4Mux_h
    port map (
            O => \N__63010\,
            I => \N__62956\
        );

    \I__15087\ : Span4Mux_v
    port map (
            O => \N__63001\,
            I => \N__62956\
        );

    \I__15086\ : InMux
    port map (
            O => \N__63000\,
            I => \N__62953\
        );

    \I__15085\ : LocalMux
    port map (
            O => \N__62997\,
            I => \N__62944\
        );

    \I__15084\ : Span4Mux_h
    port map (
            O => \N__62990\,
            I => \N__62944\
        );

    \I__15083\ : Span4Mux_v
    port map (
            O => \N__62985\,
            I => \N__62944\
        );

    \I__15082\ : Span4Mux_v
    port map (
            O => \N__62982\,
            I => \N__62944\
        );

    \I__15081\ : Span4Mux_v
    port map (
            O => \N__62979\,
            I => \N__62941\
        );

    \I__15080\ : Span4Mux_v
    port map (
            O => \N__62976\,
            I => \N__62938\
        );

    \I__15079\ : InMux
    port map (
            O => \N__62975\,
            I => \N__62935\
        );

    \I__15078\ : Span12Mux_h
    port map (
            O => \N__62972\,
            I => \N__62932\
        );

    \I__15077\ : Sp12to4
    port map (
            O => \N__62967\,
            I => \N__62929\
        );

    \I__15076\ : Span4Mux_v
    port map (
            O => \N__62964\,
            I => \N__62922\
        );

    \I__15075\ : Span4Mux_h
    port map (
            O => \N__62961\,
            I => \N__62922\
        );

    \I__15074\ : Span4Mux_v
    port map (
            O => \N__62956\,
            I => \N__62922\
        );

    \I__15073\ : LocalMux
    port map (
            O => \N__62953\,
            I => \N__62913\
        );

    \I__15072\ : Span4Mux_v
    port map (
            O => \N__62944\,
            I => \N__62913\
        );

    \I__15071\ : Span4Mux_v
    port map (
            O => \N__62941\,
            I => \N__62913\
        );

    \I__15070\ : Span4Mux_v
    port map (
            O => \N__62938\,
            I => \N__62913\
        );

    \I__15069\ : LocalMux
    port map (
            O => \N__62935\,
            I => rx_data_4
        );

    \I__15068\ : Odrv12
    port map (
            O => \N__62932\,
            I => rx_data_4
        );

    \I__15067\ : Odrv12
    port map (
            O => \N__62929\,
            I => rx_data_4
        );

    \I__15066\ : Odrv4
    port map (
            O => \N__62922\,
            I => rx_data_4
        );

    \I__15065\ : Odrv4
    port map (
            O => \N__62913\,
            I => rx_data_4
        );

    \I__15064\ : InMux
    port map (
            O => \N__62902\,
            I => \N__62897\
        );

    \I__15063\ : CascadeMux
    port map (
            O => \N__62901\,
            I => \N__62894\
        );

    \I__15062\ : InMux
    port map (
            O => \N__62900\,
            I => \N__62890\
        );

    \I__15061\ : LocalMux
    port map (
            O => \N__62897\,
            I => \N__62887\
        );

    \I__15060\ : InMux
    port map (
            O => \N__62894\,
            I => \N__62884\
        );

    \I__15059\ : InMux
    port map (
            O => \N__62893\,
            I => \N__62881\
        );

    \I__15058\ : LocalMux
    port map (
            O => \N__62890\,
            I => \N__62874\
        );

    \I__15057\ : Span4Mux_v
    port map (
            O => \N__62887\,
            I => \N__62874\
        );

    \I__15056\ : LocalMux
    port map (
            O => \N__62884\,
            I => \N__62874\
        );

    \I__15055\ : LocalMux
    port map (
            O => \N__62881\,
            I => \c0.data_in_frame_18_3\
        );

    \I__15054\ : Odrv4
    port map (
            O => \N__62874\,
            I => \c0.data_in_frame_18_3\
        );

    \I__15053\ : InMux
    port map (
            O => \N__62869\,
            I => \N__62866\
        );

    \I__15052\ : LocalMux
    port map (
            O => \N__62866\,
            I => \c0.n22095\
        );

    \I__15051\ : InMux
    port map (
            O => \N__62863\,
            I => \N__62860\
        );

    \I__15050\ : LocalMux
    port map (
            O => \N__62860\,
            I => \c0.n21124\
        );

    \I__15049\ : CascadeMux
    port map (
            O => \N__62857\,
            I => \c0.n22095_cascade_\
        );

    \I__15048\ : InMux
    port map (
            O => \N__62854\,
            I => \N__62851\
        );

    \I__15047\ : LocalMux
    port map (
            O => \N__62851\,
            I => \N__62847\
        );

    \I__15046\ : InMux
    port map (
            O => \N__62850\,
            I => \N__62844\
        );

    \I__15045\ : Odrv4
    port map (
            O => \N__62847\,
            I => \c0.n14143\
        );

    \I__15044\ : LocalMux
    port map (
            O => \N__62844\,
            I => \c0.n14143\
        );

    \I__15043\ : InMux
    port map (
            O => \N__62839\,
            I => \N__62836\
        );

    \I__15042\ : LocalMux
    port map (
            O => \N__62836\,
            I => \N__62833\
        );

    \I__15041\ : Span4Mux_h
    port map (
            O => \N__62833\,
            I => \N__62830\
        );

    \I__15040\ : Odrv4
    port map (
            O => \N__62830\,
            I => \c0.n29\
        );

    \I__15039\ : CascadeMux
    port map (
            O => \N__62827\,
            I => \N__62823\
        );

    \I__15038\ : InMux
    port map (
            O => \N__62826\,
            I => \N__62819\
        );

    \I__15037\ : InMux
    port map (
            O => \N__62823\,
            I => \N__62816\
        );

    \I__15036\ : CascadeMux
    port map (
            O => \N__62822\,
            I => \N__62812\
        );

    \I__15035\ : LocalMux
    port map (
            O => \N__62819\,
            I => \N__62807\
        );

    \I__15034\ : LocalMux
    port map (
            O => \N__62816\,
            I => \N__62807\
        );

    \I__15033\ : InMux
    port map (
            O => \N__62815\,
            I => \N__62804\
        );

    \I__15032\ : InMux
    port map (
            O => \N__62812\,
            I => \N__62801\
        );

    \I__15031\ : Span12Mux_v
    port map (
            O => \N__62807\,
            I => \N__62798\
        );

    \I__15030\ : LocalMux
    port map (
            O => \N__62804\,
            I => data_in_frame_22_0
        );

    \I__15029\ : LocalMux
    port map (
            O => \N__62801\,
            I => data_in_frame_22_0
        );

    \I__15028\ : Odrv12
    port map (
            O => \N__62798\,
            I => data_in_frame_22_0
        );

    \I__15027\ : InMux
    port map (
            O => \N__62791\,
            I => \N__62788\
        );

    \I__15026\ : LocalMux
    port map (
            O => \N__62788\,
            I => \N__62784\
        );

    \I__15025\ : InMux
    port map (
            O => \N__62787\,
            I => \N__62781\
        );

    \I__15024\ : Span4Mux_v
    port map (
            O => \N__62784\,
            I => \N__62778\
        );

    \I__15023\ : LocalMux
    port map (
            O => \N__62781\,
            I => \N__62775\
        );

    \I__15022\ : Odrv4
    port map (
            O => \N__62778\,
            I => \c0.n22267\
        );

    \I__15021\ : Odrv4
    port map (
            O => \N__62775\,
            I => \c0.n22267\
        );

    \I__15020\ : InMux
    port map (
            O => \N__62770\,
            I => \N__62767\
        );

    \I__15019\ : LocalMux
    port map (
            O => \N__62767\,
            I => \N__62762\
        );

    \I__15018\ : InMux
    port map (
            O => \N__62766\,
            I => \N__62757\
        );

    \I__15017\ : InMux
    port map (
            O => \N__62765\,
            I => \N__62757\
        );

    \I__15016\ : Odrv4
    port map (
            O => \N__62762\,
            I => \c0.data_in_frame_20_4\
        );

    \I__15015\ : LocalMux
    port map (
            O => \N__62757\,
            I => \c0.data_in_frame_20_4\
        );

    \I__15014\ : CascadeMux
    port map (
            O => \N__62752\,
            I => \N__62748\
        );

    \I__15013\ : CascadeMux
    port map (
            O => \N__62751\,
            I => \N__62745\
        );

    \I__15012\ : InMux
    port map (
            O => \N__62748\,
            I => \N__62742\
        );

    \I__15011\ : InMux
    port map (
            O => \N__62745\,
            I => \N__62739\
        );

    \I__15010\ : LocalMux
    port map (
            O => \N__62742\,
            I => \N__62736\
        );

    \I__15009\ : LocalMux
    port map (
            O => \N__62739\,
            I => \N__62733\
        );

    \I__15008\ : Span4Mux_v
    port map (
            O => \N__62736\,
            I => \N__62730\
        );

    \I__15007\ : Span4Mux_v
    port map (
            O => \N__62733\,
            I => \N__62726\
        );

    \I__15006\ : Span4Mux_h
    port map (
            O => \N__62730\,
            I => \N__62723\
        );

    \I__15005\ : InMux
    port map (
            O => \N__62729\,
            I => \N__62720\
        );

    \I__15004\ : Span4Mux_h
    port map (
            O => \N__62726\,
            I => \N__62717\
        );

    \I__15003\ : Span4Mux_v
    port map (
            O => \N__62723\,
            I => \N__62714\
        );

    \I__15002\ : LocalMux
    port map (
            O => \N__62720\,
            I => data_in_frame_22_6
        );

    \I__15001\ : Odrv4
    port map (
            O => \N__62717\,
            I => data_in_frame_22_6
        );

    \I__15000\ : Odrv4
    port map (
            O => \N__62714\,
            I => data_in_frame_22_6
        );

    \I__14999\ : InMux
    port map (
            O => \N__62707\,
            I => \N__62703\
        );

    \I__14998\ : CascadeMux
    port map (
            O => \N__62706\,
            I => \N__62699\
        );

    \I__14997\ : LocalMux
    port map (
            O => \N__62703\,
            I => \N__62695\
        );

    \I__14996\ : InMux
    port map (
            O => \N__62702\,
            I => \N__62690\
        );

    \I__14995\ : InMux
    port map (
            O => \N__62699\,
            I => \N__62690\
        );

    \I__14994\ : InMux
    port map (
            O => \N__62698\,
            I => \N__62687\
        );

    \I__14993\ : Span4Mux_v
    port map (
            O => \N__62695\,
            I => \N__62682\
        );

    \I__14992\ : LocalMux
    port map (
            O => \N__62690\,
            I => \N__62682\
        );

    \I__14991\ : LocalMux
    port map (
            O => \N__62687\,
            I => \c0.n20246\
        );

    \I__14990\ : Odrv4
    port map (
            O => \N__62682\,
            I => \c0.n20246\
        );

    \I__14989\ : InMux
    port map (
            O => \N__62677\,
            I => \N__62673\
        );

    \I__14988\ : CascadeMux
    port map (
            O => \N__62676\,
            I => \N__62668\
        );

    \I__14987\ : LocalMux
    port map (
            O => \N__62673\,
            I => \N__62665\
        );

    \I__14986\ : InMux
    port map (
            O => \N__62672\,
            I => \N__62662\
        );

    \I__14985\ : InMux
    port map (
            O => \N__62671\,
            I => \N__62658\
        );

    \I__14984\ : InMux
    port map (
            O => \N__62668\,
            I => \N__62655\
        );

    \I__14983\ : Span4Mux_v
    port map (
            O => \N__62665\,
            I => \N__62650\
        );

    \I__14982\ : LocalMux
    port map (
            O => \N__62662\,
            I => \N__62650\
        );

    \I__14981\ : InMux
    port map (
            O => \N__62661\,
            I => \N__62647\
        );

    \I__14980\ : LocalMux
    port map (
            O => \N__62658\,
            I => \N__62644\
        );

    \I__14979\ : LocalMux
    port map (
            O => \N__62655\,
            I => \c0.data_in_frame_13_6\
        );

    \I__14978\ : Odrv4
    port map (
            O => \N__62650\,
            I => \c0.data_in_frame_13_6\
        );

    \I__14977\ : LocalMux
    port map (
            O => \N__62647\,
            I => \c0.data_in_frame_13_6\
        );

    \I__14976\ : Odrv12
    port map (
            O => \N__62644\,
            I => \c0.data_in_frame_13_6\
        );

    \I__14975\ : InMux
    port map (
            O => \N__62635\,
            I => \N__62632\
        );

    \I__14974\ : LocalMux
    port map (
            O => \N__62632\,
            I => \N__62627\
        );

    \I__14973\ : InMux
    port map (
            O => \N__62631\,
            I => \N__62624\
        );

    \I__14972\ : CascadeMux
    port map (
            O => \N__62630\,
            I => \N__62621\
        );

    \I__14971\ : Span4Mux_h
    port map (
            O => \N__62627\,
            I => \N__62618\
        );

    \I__14970\ : LocalMux
    port map (
            O => \N__62624\,
            I => \N__62615\
        );

    \I__14969\ : InMux
    port map (
            O => \N__62621\,
            I => \N__62612\
        );

    \I__14968\ : Span4Mux_v
    port map (
            O => \N__62618\,
            I => \N__62609\
        );

    \I__14967\ : Span4Mux_v
    port map (
            O => \N__62615\,
            I => \N__62606\
        );

    \I__14966\ : LocalMux
    port map (
            O => \N__62612\,
            I => \c0.data_in_frame_26_5\
        );

    \I__14965\ : Odrv4
    port map (
            O => \N__62609\,
            I => \c0.data_in_frame_26_5\
        );

    \I__14964\ : Odrv4
    port map (
            O => \N__62606\,
            I => \c0.data_in_frame_26_5\
        );

    \I__14963\ : InMux
    port map (
            O => \N__62599\,
            I => \N__62595\
        );

    \I__14962\ : CascadeMux
    port map (
            O => \N__62598\,
            I => \N__62592\
        );

    \I__14961\ : LocalMux
    port map (
            O => \N__62595\,
            I => \N__62587\
        );

    \I__14960\ : InMux
    port map (
            O => \N__62592\,
            I => \N__62584\
        );

    \I__14959\ : CascadeMux
    port map (
            O => \N__62591\,
            I => \N__62581\
        );

    \I__14958\ : InMux
    port map (
            O => \N__62590\,
            I => \N__62578\
        );

    \I__14957\ : Span4Mux_v
    port map (
            O => \N__62587\,
            I => \N__62573\
        );

    \I__14956\ : LocalMux
    port map (
            O => \N__62584\,
            I => \N__62573\
        );

    \I__14955\ : InMux
    port map (
            O => \N__62581\,
            I => \N__62570\
        );

    \I__14954\ : LocalMux
    port map (
            O => \N__62578\,
            I => \N__62567\
        );

    \I__14953\ : Span4Mux_h
    port map (
            O => \N__62573\,
            I => \N__62564\
        );

    \I__14952\ : LocalMux
    port map (
            O => \N__62570\,
            I => \c0.data_in_frame_21_6\
        );

    \I__14951\ : Odrv12
    port map (
            O => \N__62567\,
            I => \c0.data_in_frame_21_6\
        );

    \I__14950\ : Odrv4
    port map (
            O => \N__62564\,
            I => \c0.data_in_frame_21_6\
        );

    \I__14949\ : InMux
    port map (
            O => \N__62557\,
            I => \N__62551\
        );

    \I__14948\ : InMux
    port map (
            O => \N__62556\,
            I => \N__62546\
        );

    \I__14947\ : InMux
    port map (
            O => \N__62555\,
            I => \N__62546\
        );

    \I__14946\ : InMux
    port map (
            O => \N__62554\,
            I => \N__62535\
        );

    \I__14945\ : LocalMux
    port map (
            O => \N__62551\,
            I => \N__62532\
        );

    \I__14944\ : LocalMux
    port map (
            O => \N__62546\,
            I => \N__62519\
        );

    \I__14943\ : InMux
    port map (
            O => \N__62545\,
            I => \N__62514\
        );

    \I__14942\ : InMux
    port map (
            O => \N__62544\,
            I => \N__62514\
        );

    \I__14941\ : InMux
    port map (
            O => \N__62543\,
            I => \N__62511\
        );

    \I__14940\ : InMux
    port map (
            O => \N__62542\,
            I => \N__62487\
        );

    \I__14939\ : InMux
    port map (
            O => \N__62541\,
            I => \N__62484\
        );

    \I__14938\ : InMux
    port map (
            O => \N__62540\,
            I => \N__62477\
        );

    \I__14937\ : InMux
    port map (
            O => \N__62539\,
            I => \N__62477\
        );

    \I__14936\ : InMux
    port map (
            O => \N__62538\,
            I => \N__62477\
        );

    \I__14935\ : LocalMux
    port map (
            O => \N__62535\,
            I => \N__62472\
        );

    \I__14934\ : Span4Mux_v
    port map (
            O => \N__62532\,
            I => \N__62472\
        );

    \I__14933\ : InMux
    port map (
            O => \N__62531\,
            I => \N__62465\
        );

    \I__14932\ : InMux
    port map (
            O => \N__62530\,
            I => \N__62465\
        );

    \I__14931\ : InMux
    port map (
            O => \N__62529\,
            I => \N__62465\
        );

    \I__14930\ : InMux
    port map (
            O => \N__62528\,
            I => \N__62458\
        );

    \I__14929\ : InMux
    port map (
            O => \N__62527\,
            I => \N__62458\
        );

    \I__14928\ : InMux
    port map (
            O => \N__62526\,
            I => \N__62458\
        );

    \I__14927\ : InMux
    port map (
            O => \N__62525\,
            I => \N__62449\
        );

    \I__14926\ : InMux
    port map (
            O => \N__62524\,
            I => \N__62449\
        );

    \I__14925\ : InMux
    port map (
            O => \N__62523\,
            I => \N__62449\
        );

    \I__14924\ : InMux
    port map (
            O => \N__62522\,
            I => \N__62449\
        );

    \I__14923\ : Span4Mux_v
    port map (
            O => \N__62519\,
            I => \N__62444\
        );

    \I__14922\ : LocalMux
    port map (
            O => \N__62514\,
            I => \N__62444\
        );

    \I__14921\ : LocalMux
    port map (
            O => \N__62511\,
            I => \N__62441\
        );

    \I__14920\ : InMux
    port map (
            O => \N__62510\,
            I => \N__62436\
        );

    \I__14919\ : InMux
    port map (
            O => \N__62509\,
            I => \N__62436\
        );

    \I__14918\ : InMux
    port map (
            O => \N__62508\,
            I => \N__62433\
        );

    \I__14917\ : InMux
    port map (
            O => \N__62507\,
            I => \N__62422\
        );

    \I__14916\ : InMux
    port map (
            O => \N__62506\,
            I => \N__62422\
        );

    \I__14915\ : InMux
    port map (
            O => \N__62505\,
            I => \N__62417\
        );

    \I__14914\ : InMux
    port map (
            O => \N__62504\,
            I => \N__62417\
        );

    \I__14913\ : InMux
    port map (
            O => \N__62503\,
            I => \N__62412\
        );

    \I__14912\ : InMux
    port map (
            O => \N__62502\,
            I => \N__62412\
        );

    \I__14911\ : InMux
    port map (
            O => \N__62501\,
            I => \N__62409\
        );

    \I__14910\ : InMux
    port map (
            O => \N__62500\,
            I => \N__62406\
        );

    \I__14909\ : InMux
    port map (
            O => \N__62499\,
            I => \N__62397\
        );

    \I__14908\ : InMux
    port map (
            O => \N__62498\,
            I => \N__62397\
        );

    \I__14907\ : InMux
    port map (
            O => \N__62497\,
            I => \N__62397\
        );

    \I__14906\ : InMux
    port map (
            O => \N__62496\,
            I => \N__62397\
        );

    \I__14905\ : InMux
    port map (
            O => \N__62495\,
            I => \N__62383\
        );

    \I__14904\ : InMux
    port map (
            O => \N__62494\,
            I => \N__62383\
        );

    \I__14903\ : InMux
    port map (
            O => \N__62493\,
            I => \N__62383\
        );

    \I__14902\ : InMux
    port map (
            O => \N__62492\,
            I => \N__62383\
        );

    \I__14901\ : InMux
    port map (
            O => \N__62491\,
            I => \N__62383\
        );

    \I__14900\ : InMux
    port map (
            O => \N__62490\,
            I => \N__62383\
        );

    \I__14899\ : LocalMux
    port map (
            O => \N__62487\,
            I => \N__62380\
        );

    \I__14898\ : LocalMux
    port map (
            O => \N__62484\,
            I => \N__62365\
        );

    \I__14897\ : LocalMux
    port map (
            O => \N__62477\,
            I => \N__62365\
        );

    \I__14896\ : Span4Mux_h
    port map (
            O => \N__62472\,
            I => \N__62365\
        );

    \I__14895\ : LocalMux
    port map (
            O => \N__62465\,
            I => \N__62365\
        );

    \I__14894\ : LocalMux
    port map (
            O => \N__62458\,
            I => \N__62360\
        );

    \I__14893\ : LocalMux
    port map (
            O => \N__62449\,
            I => \N__62360\
        );

    \I__14892\ : Span4Mux_v
    port map (
            O => \N__62444\,
            I => \N__62357\
        );

    \I__14891\ : Span4Mux_v
    port map (
            O => \N__62441\,
            I => \N__62352\
        );

    \I__14890\ : LocalMux
    port map (
            O => \N__62436\,
            I => \N__62352\
        );

    \I__14889\ : LocalMux
    port map (
            O => \N__62433\,
            I => \N__62348\
        );

    \I__14888\ : InMux
    port map (
            O => \N__62432\,
            I => \N__62343\
        );

    \I__14887\ : InMux
    port map (
            O => \N__62431\,
            I => \N__62343\
        );

    \I__14886\ : InMux
    port map (
            O => \N__62430\,
            I => \N__62340\
        );

    \I__14885\ : InMux
    port map (
            O => \N__62429\,
            I => \N__62333\
        );

    \I__14884\ : InMux
    port map (
            O => \N__62428\,
            I => \N__62333\
        );

    \I__14883\ : InMux
    port map (
            O => \N__62427\,
            I => \N__62333\
        );

    \I__14882\ : LocalMux
    port map (
            O => \N__62422\,
            I => \N__62330\
        );

    \I__14881\ : LocalMux
    port map (
            O => \N__62417\,
            I => \N__62327\
        );

    \I__14880\ : LocalMux
    port map (
            O => \N__62412\,
            I => \N__62324\
        );

    \I__14879\ : LocalMux
    port map (
            O => \N__62409\,
            I => \N__62317\
        );

    \I__14878\ : LocalMux
    port map (
            O => \N__62406\,
            I => \N__62317\
        );

    \I__14877\ : LocalMux
    port map (
            O => \N__62397\,
            I => \N__62317\
        );

    \I__14876\ : InMux
    port map (
            O => \N__62396\,
            I => \N__62314\
        );

    \I__14875\ : LocalMux
    port map (
            O => \N__62383\,
            I => \N__62311\
        );

    \I__14874\ : Span4Mux_v
    port map (
            O => \N__62380\,
            I => \N__62308\
        );

    \I__14873\ : InMux
    port map (
            O => \N__62379\,
            I => \N__62305\
        );

    \I__14872\ : InMux
    port map (
            O => \N__62378\,
            I => \N__62302\
        );

    \I__14871\ : InMux
    port map (
            O => \N__62377\,
            I => \N__62299\
        );

    \I__14870\ : InMux
    port map (
            O => \N__62376\,
            I => \N__62292\
        );

    \I__14869\ : InMux
    port map (
            O => \N__62375\,
            I => \N__62292\
        );

    \I__14868\ : InMux
    port map (
            O => \N__62374\,
            I => \N__62292\
        );

    \I__14867\ : Span4Mux_v
    port map (
            O => \N__62365\,
            I => \N__62289\
        );

    \I__14866\ : Span4Mux_v
    port map (
            O => \N__62360\,
            I => \N__62282\
        );

    \I__14865\ : Span4Mux_h
    port map (
            O => \N__62357\,
            I => \N__62282\
        );

    \I__14864\ : Span4Mux_v
    port map (
            O => \N__62352\,
            I => \N__62282\
        );

    \I__14863\ : InMux
    port map (
            O => \N__62351\,
            I => \N__62279\
        );

    \I__14862\ : Span4Mux_v
    port map (
            O => \N__62348\,
            I => \N__62276\
        );

    \I__14861\ : LocalMux
    port map (
            O => \N__62343\,
            I => \N__62273\
        );

    \I__14860\ : LocalMux
    port map (
            O => \N__62340\,
            I => \N__62260\
        );

    \I__14859\ : LocalMux
    port map (
            O => \N__62333\,
            I => \N__62260\
        );

    \I__14858\ : Span4Mux_h
    port map (
            O => \N__62330\,
            I => \N__62260\
        );

    \I__14857\ : Span4Mux_v
    port map (
            O => \N__62327\,
            I => \N__62260\
        );

    \I__14856\ : Span4Mux_h
    port map (
            O => \N__62324\,
            I => \N__62260\
        );

    \I__14855\ : Span4Mux_v
    port map (
            O => \N__62317\,
            I => \N__62260\
        );

    \I__14854\ : LocalMux
    port map (
            O => \N__62314\,
            I => \N__62257\
        );

    \I__14853\ : Span4Mux_v
    port map (
            O => \N__62311\,
            I => \N__62252\
        );

    \I__14852\ : Span4Mux_h
    port map (
            O => \N__62308\,
            I => \N__62252\
        );

    \I__14851\ : LocalMux
    port map (
            O => \N__62305\,
            I => \N__62249\
        );

    \I__14850\ : LocalMux
    port map (
            O => \N__62302\,
            I => \N__62236\
        );

    \I__14849\ : LocalMux
    port map (
            O => \N__62299\,
            I => \N__62236\
        );

    \I__14848\ : LocalMux
    port map (
            O => \N__62292\,
            I => \N__62236\
        );

    \I__14847\ : Sp12to4
    port map (
            O => \N__62289\,
            I => \N__62236\
        );

    \I__14846\ : Sp12to4
    port map (
            O => \N__62282\,
            I => \N__62236\
        );

    \I__14845\ : LocalMux
    port map (
            O => \N__62279\,
            I => \N__62236\
        );

    \I__14844\ : Span4Mux_h
    port map (
            O => \N__62276\,
            I => \N__62233\
        );

    \I__14843\ : Span12Mux_v
    port map (
            O => \N__62273\,
            I => \N__62230\
        );

    \I__14842\ : Span4Mux_h
    port map (
            O => \N__62260\,
            I => \N__62227\
        );

    \I__14841\ : Span4Mux_v
    port map (
            O => \N__62257\,
            I => \N__62222\
        );

    \I__14840\ : Span4Mux_v
    port map (
            O => \N__62252\,
            I => \N__62222\
        );

    \I__14839\ : Sp12to4
    port map (
            O => \N__62249\,
            I => \N__62217\
        );

    \I__14838\ : Span12Mux_h
    port map (
            O => \N__62236\,
            I => \N__62217\
        );

    \I__14837\ : Odrv4
    port map (
            O => \N__62233\,
            I => \c0.n21749\
        );

    \I__14836\ : Odrv12
    port map (
            O => \N__62230\,
            I => \c0.n21749\
        );

    \I__14835\ : Odrv4
    port map (
            O => \N__62227\,
            I => \c0.n21749\
        );

    \I__14834\ : Odrv4
    port map (
            O => \N__62222\,
            I => \c0.n21749\
        );

    \I__14833\ : Odrv12
    port map (
            O => \N__62217\,
            I => \c0.n21749\
        );

    \I__14832\ : CascadeMux
    port map (
            O => \N__62206\,
            I => \N__62199\
        );

    \I__14831\ : CascadeMux
    port map (
            O => \N__62205\,
            I => \N__62194\
        );

    \I__14830\ : CascadeMux
    port map (
            O => \N__62204\,
            I => \N__62191\
        );

    \I__14829\ : CascadeMux
    port map (
            O => \N__62203\,
            I => \N__62178\
        );

    \I__14828\ : CascadeMux
    port map (
            O => \N__62202\,
            I => \N__62174\
        );

    \I__14827\ : InMux
    port map (
            O => \N__62199\,
            I => \N__62171\
        );

    \I__14826\ : InMux
    port map (
            O => \N__62198\,
            I => \N__62168\
        );

    \I__14825\ : InMux
    port map (
            O => \N__62197\,
            I => \N__62161\
        );

    \I__14824\ : InMux
    port map (
            O => \N__62194\,
            I => \N__62161\
        );

    \I__14823\ : InMux
    port map (
            O => \N__62191\,
            I => \N__62157\
        );

    \I__14822\ : CascadeMux
    port map (
            O => \N__62190\,
            I => \N__62154\
        );

    \I__14821\ : InMux
    port map (
            O => \N__62189\,
            I => \N__62151\
        );

    \I__14820\ : InMux
    port map (
            O => \N__62188\,
            I => \N__62145\
        );

    \I__14819\ : InMux
    port map (
            O => \N__62187\,
            I => \N__62142\
        );

    \I__14818\ : InMux
    port map (
            O => \N__62186\,
            I => \N__62137\
        );

    \I__14817\ : InMux
    port map (
            O => \N__62185\,
            I => \N__62137\
        );

    \I__14816\ : InMux
    port map (
            O => \N__62184\,
            I => \N__62132\
        );

    \I__14815\ : InMux
    port map (
            O => \N__62183\,
            I => \N__62132\
        );

    \I__14814\ : InMux
    port map (
            O => \N__62182\,
            I => \N__62125\
        );

    \I__14813\ : InMux
    port map (
            O => \N__62181\,
            I => \N__62125\
        );

    \I__14812\ : InMux
    port map (
            O => \N__62178\,
            I => \N__62125\
        );

    \I__14811\ : CascadeMux
    port map (
            O => \N__62177\,
            I => \N__62122\
        );

    \I__14810\ : InMux
    port map (
            O => \N__62174\,
            I => \N__62117\
        );

    \I__14809\ : LocalMux
    port map (
            O => \N__62171\,
            I => \N__62112\
        );

    \I__14808\ : LocalMux
    port map (
            O => \N__62168\,
            I => \N__62112\
        );

    \I__14807\ : InMux
    port map (
            O => \N__62167\,
            I => \N__62107\
        );

    \I__14806\ : InMux
    port map (
            O => \N__62166\,
            I => \N__62107\
        );

    \I__14805\ : LocalMux
    port map (
            O => \N__62161\,
            I => \N__62104\
        );

    \I__14804\ : InMux
    port map (
            O => \N__62160\,
            I => \N__62101\
        );

    \I__14803\ : LocalMux
    port map (
            O => \N__62157\,
            I => \N__62098\
        );

    \I__14802\ : InMux
    port map (
            O => \N__62154\,
            I => \N__62095\
        );

    \I__14801\ : LocalMux
    port map (
            O => \N__62151\,
            I => \N__62092\
        );

    \I__14800\ : InMux
    port map (
            O => \N__62150\,
            I => \N__62089\
        );

    \I__14799\ : CascadeMux
    port map (
            O => \N__62149\,
            I => \N__62083\
        );

    \I__14798\ : InMux
    port map (
            O => \N__62148\,
            I => \N__62080\
        );

    \I__14797\ : LocalMux
    port map (
            O => \N__62145\,
            I => \N__62077\
        );

    \I__14796\ : LocalMux
    port map (
            O => \N__62142\,
            I => \N__62074\
        );

    \I__14795\ : LocalMux
    port map (
            O => \N__62137\,
            I => \N__62071\
        );

    \I__14794\ : LocalMux
    port map (
            O => \N__62132\,
            I => \N__62068\
        );

    \I__14793\ : LocalMux
    port map (
            O => \N__62125\,
            I => \N__62065\
        );

    \I__14792\ : InMux
    port map (
            O => \N__62122\,
            I => \N__62062\
        );

    \I__14791\ : CascadeMux
    port map (
            O => \N__62121\,
            I => \N__62059\
        );

    \I__14790\ : InMux
    port map (
            O => \N__62120\,
            I => \N__62055\
        );

    \I__14789\ : LocalMux
    port map (
            O => \N__62117\,
            I => \N__62052\
        );

    \I__14788\ : Span4Mux_v
    port map (
            O => \N__62112\,
            I => \N__62049\
        );

    \I__14787\ : LocalMux
    port map (
            O => \N__62107\,
            I => \N__62046\
        );

    \I__14786\ : Span4Mux_h
    port map (
            O => \N__62104\,
            I => \N__62043\
        );

    \I__14785\ : LocalMux
    port map (
            O => \N__62101\,
            I => \N__62038\
        );

    \I__14784\ : Span4Mux_h
    port map (
            O => \N__62098\,
            I => \N__62038\
        );

    \I__14783\ : LocalMux
    port map (
            O => \N__62095\,
            I => \N__62033\
        );

    \I__14782\ : Span4Mux_h
    port map (
            O => \N__62092\,
            I => \N__62033\
        );

    \I__14781\ : LocalMux
    port map (
            O => \N__62089\,
            I => \N__62030\
        );

    \I__14780\ : InMux
    port map (
            O => \N__62088\,
            I => \N__62027\
        );

    \I__14779\ : InMux
    port map (
            O => \N__62087\,
            I => \N__62024\
        );

    \I__14778\ : InMux
    port map (
            O => \N__62086\,
            I => \N__62021\
        );

    \I__14777\ : InMux
    port map (
            O => \N__62083\,
            I => \N__62018\
        );

    \I__14776\ : LocalMux
    port map (
            O => \N__62080\,
            I => \N__62015\
        );

    \I__14775\ : Span4Mux_v
    port map (
            O => \N__62077\,
            I => \N__62010\
        );

    \I__14774\ : Span4Mux_h
    port map (
            O => \N__62074\,
            I => \N__62010\
        );

    \I__14773\ : Span4Mux_h
    port map (
            O => \N__62071\,
            I => \N__62007\
        );

    \I__14772\ : Span4Mux_h
    port map (
            O => \N__62068\,
            I => \N__62004\
        );

    \I__14771\ : Span4Mux_h
    port map (
            O => \N__62065\,
            I => \N__62001\
        );

    \I__14770\ : LocalMux
    port map (
            O => \N__62062\,
            I => \N__61998\
        );

    \I__14769\ : InMux
    port map (
            O => \N__62059\,
            I => \N__61995\
        );

    \I__14768\ : InMux
    port map (
            O => \N__62058\,
            I => \N__61992\
        );

    \I__14767\ : LocalMux
    port map (
            O => \N__62055\,
            I => \N__61989\
        );

    \I__14766\ : Span4Mux_h
    port map (
            O => \N__62052\,
            I => \N__61982\
        );

    \I__14765\ : Span4Mux_h
    port map (
            O => \N__62049\,
            I => \N__61982\
        );

    \I__14764\ : Span4Mux_h
    port map (
            O => \N__62046\,
            I => \N__61982\
        );

    \I__14763\ : Span4Mux_h
    port map (
            O => \N__62043\,
            I => \N__61977\
        );

    \I__14762\ : Span4Mux_h
    port map (
            O => \N__62038\,
            I => \N__61977\
        );

    \I__14761\ : Span4Mux_v
    port map (
            O => \N__62033\,
            I => \N__61974\
        );

    \I__14760\ : Span4Mux_h
    port map (
            O => \N__62030\,
            I => \N__61971\
        );

    \I__14759\ : LocalMux
    port map (
            O => \N__62027\,
            I => \N__61966\
        );

    \I__14758\ : LocalMux
    port map (
            O => \N__62024\,
            I => \N__61961\
        );

    \I__14757\ : LocalMux
    port map (
            O => \N__62021\,
            I => \N__61961\
        );

    \I__14756\ : LocalMux
    port map (
            O => \N__62018\,
            I => \N__61950\
        );

    \I__14755\ : Span4Mux_h
    port map (
            O => \N__62015\,
            I => \N__61950\
        );

    \I__14754\ : Span4Mux_h
    port map (
            O => \N__62010\,
            I => \N__61950\
        );

    \I__14753\ : Span4Mux_h
    port map (
            O => \N__62007\,
            I => \N__61950\
        );

    \I__14752\ : Span4Mux_v
    port map (
            O => \N__62004\,
            I => \N__61950\
        );

    \I__14751\ : Span4Mux_v
    port map (
            O => \N__62001\,
            I => \N__61945\
        );

    \I__14750\ : Span4Mux_h
    port map (
            O => \N__61998\,
            I => \N__61945\
        );

    \I__14749\ : LocalMux
    port map (
            O => \N__61995\,
            I => \N__61934\
        );

    \I__14748\ : LocalMux
    port map (
            O => \N__61992\,
            I => \N__61934\
        );

    \I__14747\ : Span12Mux_s9_h
    port map (
            O => \N__61989\,
            I => \N__61934\
        );

    \I__14746\ : Sp12to4
    port map (
            O => \N__61982\,
            I => \N__61934\
        );

    \I__14745\ : Sp12to4
    port map (
            O => \N__61977\,
            I => \N__61934\
        );

    \I__14744\ : Span4Mux_v
    port map (
            O => \N__61974\,
            I => \N__61929\
        );

    \I__14743\ : Span4Mux_v
    port map (
            O => \N__61971\,
            I => \N__61929\
        );

    \I__14742\ : InMux
    port map (
            O => \N__61970\,
            I => \N__61924\
        );

    \I__14741\ : InMux
    port map (
            O => \N__61969\,
            I => \N__61924\
        );

    \I__14740\ : Span4Mux_h
    port map (
            O => \N__61966\,
            I => \N__61921\
        );

    \I__14739\ : Span4Mux_v
    port map (
            O => \N__61961\,
            I => \N__61918\
        );

    \I__14738\ : Span4Mux_v
    port map (
            O => \N__61950\,
            I => \N__61915\
        );

    \I__14737\ : Sp12to4
    port map (
            O => \N__61945\,
            I => \N__61910\
        );

    \I__14736\ : Span12Mux_v
    port map (
            O => \N__61934\,
            I => \N__61910\
        );

    \I__14735\ : Span4Mux_h
    port map (
            O => \N__61929\,
            I => \N__61907\
        );

    \I__14734\ : LocalMux
    port map (
            O => \N__61924\,
            I => \c0.n9_adj_4237\
        );

    \I__14733\ : Odrv4
    port map (
            O => \N__61921\,
            I => \c0.n9_adj_4237\
        );

    \I__14732\ : Odrv4
    port map (
            O => \N__61918\,
            I => \c0.n9_adj_4237\
        );

    \I__14731\ : Odrv4
    port map (
            O => \N__61915\,
            I => \c0.n9_adj_4237\
        );

    \I__14730\ : Odrv12
    port map (
            O => \N__61910\,
            I => \c0.n9_adj_4237\
        );

    \I__14729\ : Odrv4
    port map (
            O => \N__61907\,
            I => \c0.n9_adj_4237\
        );

    \I__14728\ : CascadeMux
    port map (
            O => \N__61894\,
            I => \N__61891\
        );

    \I__14727\ : InMux
    port map (
            O => \N__61891\,
            I => \N__61888\
        );

    \I__14726\ : LocalMux
    port map (
            O => \N__61888\,
            I => \N__61881\
        );

    \I__14725\ : InMux
    port map (
            O => \N__61887\,
            I => \N__61878\
        );

    \I__14724\ : InMux
    port map (
            O => \N__61886\,
            I => \N__61875\
        );

    \I__14723\ : InMux
    port map (
            O => \N__61885\,
            I => \N__61872\
        );

    \I__14722\ : InMux
    port map (
            O => \N__61884\,
            I => \N__61869\
        );

    \I__14721\ : Span12Mux_v
    port map (
            O => \N__61881\,
            I => \N__61866\
        );

    \I__14720\ : LocalMux
    port map (
            O => \N__61878\,
            I => \N__61861\
        );

    \I__14719\ : LocalMux
    port map (
            O => \N__61875\,
            I => \N__61861\
        );

    \I__14718\ : LocalMux
    port map (
            O => \N__61872\,
            I => \c0.data_in_frame_13_7\
        );

    \I__14717\ : LocalMux
    port map (
            O => \N__61869\,
            I => \c0.data_in_frame_13_7\
        );

    \I__14716\ : Odrv12
    port map (
            O => \N__61866\,
            I => \c0.data_in_frame_13_7\
        );

    \I__14715\ : Odrv12
    port map (
            O => \N__61861\,
            I => \c0.data_in_frame_13_7\
        );

    \I__14714\ : InMux
    port map (
            O => \N__61852\,
            I => \N__61849\
        );

    \I__14713\ : LocalMux
    port map (
            O => \N__61849\,
            I => \N__61845\
        );

    \I__14712\ : InMux
    port map (
            O => \N__61848\,
            I => \N__61842\
        );

    \I__14711\ : Span4Mux_v
    port map (
            O => \N__61845\,
            I => \N__61839\
        );

    \I__14710\ : LocalMux
    port map (
            O => \N__61842\,
            I => \N__61836\
        );

    \I__14709\ : Span4Mux_v
    port map (
            O => \N__61839\,
            I => \N__61833\
        );

    \I__14708\ : Odrv12
    port map (
            O => \N__61836\,
            I => \c0.n22388\
        );

    \I__14707\ : Odrv4
    port map (
            O => \N__61833\,
            I => \c0.n22388\
        );

    \I__14706\ : InMux
    port map (
            O => \N__61828\,
            I => \N__61825\
        );

    \I__14705\ : LocalMux
    port map (
            O => \N__61825\,
            I => \N__61820\
        );

    \I__14704\ : InMux
    port map (
            O => \N__61824\,
            I => \N__61817\
        );

    \I__14703\ : CascadeMux
    port map (
            O => \N__61823\,
            I => \N__61814\
        );

    \I__14702\ : Span4Mux_v
    port map (
            O => \N__61820\,
            I => \N__61808\
        );

    \I__14701\ : LocalMux
    port map (
            O => \N__61817\,
            I => \N__61808\
        );

    \I__14700\ : InMux
    port map (
            O => \N__61814\,
            I => \N__61804\
        );

    \I__14699\ : InMux
    port map (
            O => \N__61813\,
            I => \N__61801\
        );

    \I__14698\ : Span4Mux_h
    port map (
            O => \N__61808\,
            I => \N__61798\
        );

    \I__14697\ : InMux
    port map (
            O => \N__61807\,
            I => \N__61795\
        );

    \I__14696\ : LocalMux
    port map (
            O => \N__61804\,
            I => \c0.data_in_frame_17_6\
        );

    \I__14695\ : LocalMux
    port map (
            O => \N__61801\,
            I => \c0.data_in_frame_17_6\
        );

    \I__14694\ : Odrv4
    port map (
            O => \N__61798\,
            I => \c0.data_in_frame_17_6\
        );

    \I__14693\ : LocalMux
    port map (
            O => \N__61795\,
            I => \c0.data_in_frame_17_6\
        );

    \I__14692\ : InMux
    port map (
            O => \N__61786\,
            I => \N__61783\
        );

    \I__14691\ : LocalMux
    port map (
            O => \N__61783\,
            I => \N__61780\
        );

    \I__14690\ : Span4Mux_v
    port map (
            O => \N__61780\,
            I => \N__61777\
        );

    \I__14689\ : Odrv4
    port map (
            O => \N__61777\,
            I => \c0.n20_adj_4247\
        );

    \I__14688\ : InMux
    port map (
            O => \N__61774\,
            I => \N__61770\
        );

    \I__14687\ : CascadeMux
    port map (
            O => \N__61773\,
            I => \N__61767\
        );

    \I__14686\ : LocalMux
    port map (
            O => \N__61770\,
            I => \N__61764\
        );

    \I__14685\ : InMux
    port map (
            O => \N__61767\,
            I => \N__61760\
        );

    \I__14684\ : Span4Mux_h
    port map (
            O => \N__61764\,
            I => \N__61757\
        );

    \I__14683\ : InMux
    port map (
            O => \N__61763\,
            I => \N__61754\
        );

    \I__14682\ : LocalMux
    port map (
            O => \N__61760\,
            I => \c0.data_in_frame_20_2\
        );

    \I__14681\ : Odrv4
    port map (
            O => \N__61757\,
            I => \c0.data_in_frame_20_2\
        );

    \I__14680\ : LocalMux
    port map (
            O => \N__61754\,
            I => \c0.data_in_frame_20_2\
        );

    \I__14679\ : InMux
    port map (
            O => \N__61747\,
            I => \N__61742\
        );

    \I__14678\ : InMux
    port map (
            O => \N__61746\,
            I => \N__61738\
        );

    \I__14677\ : InMux
    port map (
            O => \N__61745\,
            I => \N__61734\
        );

    \I__14676\ : LocalMux
    port map (
            O => \N__61742\,
            I => \N__61731\
        );

    \I__14675\ : InMux
    port map (
            O => \N__61741\,
            I => \N__61728\
        );

    \I__14674\ : LocalMux
    port map (
            O => \N__61738\,
            I => \N__61725\
        );

    \I__14673\ : InMux
    port map (
            O => \N__61737\,
            I => \N__61722\
        );

    \I__14672\ : LocalMux
    port map (
            O => \N__61734\,
            I => \N__61715\
        );

    \I__14671\ : Span4Mux_h
    port map (
            O => \N__61731\,
            I => \N__61715\
        );

    \I__14670\ : LocalMux
    port map (
            O => \N__61728\,
            I => \N__61715\
        );

    \I__14669\ : Odrv4
    port map (
            O => \N__61725\,
            I => \c0.n13544\
        );

    \I__14668\ : LocalMux
    port map (
            O => \N__61722\,
            I => \c0.n13544\
        );

    \I__14667\ : Odrv4
    port map (
            O => \N__61715\,
            I => \c0.n13544\
        );

    \I__14666\ : CascadeMux
    port map (
            O => \N__61708\,
            I => \N__61705\
        );

    \I__14665\ : InMux
    port map (
            O => \N__61705\,
            I => \N__61702\
        );

    \I__14664\ : LocalMux
    port map (
            O => \N__61702\,
            I => \N__61699\
        );

    \I__14663\ : Span4Mux_v
    port map (
            O => \N__61699\,
            I => \N__61696\
        );

    \I__14662\ : Span4Mux_v
    port map (
            O => \N__61696\,
            I => \N__61691\
        );

    \I__14661\ : InMux
    port map (
            O => \N__61695\,
            I => \N__61688\
        );

    \I__14660\ : InMux
    port map (
            O => \N__61694\,
            I => \N__61685\
        );

    \I__14659\ : Span4Mux_h
    port map (
            O => \N__61691\,
            I => \N__61682\
        );

    \I__14658\ : LocalMux
    port map (
            O => \N__61688\,
            I => \N__61679\
        );

    \I__14657\ : LocalMux
    port map (
            O => \N__61685\,
            I => data_in_frame_22_3
        );

    \I__14656\ : Odrv4
    port map (
            O => \N__61682\,
            I => data_in_frame_22_3
        );

    \I__14655\ : Odrv4
    port map (
            O => \N__61679\,
            I => data_in_frame_22_3
        );

    \I__14654\ : InMux
    port map (
            O => \N__61672\,
            I => \N__61669\
        );

    \I__14653\ : LocalMux
    port map (
            O => \N__61669\,
            I => \N__61663\
        );

    \I__14652\ : InMux
    port map (
            O => \N__61668\,
            I => \N__61660\
        );

    \I__14651\ : InMux
    port map (
            O => \N__61667\,
            I => \N__61655\
        );

    \I__14650\ : InMux
    port map (
            O => \N__61666\,
            I => \N__61655\
        );

    \I__14649\ : Span4Mux_v
    port map (
            O => \N__61663\,
            I => \N__61652\
        );

    \I__14648\ : LocalMux
    port map (
            O => \N__61660\,
            I => \N__61647\
        );

    \I__14647\ : LocalMux
    port map (
            O => \N__61655\,
            I => \N__61647\
        );

    \I__14646\ : Odrv4
    port map (
            O => \N__61652\,
            I => \c0.n23426\
        );

    \I__14645\ : Odrv12
    port map (
            O => \N__61647\,
            I => \c0.n23426\
        );

    \I__14644\ : InMux
    port map (
            O => \N__61642\,
            I => \N__61638\
        );

    \I__14643\ : InMux
    port map (
            O => \N__61641\,
            I => \N__61635\
        );

    \I__14642\ : LocalMux
    port map (
            O => \N__61638\,
            I => \N__61632\
        );

    \I__14641\ : LocalMux
    port map (
            O => \N__61635\,
            I => \N__61629\
        );

    \I__14640\ : Span4Mux_v
    port map (
            O => \N__61632\,
            I => \N__61626\
        );

    \I__14639\ : Span4Mux_v
    port map (
            O => \N__61629\,
            I => \N__61623\
        );

    \I__14638\ : Odrv4
    port map (
            O => \N__61626\,
            I => \c0.n22007\
        );

    \I__14637\ : Odrv4
    port map (
            O => \N__61623\,
            I => \c0.n22007\
        );

    \I__14636\ : InMux
    port map (
            O => \N__61618\,
            I => \N__61612\
        );

    \I__14635\ : CascadeMux
    port map (
            O => \N__61617\,
            I => \N__61609\
        );

    \I__14634\ : InMux
    port map (
            O => \N__61616\,
            I => \N__61604\
        );

    \I__14633\ : InMux
    port map (
            O => \N__61615\,
            I => \N__61604\
        );

    \I__14632\ : LocalMux
    port map (
            O => \N__61612\,
            I => \N__61600\
        );

    \I__14631\ : InMux
    port map (
            O => \N__61609\,
            I => \N__61597\
        );

    \I__14630\ : LocalMux
    port map (
            O => \N__61604\,
            I => \N__61594\
        );

    \I__14629\ : InMux
    port map (
            O => \N__61603\,
            I => \N__61591\
        );

    \I__14628\ : Span4Mux_h
    port map (
            O => \N__61600\,
            I => \N__61588\
        );

    \I__14627\ : LocalMux
    port map (
            O => \N__61597\,
            I => \c0.data_in_frame_19_6\
        );

    \I__14626\ : Odrv12
    port map (
            O => \N__61594\,
            I => \c0.data_in_frame_19_6\
        );

    \I__14625\ : LocalMux
    port map (
            O => \N__61591\,
            I => \c0.data_in_frame_19_6\
        );

    \I__14624\ : Odrv4
    port map (
            O => \N__61588\,
            I => \c0.data_in_frame_19_6\
        );

    \I__14623\ : CascadeMux
    port map (
            O => \N__61579\,
            I => \N__61575\
        );

    \I__14622\ : InMux
    port map (
            O => \N__61578\,
            I => \N__61572\
        );

    \I__14621\ : InMux
    port map (
            O => \N__61575\,
            I => \N__61569\
        );

    \I__14620\ : LocalMux
    port map (
            O => \N__61572\,
            I => \N__61566\
        );

    \I__14619\ : LocalMux
    port map (
            O => \N__61569\,
            I => \c0.data_in_frame_18_5\
        );

    \I__14618\ : Odrv12
    port map (
            O => \N__61566\,
            I => \c0.data_in_frame_18_5\
        );

    \I__14617\ : InMux
    port map (
            O => \N__61561\,
            I => \N__61558\
        );

    \I__14616\ : LocalMux
    port map (
            O => \N__61558\,
            I => \N__61555\
        );

    \I__14615\ : Span4Mux_h
    port map (
            O => \N__61555\,
            I => \N__61552\
        );

    \I__14614\ : Span4Mux_v
    port map (
            O => \N__61552\,
            I => \N__61549\
        );

    \I__14613\ : Odrv4
    port map (
            O => \N__61549\,
            I => \c0.n22385\
        );

    \I__14612\ : InMux
    port map (
            O => \N__61546\,
            I => \N__61543\
        );

    \I__14611\ : LocalMux
    port map (
            O => \N__61543\,
            I => \N__61539\
        );

    \I__14610\ : InMux
    port map (
            O => \N__61542\,
            I => \N__61536\
        );

    \I__14609\ : Span12Mux_v
    port map (
            O => \N__61539\,
            I => \N__61533\
        );

    \I__14608\ : LocalMux
    port map (
            O => \N__61536\,
            I => \N__61530\
        );

    \I__14607\ : Odrv12
    port map (
            O => \N__61533\,
            I => \c0.n21126\
        );

    \I__14606\ : Odrv12
    port map (
            O => \N__61530\,
            I => \c0.n21126\
        );

    \I__14605\ : CascadeMux
    port map (
            O => \N__61525\,
            I => \N__61522\
        );

    \I__14604\ : InMux
    port map (
            O => \N__61522\,
            I => \N__61519\
        );

    \I__14603\ : LocalMux
    port map (
            O => \N__61519\,
            I => \N__61514\
        );

    \I__14602\ : InMux
    port map (
            O => \N__61518\,
            I => \N__61511\
        );

    \I__14601\ : InMux
    port map (
            O => \N__61517\,
            I => \N__61508\
        );

    \I__14600\ : Odrv4
    port map (
            O => \N__61514\,
            I => \c0.data_in_frame_16_1\
        );

    \I__14599\ : LocalMux
    port map (
            O => \N__61511\,
            I => \c0.data_in_frame_16_1\
        );

    \I__14598\ : LocalMux
    port map (
            O => \N__61508\,
            I => \c0.data_in_frame_16_1\
        );

    \I__14597\ : CascadeMux
    port map (
            O => \N__61501\,
            I => \N__61497\
        );

    \I__14596\ : CascadeMux
    port map (
            O => \N__61500\,
            I => \N__61493\
        );

    \I__14595\ : InMux
    port map (
            O => \N__61497\,
            I => \N__61488\
        );

    \I__14594\ : InMux
    port map (
            O => \N__61496\,
            I => \N__61488\
        );

    \I__14593\ : InMux
    port map (
            O => \N__61493\,
            I => \N__61485\
        );

    \I__14592\ : LocalMux
    port map (
            O => \N__61488\,
            I => \N__61482\
        );

    \I__14591\ : LocalMux
    port map (
            O => \N__61485\,
            I => \N__61476\
        );

    \I__14590\ : Span4Mux_v
    port map (
            O => \N__61482\,
            I => \N__61476\
        );

    \I__14589\ : InMux
    port map (
            O => \N__61481\,
            I => \N__61473\
        );

    \I__14588\ : Odrv4
    port map (
            O => \N__61476\,
            I => \c0.data_in_frame_12_3\
        );

    \I__14587\ : LocalMux
    port map (
            O => \N__61473\,
            I => \c0.data_in_frame_12_3\
        );

    \I__14586\ : InMux
    port map (
            O => \N__61468\,
            I => \N__61464\
        );

    \I__14585\ : InMux
    port map (
            O => \N__61467\,
            I => \N__61461\
        );

    \I__14584\ : LocalMux
    port map (
            O => \N__61464\,
            I => \N__61458\
        );

    \I__14583\ : LocalMux
    port map (
            O => \N__61461\,
            I => \N__61455\
        );

    \I__14582\ : Span4Mux_v
    port map (
            O => \N__61458\,
            I => \N__61452\
        );

    \I__14581\ : Span4Mux_h
    port map (
            O => \N__61455\,
            I => \N__61449\
        );

    \I__14580\ : Span4Mux_h
    port map (
            O => \N__61452\,
            I => \N__61443\
        );

    \I__14579\ : Span4Mux_v
    port map (
            O => \N__61449\,
            I => \N__61443\
        );

    \I__14578\ : InMux
    port map (
            O => \N__61448\,
            I => \N__61440\
        );

    \I__14577\ : Odrv4
    port map (
            O => \N__61443\,
            I => \c0.n21975\
        );

    \I__14576\ : LocalMux
    port map (
            O => \N__61440\,
            I => \c0.n21975\
        );

    \I__14575\ : InMux
    port map (
            O => \N__61435\,
            I => \N__61431\
        );

    \I__14574\ : InMux
    port map (
            O => \N__61434\,
            I => \N__61427\
        );

    \I__14573\ : LocalMux
    port map (
            O => \N__61431\,
            I => \N__61424\
        );

    \I__14572\ : InMux
    port map (
            O => \N__61430\,
            I => \N__61421\
        );

    \I__14571\ : LocalMux
    port map (
            O => \N__61427\,
            I => \N__61417\
        );

    \I__14570\ : Span4Mux_v
    port map (
            O => \N__61424\,
            I => \N__61410\
        );

    \I__14569\ : LocalMux
    port map (
            O => \N__61421\,
            I => \N__61410\
        );

    \I__14568\ : InMux
    port map (
            O => \N__61420\,
            I => \N__61407\
        );

    \I__14567\ : Span4Mux_h
    port map (
            O => \N__61417\,
            I => \N__61404\
        );

    \I__14566\ : InMux
    port map (
            O => \N__61416\,
            I => \N__61399\
        );

    \I__14565\ : InMux
    port map (
            O => \N__61415\,
            I => \N__61399\
        );

    \I__14564\ : Odrv4
    port map (
            O => \N__61410\,
            I => \c0.data_in_frame_17_2\
        );

    \I__14563\ : LocalMux
    port map (
            O => \N__61407\,
            I => \c0.data_in_frame_17_2\
        );

    \I__14562\ : Odrv4
    port map (
            O => \N__61404\,
            I => \c0.data_in_frame_17_2\
        );

    \I__14561\ : LocalMux
    port map (
            O => \N__61399\,
            I => \c0.data_in_frame_17_2\
        );

    \I__14560\ : InMux
    port map (
            O => \N__61390\,
            I => \N__61386\
        );

    \I__14559\ : InMux
    port map (
            O => \N__61389\,
            I => \N__61383\
        );

    \I__14558\ : LocalMux
    port map (
            O => \N__61386\,
            I => \N__61379\
        );

    \I__14557\ : LocalMux
    port map (
            O => \N__61383\,
            I => \N__61376\
        );

    \I__14556\ : InMux
    port map (
            O => \N__61382\,
            I => \N__61373\
        );

    \I__14555\ : Span4Mux_h
    port map (
            O => \N__61379\,
            I => \N__61370\
        );

    \I__14554\ : Span12Mux_v
    port map (
            O => \N__61376\,
            I => \N__61367\
        );

    \I__14553\ : LocalMux
    port map (
            O => \N__61373\,
            I => \c0.data_in_frame_15_1\
        );

    \I__14552\ : Odrv4
    port map (
            O => \N__61370\,
            I => \c0.data_in_frame_15_1\
        );

    \I__14551\ : Odrv12
    port map (
            O => \N__61367\,
            I => \c0.data_in_frame_15_1\
        );

    \I__14550\ : CascadeMux
    port map (
            O => \N__61360\,
            I => \N__61356\
        );

    \I__14549\ : CascadeMux
    port map (
            O => \N__61359\,
            I => \N__61353\
        );

    \I__14548\ : InMux
    port map (
            O => \N__61356\,
            I => \N__61350\
        );

    \I__14547\ : InMux
    port map (
            O => \N__61353\,
            I => \N__61347\
        );

    \I__14546\ : LocalMux
    port map (
            O => \N__61350\,
            I => \N__61344\
        );

    \I__14545\ : LocalMux
    port map (
            O => \N__61347\,
            I => \N__61338\
        );

    \I__14544\ : Span4Mux_h
    port map (
            O => \N__61344\,
            I => \N__61338\
        );

    \I__14543\ : InMux
    port map (
            O => \N__61343\,
            I => \N__61335\
        );

    \I__14542\ : Odrv4
    port map (
            O => \N__61338\,
            I => \c0.data_in_frame_12_4\
        );

    \I__14541\ : LocalMux
    port map (
            O => \N__61335\,
            I => \c0.data_in_frame_12_4\
        );

    \I__14540\ : CascadeMux
    port map (
            O => \N__61330\,
            I => \N__61326\
        );

    \I__14539\ : InMux
    port map (
            O => \N__61329\,
            I => \N__61323\
        );

    \I__14538\ : InMux
    port map (
            O => \N__61326\,
            I => \N__61319\
        );

    \I__14537\ : LocalMux
    port map (
            O => \N__61323\,
            I => \N__61316\
        );

    \I__14536\ : InMux
    port map (
            O => \N__61322\,
            I => \N__61313\
        );

    \I__14535\ : LocalMux
    port map (
            O => \N__61319\,
            I => \N__61307\
        );

    \I__14534\ : Span4Mux_v
    port map (
            O => \N__61316\,
            I => \N__61307\
        );

    \I__14533\ : LocalMux
    port map (
            O => \N__61313\,
            I => \N__61304\
        );

    \I__14532\ : InMux
    port map (
            O => \N__61312\,
            I => \N__61301\
        );

    \I__14531\ : Odrv4
    port map (
            O => \N__61307\,
            I => \c0.data_in_frame_13_3\
        );

    \I__14530\ : Odrv4
    port map (
            O => \N__61304\,
            I => \c0.data_in_frame_13_3\
        );

    \I__14529\ : LocalMux
    port map (
            O => \N__61301\,
            I => \c0.data_in_frame_13_3\
        );

    \I__14528\ : InMux
    port map (
            O => \N__61294\,
            I => \N__61291\
        );

    \I__14527\ : LocalMux
    port map (
            O => \N__61291\,
            I => \N__61286\
        );

    \I__14526\ : CascadeMux
    port map (
            O => \N__61290\,
            I => \N__61281\
        );

    \I__14525\ : InMux
    port map (
            O => \N__61289\,
            I => \N__61278\
        );

    \I__14524\ : Span4Mux_h
    port map (
            O => \N__61286\,
            I => \N__61275\
        );

    \I__14523\ : InMux
    port map (
            O => \N__61285\,
            I => \N__61268\
        );

    \I__14522\ : InMux
    port map (
            O => \N__61284\,
            I => \N__61268\
        );

    \I__14521\ : InMux
    port map (
            O => \N__61281\,
            I => \N__61268\
        );

    \I__14520\ : LocalMux
    port map (
            O => \N__61278\,
            I => \c0.data_in_frame_13_5\
        );

    \I__14519\ : Odrv4
    port map (
            O => \N__61275\,
            I => \c0.data_in_frame_13_5\
        );

    \I__14518\ : LocalMux
    port map (
            O => \N__61268\,
            I => \c0.data_in_frame_13_5\
        );

    \I__14517\ : CascadeMux
    port map (
            O => \N__61261\,
            I => \N__61258\
        );

    \I__14516\ : InMux
    port map (
            O => \N__61258\,
            I => \N__61255\
        );

    \I__14515\ : LocalMux
    port map (
            O => \N__61255\,
            I => \N__61251\
        );

    \I__14514\ : InMux
    port map (
            O => \N__61254\,
            I => \N__61248\
        );

    \I__14513\ : Odrv12
    port map (
            O => \N__61251\,
            I => \c0.n14081\
        );

    \I__14512\ : LocalMux
    port map (
            O => \N__61248\,
            I => \c0.n14081\
        );

    \I__14511\ : CascadeMux
    port map (
            O => \N__61243\,
            I => \N__61239\
        );

    \I__14510\ : InMux
    port map (
            O => \N__61242\,
            I => \N__61236\
        );

    \I__14509\ : InMux
    port map (
            O => \N__61239\,
            I => \N__61232\
        );

    \I__14508\ : LocalMux
    port map (
            O => \N__61236\,
            I => \N__61229\
        );

    \I__14507\ : InMux
    port map (
            O => \N__61235\,
            I => \N__61226\
        );

    \I__14506\ : LocalMux
    port map (
            O => \N__61232\,
            I => \N__61219\
        );

    \I__14505\ : Span4Mux_h
    port map (
            O => \N__61229\,
            I => \N__61219\
        );

    \I__14504\ : LocalMux
    port map (
            O => \N__61226\,
            I => \N__61219\
        );

    \I__14503\ : Odrv4
    port map (
            O => \N__61219\,
            I => \c0.data_in_frame_16_0\
        );

    \I__14502\ : CascadeMux
    port map (
            O => \N__61216\,
            I => \N__61213\
        );

    \I__14501\ : InMux
    port map (
            O => \N__61213\,
            I => \N__61210\
        );

    \I__14500\ : LocalMux
    port map (
            O => \N__61210\,
            I => \N__61206\
        );

    \I__14499\ : CascadeMux
    port map (
            O => \N__61209\,
            I => \N__61203\
        );

    \I__14498\ : Span4Mux_v
    port map (
            O => \N__61206\,
            I => \N__61199\
        );

    \I__14497\ : InMux
    port map (
            O => \N__61203\,
            I => \N__61196\
        );

    \I__14496\ : CascadeMux
    port map (
            O => \N__61202\,
            I => \N__61193\
        );

    \I__14495\ : Span4Mux_h
    port map (
            O => \N__61199\,
            I => \N__61188\
        );

    \I__14494\ : LocalMux
    port map (
            O => \N__61196\,
            I => \N__61188\
        );

    \I__14493\ : InMux
    port map (
            O => \N__61193\,
            I => \N__61185\
        );

    \I__14492\ : Span4Mux_v
    port map (
            O => \N__61188\,
            I => \N__61182\
        );

    \I__14491\ : LocalMux
    port map (
            O => \N__61185\,
            I => \c0.data_in_frame_21_7\
        );

    \I__14490\ : Odrv4
    port map (
            O => \N__61182\,
            I => \c0.data_in_frame_21_7\
        );

    \I__14489\ : InMux
    port map (
            O => \N__61177\,
            I => \N__61173\
        );

    \I__14488\ : InMux
    port map (
            O => \N__61176\,
            I => \N__61169\
        );

    \I__14487\ : LocalMux
    port map (
            O => \N__61173\,
            I => \N__61166\
        );

    \I__14486\ : InMux
    port map (
            O => \N__61172\,
            I => \N__61163\
        );

    \I__14485\ : LocalMux
    port map (
            O => \N__61169\,
            I => \c0.n13210\
        );

    \I__14484\ : Odrv4
    port map (
            O => \N__61166\,
            I => \c0.n13210\
        );

    \I__14483\ : LocalMux
    port map (
            O => \N__61163\,
            I => \c0.n13210\
        );

    \I__14482\ : InMux
    port map (
            O => \N__61156\,
            I => \N__61153\
        );

    \I__14481\ : LocalMux
    port map (
            O => \N__61153\,
            I => \N__61150\
        );

    \I__14480\ : Span4Mux_h
    port map (
            O => \N__61150\,
            I => \N__61146\
        );

    \I__14479\ : InMux
    port map (
            O => \N__61149\,
            I => \N__61143\
        );

    \I__14478\ : Odrv4
    port map (
            O => \N__61146\,
            I => \c0.n22091\
        );

    \I__14477\ : LocalMux
    port map (
            O => \N__61143\,
            I => \c0.n22091\
        );

    \I__14476\ : InMux
    port map (
            O => \N__61138\,
            I => \N__61135\
        );

    \I__14475\ : LocalMux
    port map (
            O => \N__61135\,
            I => \N__61132\
        );

    \I__14474\ : Span4Mux_v
    port map (
            O => \N__61132\,
            I => \N__61128\
        );

    \I__14473\ : InMux
    port map (
            O => \N__61131\,
            I => \N__61125\
        );

    \I__14472\ : Sp12to4
    port map (
            O => \N__61128\,
            I => \N__61119\
        );

    \I__14471\ : LocalMux
    port map (
            O => \N__61125\,
            I => \N__61119\
        );

    \I__14470\ : InMux
    port map (
            O => \N__61124\,
            I => \N__61116\
        );

    \I__14469\ : Odrv12
    port map (
            O => \N__61119\,
            I => \c0.n21934\
        );

    \I__14468\ : LocalMux
    port map (
            O => \N__61116\,
            I => \c0.n21934\
        );

    \I__14467\ : InMux
    port map (
            O => \N__61111\,
            I => \N__61108\
        );

    \I__14466\ : LocalMux
    port map (
            O => \N__61108\,
            I => \N__61104\
        );

    \I__14465\ : InMux
    port map (
            O => \N__61107\,
            I => \N__61100\
        );

    \I__14464\ : Span4Mux_h
    port map (
            O => \N__61104\,
            I => \N__61097\
        );

    \I__14463\ : InMux
    port map (
            O => \N__61103\,
            I => \N__61094\
        );

    \I__14462\ : LocalMux
    port map (
            O => \N__61100\,
            I => \N__61089\
        );

    \I__14461\ : Span4Mux_h
    port map (
            O => \N__61097\,
            I => \N__61084\
        );

    \I__14460\ : LocalMux
    port map (
            O => \N__61094\,
            I => \N__61084\
        );

    \I__14459\ : InMux
    port map (
            O => \N__61093\,
            I => \N__61079\
        );

    \I__14458\ : InMux
    port map (
            O => \N__61092\,
            I => \N__61079\
        );

    \I__14457\ : Odrv12
    port map (
            O => \N__61089\,
            I => \c0.data_in_frame_4_5\
        );

    \I__14456\ : Odrv4
    port map (
            O => \N__61084\,
            I => \c0.data_in_frame_4_5\
        );

    \I__14455\ : LocalMux
    port map (
            O => \N__61079\,
            I => \c0.data_in_frame_4_5\
        );

    \I__14454\ : CascadeMux
    port map (
            O => \N__61072\,
            I => \N__61069\
        );

    \I__14453\ : InMux
    port map (
            O => \N__61069\,
            I => \N__61066\
        );

    \I__14452\ : LocalMux
    port map (
            O => \N__61066\,
            I => \N__61063\
        );

    \I__14451\ : Span4Mux_v
    port map (
            O => \N__61063\,
            I => \N__61059\
        );

    \I__14450\ : InMux
    port map (
            O => \N__61062\,
            I => \N__61056\
        );

    \I__14449\ : Span4Mux_h
    port map (
            O => \N__61059\,
            I => \N__61051\
        );

    \I__14448\ : LocalMux
    port map (
            O => \N__61056\,
            I => \N__61051\
        );

    \I__14447\ : Span4Mux_h
    port map (
            O => \N__61051\,
            I => \N__61048\
        );

    \I__14446\ : Odrv4
    port map (
            O => \N__61048\,
            I => \c0.n13421\
        );

    \I__14445\ : CascadeMux
    port map (
            O => \N__61045\,
            I => \N__61041\
        );

    \I__14444\ : InMux
    port map (
            O => \N__61044\,
            I => \N__61037\
        );

    \I__14443\ : InMux
    port map (
            O => \N__61041\,
            I => \N__61032\
        );

    \I__14442\ : InMux
    port map (
            O => \N__61040\,
            I => \N__61032\
        );

    \I__14441\ : LocalMux
    port map (
            O => \N__61037\,
            I => \c0.data_in_frame_11_4\
        );

    \I__14440\ : LocalMux
    port map (
            O => \N__61032\,
            I => \c0.data_in_frame_11_4\
        );

    \I__14439\ : CascadeMux
    port map (
            O => \N__61027\,
            I => \c0.n13421_cascade_\
        );

    \I__14438\ : InMux
    port map (
            O => \N__61024\,
            I => \N__61020\
        );

    \I__14437\ : InMux
    port map (
            O => \N__61023\,
            I => \N__61017\
        );

    \I__14436\ : LocalMux
    port map (
            O => \N__61020\,
            I => \N__61014\
        );

    \I__14435\ : LocalMux
    port map (
            O => \N__61017\,
            I => \N__61011\
        );

    \I__14434\ : Span4Mux_h
    port map (
            O => \N__61014\,
            I => \N__61008\
        );

    \I__14433\ : Odrv12
    port map (
            O => \N__61011\,
            I => \c0.n22069\
        );

    \I__14432\ : Odrv4
    port map (
            O => \N__61008\,
            I => \c0.n22069\
        );

    \I__14431\ : InMux
    port map (
            O => \N__61003\,
            I => \N__61000\
        );

    \I__14430\ : LocalMux
    port map (
            O => \N__61000\,
            I => \c0.n10_adj_4252\
        );

    \I__14429\ : CascadeMux
    port map (
            O => \N__60997\,
            I => \N__60993\
        );

    \I__14428\ : InMux
    port map (
            O => \N__60996\,
            I => \N__60990\
        );

    \I__14427\ : InMux
    port map (
            O => \N__60993\,
            I => \N__60986\
        );

    \I__14426\ : LocalMux
    port map (
            O => \N__60990\,
            I => \N__60983\
        );

    \I__14425\ : InMux
    port map (
            O => \N__60989\,
            I => \N__60980\
        );

    \I__14424\ : LocalMux
    port map (
            O => \N__60986\,
            I => \c0.data_in_frame_7_2\
        );

    \I__14423\ : Odrv4
    port map (
            O => \N__60983\,
            I => \c0.data_in_frame_7_2\
        );

    \I__14422\ : LocalMux
    port map (
            O => \N__60980\,
            I => \c0.data_in_frame_7_2\
        );

    \I__14421\ : InMux
    port map (
            O => \N__60973\,
            I => \N__60969\
        );

    \I__14420\ : InMux
    port map (
            O => \N__60972\,
            I => \N__60966\
        );

    \I__14419\ : LocalMux
    port map (
            O => \N__60969\,
            I => \N__60963\
        );

    \I__14418\ : LocalMux
    port map (
            O => \N__60966\,
            I => \c0.n22343\
        );

    \I__14417\ : Odrv12
    port map (
            O => \N__60963\,
            I => \c0.n22343\
        );

    \I__14416\ : InMux
    port map (
            O => \N__60958\,
            I => \N__60955\
        );

    \I__14415\ : LocalMux
    port map (
            O => \N__60955\,
            I => \N__60952\
        );

    \I__14414\ : Odrv4
    port map (
            O => \N__60952\,
            I => \c0.n10_adj_4267\
        );

    \I__14413\ : CascadeMux
    port map (
            O => \N__60949\,
            I => \N__60944\
        );

    \I__14412\ : CascadeMux
    port map (
            O => \N__60948\,
            I => \N__60941\
        );

    \I__14411\ : InMux
    port map (
            O => \N__60947\,
            I => \N__60938\
        );

    \I__14410\ : InMux
    port map (
            O => \N__60944\,
            I => \N__60934\
        );

    \I__14409\ : InMux
    port map (
            O => \N__60941\,
            I => \N__60931\
        );

    \I__14408\ : LocalMux
    port map (
            O => \N__60938\,
            I => \N__60928\
        );

    \I__14407\ : InMux
    port map (
            O => \N__60937\,
            I => \N__60925\
        );

    \I__14406\ : LocalMux
    port map (
            O => \N__60934\,
            I => \N__60922\
        );

    \I__14405\ : LocalMux
    port map (
            O => \N__60931\,
            I => \N__60915\
        );

    \I__14404\ : Span4Mux_v
    port map (
            O => \N__60928\,
            I => \N__60915\
        );

    \I__14403\ : LocalMux
    port map (
            O => \N__60925\,
            I => \N__60915\
        );

    \I__14402\ : Span4Mux_h
    port map (
            O => \N__60922\,
            I => \N__60912\
        );

    \I__14401\ : Odrv4
    port map (
            O => \N__60915\,
            I => \c0.data_in_frame_12_5\
        );

    \I__14400\ : Odrv4
    port map (
            O => \N__60912\,
            I => \c0.data_in_frame_12_5\
        );

    \I__14399\ : InMux
    port map (
            O => \N__60907\,
            I => \N__60904\
        );

    \I__14398\ : LocalMux
    port map (
            O => \N__60904\,
            I => \N__60901\
        );

    \I__14397\ : Odrv4
    port map (
            O => \N__60901\,
            I => \c0.n16_adj_4268\
        );

    \I__14396\ : InMux
    port map (
            O => \N__60898\,
            I => \N__60884\
        );

    \I__14395\ : InMux
    port map (
            O => \N__60897\,
            I => \N__60878\
        );

    \I__14394\ : InMux
    port map (
            O => \N__60896\,
            I => \N__60871\
        );

    \I__14393\ : InMux
    port map (
            O => \N__60895\,
            I => \N__60871\
        );

    \I__14392\ : InMux
    port map (
            O => \N__60894\,
            I => \N__60871\
        );

    \I__14391\ : CascadeMux
    port map (
            O => \N__60893\,
            I => \N__60864\
        );

    \I__14390\ : InMux
    port map (
            O => \N__60892\,
            I => \N__60856\
        );

    \I__14389\ : InMux
    port map (
            O => \N__60891\,
            I => \N__60856\
        );

    \I__14388\ : InMux
    port map (
            O => \N__60890\,
            I => \N__60856\
        );

    \I__14387\ : InMux
    port map (
            O => \N__60889\,
            I => \N__60853\
        );

    \I__14386\ : InMux
    port map (
            O => \N__60888\,
            I => \N__60839\
        );

    \I__14385\ : CascadeMux
    port map (
            O => \N__60887\,
            I => \N__60836\
        );

    \I__14384\ : LocalMux
    port map (
            O => \N__60884\,
            I => \N__60831\
        );

    \I__14383\ : InMux
    port map (
            O => \N__60883\,
            I => \N__60824\
        );

    \I__14382\ : InMux
    port map (
            O => \N__60882\,
            I => \N__60824\
        );

    \I__14381\ : InMux
    port map (
            O => \N__60881\,
            I => \N__60824\
        );

    \I__14380\ : LocalMux
    port map (
            O => \N__60878\,
            I => \N__60820\
        );

    \I__14379\ : LocalMux
    port map (
            O => \N__60871\,
            I => \N__60817\
        );

    \I__14378\ : InMux
    port map (
            O => \N__60870\,
            I => \N__60808\
        );

    \I__14377\ : InMux
    port map (
            O => \N__60869\,
            I => \N__60808\
        );

    \I__14376\ : InMux
    port map (
            O => \N__60868\,
            I => \N__60808\
        );

    \I__14375\ : InMux
    port map (
            O => \N__60867\,
            I => \N__60808\
        );

    \I__14374\ : InMux
    port map (
            O => \N__60864\,
            I => \N__60803\
        );

    \I__14373\ : InMux
    port map (
            O => \N__60863\,
            I => \N__60800\
        );

    \I__14372\ : LocalMux
    port map (
            O => \N__60856\,
            I => \N__60795\
        );

    \I__14371\ : LocalMux
    port map (
            O => \N__60853\,
            I => \N__60795\
        );

    \I__14370\ : InMux
    port map (
            O => \N__60852\,
            I => \N__60784\
        );

    \I__14369\ : InMux
    port map (
            O => \N__60851\,
            I => \N__60784\
        );

    \I__14368\ : InMux
    port map (
            O => \N__60850\,
            I => \N__60784\
        );

    \I__14367\ : InMux
    port map (
            O => \N__60849\,
            I => \N__60784\
        );

    \I__14366\ : InMux
    port map (
            O => \N__60848\,
            I => \N__60784\
        );

    \I__14365\ : InMux
    port map (
            O => \N__60847\,
            I => \N__60777\
        );

    \I__14364\ : InMux
    port map (
            O => \N__60846\,
            I => \N__60777\
        );

    \I__14363\ : InMux
    port map (
            O => \N__60845\,
            I => \N__60777\
        );

    \I__14362\ : InMux
    port map (
            O => \N__60844\,
            I => \N__60770\
        );

    \I__14361\ : InMux
    port map (
            O => \N__60843\,
            I => \N__60770\
        );

    \I__14360\ : InMux
    port map (
            O => \N__60842\,
            I => \N__60770\
        );

    \I__14359\ : LocalMux
    port map (
            O => \N__60839\,
            I => \N__60767\
        );

    \I__14358\ : InMux
    port map (
            O => \N__60836\,
            I => \N__60752\
        );

    \I__14357\ : InMux
    port map (
            O => \N__60835\,
            I => \N__60747\
        );

    \I__14356\ : InMux
    port map (
            O => \N__60834\,
            I => \N__60747\
        );

    \I__14355\ : Span4Mux_h
    port map (
            O => \N__60831\,
            I => \N__60742\
        );

    \I__14354\ : LocalMux
    port map (
            O => \N__60824\,
            I => \N__60742\
        );

    \I__14353\ : InMux
    port map (
            O => \N__60823\,
            I => \N__60739\
        );

    \I__14352\ : Span4Mux_h
    port map (
            O => \N__60820\,
            I => \N__60734\
        );

    \I__14351\ : Span4Mux_v
    port map (
            O => \N__60817\,
            I => \N__60734\
        );

    \I__14350\ : LocalMux
    port map (
            O => \N__60808\,
            I => \N__60731\
        );

    \I__14349\ : InMux
    port map (
            O => \N__60807\,
            I => \N__60728\
        );

    \I__14348\ : InMux
    port map (
            O => \N__60806\,
            I => \N__60724\
        );

    \I__14347\ : LocalMux
    port map (
            O => \N__60803\,
            I => \N__60719\
        );

    \I__14346\ : LocalMux
    port map (
            O => \N__60800\,
            I => \N__60719\
        );

    \I__14345\ : Span4Mux_v
    port map (
            O => \N__60795\,
            I => \N__60716\
        );

    \I__14344\ : LocalMux
    port map (
            O => \N__60784\,
            I => \N__60708\
        );

    \I__14343\ : LocalMux
    port map (
            O => \N__60777\,
            I => \N__60708\
        );

    \I__14342\ : LocalMux
    port map (
            O => \N__60770\,
            I => \N__60703\
        );

    \I__14341\ : Span4Mux_h
    port map (
            O => \N__60767\,
            I => \N__60703\
        );

    \I__14340\ : InMux
    port map (
            O => \N__60766\,
            I => \N__60688\
        );

    \I__14339\ : InMux
    port map (
            O => \N__60765\,
            I => \N__60688\
        );

    \I__14338\ : InMux
    port map (
            O => \N__60764\,
            I => \N__60688\
        );

    \I__14337\ : InMux
    port map (
            O => \N__60763\,
            I => \N__60688\
        );

    \I__14336\ : InMux
    port map (
            O => \N__60762\,
            I => \N__60688\
        );

    \I__14335\ : InMux
    port map (
            O => \N__60761\,
            I => \N__60688\
        );

    \I__14334\ : InMux
    port map (
            O => \N__60760\,
            I => \N__60688\
        );

    \I__14333\ : InMux
    port map (
            O => \N__60759\,
            I => \N__60685\
        );

    \I__14332\ : InMux
    port map (
            O => \N__60758\,
            I => \N__60676\
        );

    \I__14331\ : InMux
    port map (
            O => \N__60757\,
            I => \N__60676\
        );

    \I__14330\ : InMux
    port map (
            O => \N__60756\,
            I => \N__60676\
        );

    \I__14329\ : InMux
    port map (
            O => \N__60755\,
            I => \N__60676\
        );

    \I__14328\ : LocalMux
    port map (
            O => \N__60752\,
            I => \N__60673\
        );

    \I__14327\ : LocalMux
    port map (
            O => \N__60747\,
            I => \N__60668\
        );

    \I__14326\ : Span4Mux_h
    port map (
            O => \N__60742\,
            I => \N__60668\
        );

    \I__14325\ : LocalMux
    port map (
            O => \N__60739\,
            I => \N__60661\
        );

    \I__14324\ : Span4Mux_h
    port map (
            O => \N__60734\,
            I => \N__60661\
        );

    \I__14323\ : Span4Mux_v
    port map (
            O => \N__60731\,
            I => \N__60661\
        );

    \I__14322\ : LocalMux
    port map (
            O => \N__60728\,
            I => \N__60658\
        );

    \I__14321\ : InMux
    port map (
            O => \N__60727\,
            I => \N__60655\
        );

    \I__14320\ : LocalMux
    port map (
            O => \N__60724\,
            I => \N__60652\
        );

    \I__14319\ : Span4Mux_v
    port map (
            O => \N__60719\,
            I => \N__60649\
        );

    \I__14318\ : Span4Mux_v
    port map (
            O => \N__60716\,
            I => \N__60646\
        );

    \I__14317\ : InMux
    port map (
            O => \N__60715\,
            I => \N__60639\
        );

    \I__14316\ : InMux
    port map (
            O => \N__60714\,
            I => \N__60634\
        );

    \I__14315\ : InMux
    port map (
            O => \N__60713\,
            I => \N__60634\
        );

    \I__14314\ : Span4Mux_v
    port map (
            O => \N__60708\,
            I => \N__60629\
        );

    \I__14313\ : Span4Mux_v
    port map (
            O => \N__60703\,
            I => \N__60629\
        );

    \I__14312\ : LocalMux
    port map (
            O => \N__60688\,
            I => \N__60624\
        );

    \I__14311\ : LocalMux
    port map (
            O => \N__60685\,
            I => \N__60624\
        );

    \I__14310\ : LocalMux
    port map (
            O => \N__60676\,
            I => \N__60617\
        );

    \I__14309\ : Span4Mux_h
    port map (
            O => \N__60673\,
            I => \N__60617\
        );

    \I__14308\ : Span4Mux_v
    port map (
            O => \N__60668\,
            I => \N__60617\
        );

    \I__14307\ : Span4Mux_v
    port map (
            O => \N__60661\,
            I => \N__60614\
        );

    \I__14306\ : Span12Mux_v
    port map (
            O => \N__60658\,
            I => \N__60611\
        );

    \I__14305\ : LocalMux
    port map (
            O => \N__60655\,
            I => \N__60602\
        );

    \I__14304\ : Span4Mux_v
    port map (
            O => \N__60652\,
            I => \N__60602\
        );

    \I__14303\ : Span4Mux_h
    port map (
            O => \N__60649\,
            I => \N__60602\
        );

    \I__14302\ : Span4Mux_h
    port map (
            O => \N__60646\,
            I => \N__60602\
        );

    \I__14301\ : InMux
    port map (
            O => \N__60645\,
            I => \N__60593\
        );

    \I__14300\ : InMux
    port map (
            O => \N__60644\,
            I => \N__60593\
        );

    \I__14299\ : InMux
    port map (
            O => \N__60643\,
            I => \N__60593\
        );

    \I__14298\ : InMux
    port map (
            O => \N__60642\,
            I => \N__60593\
        );

    \I__14297\ : LocalMux
    port map (
            O => \N__60639\,
            I => \c0.n21740\
        );

    \I__14296\ : LocalMux
    port map (
            O => \N__60634\,
            I => \c0.n21740\
        );

    \I__14295\ : Odrv4
    port map (
            O => \N__60629\,
            I => \c0.n21740\
        );

    \I__14294\ : Odrv12
    port map (
            O => \N__60624\,
            I => \c0.n21740\
        );

    \I__14293\ : Odrv4
    port map (
            O => \N__60617\,
            I => \c0.n21740\
        );

    \I__14292\ : Odrv4
    port map (
            O => \N__60614\,
            I => \c0.n21740\
        );

    \I__14291\ : Odrv12
    port map (
            O => \N__60611\,
            I => \c0.n21740\
        );

    \I__14290\ : Odrv4
    port map (
            O => \N__60602\,
            I => \c0.n21740\
        );

    \I__14289\ : LocalMux
    port map (
            O => \N__60593\,
            I => \c0.n21740\
        );

    \I__14288\ : InMux
    port map (
            O => \N__60574\,
            I => \N__60571\
        );

    \I__14287\ : LocalMux
    port map (
            O => \N__60571\,
            I => \N__60568\
        );

    \I__14286\ : Span4Mux_h
    port map (
            O => \N__60568\,
            I => \N__60563\
        );

    \I__14285\ : InMux
    port map (
            O => \N__60567\,
            I => \N__60558\
        );

    \I__14284\ : InMux
    port map (
            O => \N__60566\,
            I => \N__60558\
        );

    \I__14283\ : Odrv4
    port map (
            O => \N__60563\,
            I => \c0.data_in_frame_7_0\
        );

    \I__14282\ : LocalMux
    port map (
            O => \N__60558\,
            I => \c0.data_in_frame_7_0\
        );

    \I__14281\ : InMux
    port map (
            O => \N__60553\,
            I => \N__60550\
        );

    \I__14280\ : LocalMux
    port map (
            O => \N__60550\,
            I => \N__60547\
        );

    \I__14279\ : Span4Mux_h
    port map (
            O => \N__60547\,
            I => \N__60543\
        );

    \I__14278\ : InMux
    port map (
            O => \N__60546\,
            I => \N__60540\
        );

    \I__14277\ : Odrv4
    port map (
            O => \N__60543\,
            I => \c0.n21845\
        );

    \I__14276\ : LocalMux
    port map (
            O => \N__60540\,
            I => \c0.n21845\
        );

    \I__14275\ : InMux
    port map (
            O => \N__60535\,
            I => \N__60532\
        );

    \I__14274\ : LocalMux
    port map (
            O => \N__60532\,
            I => \N__60528\
        );

    \I__14273\ : InMux
    port map (
            O => \N__60531\,
            I => \N__60525\
        );

    \I__14272\ : Odrv4
    port map (
            O => \N__60528\,
            I => \c0.n22781\
        );

    \I__14271\ : LocalMux
    port map (
            O => \N__60525\,
            I => \c0.n22781\
        );

    \I__14270\ : InMux
    port map (
            O => \N__60520\,
            I => \N__60516\
        );

    \I__14269\ : CascadeMux
    port map (
            O => \N__60519\,
            I => \N__60513\
        );

    \I__14268\ : LocalMux
    port map (
            O => \N__60516\,
            I => \N__60508\
        );

    \I__14267\ : InMux
    port map (
            O => \N__60513\,
            I => \N__60503\
        );

    \I__14266\ : InMux
    port map (
            O => \N__60512\,
            I => \N__60503\
        );

    \I__14265\ : InMux
    port map (
            O => \N__60511\,
            I => \N__60500\
        );

    \I__14264\ : Span4Mux_h
    port map (
            O => \N__60508\,
            I => \N__60497\
        );

    \I__14263\ : LocalMux
    port map (
            O => \N__60503\,
            I => \c0.data_in_frame_11_1\
        );

    \I__14262\ : LocalMux
    port map (
            O => \N__60500\,
            I => \c0.data_in_frame_11_1\
        );

    \I__14261\ : Odrv4
    port map (
            O => \N__60497\,
            I => \c0.data_in_frame_11_1\
        );

    \I__14260\ : InMux
    port map (
            O => \N__60490\,
            I => \N__60486\
        );

    \I__14259\ : InMux
    port map (
            O => \N__60489\,
            I => \N__60483\
        );

    \I__14258\ : LocalMux
    port map (
            O => \N__60486\,
            I => \N__60479\
        );

    \I__14257\ : LocalMux
    port map (
            O => \N__60483\,
            I => \N__60476\
        );

    \I__14256\ : CascadeMux
    port map (
            O => \N__60482\,
            I => \N__60473\
        );

    \I__14255\ : Span4Mux_v
    port map (
            O => \N__60479\,
            I => \N__60470\
        );

    \I__14254\ : Span4Mux_v
    port map (
            O => \N__60476\,
            I => \N__60467\
        );

    \I__14253\ : InMux
    port map (
            O => \N__60473\,
            I => \N__60464\
        );

    \I__14252\ : Span4Mux_v
    port map (
            O => \N__60470\,
            I => \N__60461\
        );

    \I__14251\ : Span4Mux_v
    port map (
            O => \N__60467\,
            I => \N__60458\
        );

    \I__14250\ : LocalMux
    port map (
            O => \N__60464\,
            I => \c0.data_in_frame_23_3\
        );

    \I__14249\ : Odrv4
    port map (
            O => \N__60461\,
            I => \c0.data_in_frame_23_3\
        );

    \I__14248\ : Odrv4
    port map (
            O => \N__60458\,
            I => \c0.data_in_frame_23_3\
        );

    \I__14247\ : InMux
    port map (
            O => \N__60451\,
            I => \N__60447\
        );

    \I__14246\ : InMux
    port map (
            O => \N__60450\,
            I => \N__60444\
        );

    \I__14245\ : LocalMux
    port map (
            O => \N__60447\,
            I => \N__60441\
        );

    \I__14244\ : LocalMux
    port map (
            O => \N__60444\,
            I => \c0.n22236\
        );

    \I__14243\ : Odrv4
    port map (
            O => \N__60441\,
            I => \c0.n22236\
        );

    \I__14242\ : InMux
    port map (
            O => \N__60436\,
            I => \N__60432\
        );

    \I__14241\ : InMux
    port map (
            O => \N__60435\,
            I => \N__60429\
        );

    \I__14240\ : LocalMux
    port map (
            O => \N__60432\,
            I => \N__60426\
        );

    \I__14239\ : LocalMux
    port map (
            O => \N__60429\,
            I => \c0.n4\
        );

    \I__14238\ : Odrv12
    port map (
            O => \N__60426\,
            I => \c0.n4\
        );

    \I__14237\ : CascadeMux
    port map (
            O => \N__60421\,
            I => \N__60418\
        );

    \I__14236\ : InMux
    port map (
            O => \N__60418\,
            I => \N__60415\
        );

    \I__14235\ : LocalMux
    port map (
            O => \N__60415\,
            I => \c0.n5965\
        );

    \I__14234\ : InMux
    port map (
            O => \N__60412\,
            I => \N__60409\
        );

    \I__14233\ : LocalMux
    port map (
            O => \N__60409\,
            I => \c0.n8_adj_4275\
        );

    \I__14232\ : InMux
    port map (
            O => \N__60406\,
            I => \N__60403\
        );

    \I__14231\ : LocalMux
    port map (
            O => \N__60403\,
            I => \c0.n8_adj_4276\
        );

    \I__14230\ : InMux
    port map (
            O => \N__60400\,
            I => \N__60395\
        );

    \I__14229\ : InMux
    port map (
            O => \N__60399\,
            I => \N__60392\
        );

    \I__14228\ : CascadeMux
    port map (
            O => \N__60398\,
            I => \N__60389\
        );

    \I__14227\ : LocalMux
    port map (
            O => \N__60395\,
            I => \N__60384\
        );

    \I__14226\ : LocalMux
    port map (
            O => \N__60392\,
            I => \N__60384\
        );

    \I__14225\ : InMux
    port map (
            O => \N__60389\,
            I => \N__60380\
        );

    \I__14224\ : Span4Mux_v
    port map (
            O => \N__60384\,
            I => \N__60377\
        );

    \I__14223\ : InMux
    port map (
            O => \N__60383\,
            I => \N__60374\
        );

    \I__14222\ : LocalMux
    port map (
            O => \N__60380\,
            I => \c0.data_in_frame_13_0\
        );

    \I__14221\ : Odrv4
    port map (
            O => \N__60377\,
            I => \c0.data_in_frame_13_0\
        );

    \I__14220\ : LocalMux
    port map (
            O => \N__60374\,
            I => \c0.data_in_frame_13_0\
        );

    \I__14219\ : InMux
    port map (
            O => \N__60367\,
            I => \N__60364\
        );

    \I__14218\ : LocalMux
    port map (
            O => \N__60364\,
            I => \N__60360\
        );

    \I__14217\ : InMux
    port map (
            O => \N__60363\,
            I => \N__60357\
        );

    \I__14216\ : Span4Mux_v
    port map (
            O => \N__60360\,
            I => \N__60351\
        );

    \I__14215\ : LocalMux
    port map (
            O => \N__60357\,
            I => \N__60351\
        );

    \I__14214\ : InMux
    port map (
            O => \N__60356\,
            I => \N__60348\
        );

    \I__14213\ : Span4Mux_h
    port map (
            O => \N__60351\,
            I => \N__60345\
        );

    \I__14212\ : LocalMux
    port map (
            O => \N__60348\,
            I => \c0.data_in_frame_12_7\
        );

    \I__14211\ : Odrv4
    port map (
            O => \N__60345\,
            I => \c0.data_in_frame_12_7\
        );

    \I__14210\ : InMux
    port map (
            O => \N__60340\,
            I => \N__60337\
        );

    \I__14209\ : LocalMux
    port map (
            O => \N__60337\,
            I => \N__60334\
        );

    \I__14208\ : Span4Mux_h
    port map (
            O => \N__60334\,
            I => \N__60330\
        );

    \I__14207\ : InMux
    port map (
            O => \N__60333\,
            I => \N__60326\
        );

    \I__14206\ : Span4Mux_v
    port map (
            O => \N__60330\,
            I => \N__60323\
        );

    \I__14205\ : InMux
    port map (
            O => \N__60329\,
            I => \N__60320\
        );

    \I__14204\ : LocalMux
    port map (
            O => \N__60326\,
            I => \c0.data_in_frame_23_1\
        );

    \I__14203\ : Odrv4
    port map (
            O => \N__60323\,
            I => \c0.data_in_frame_23_1\
        );

    \I__14202\ : LocalMux
    port map (
            O => \N__60320\,
            I => \c0.data_in_frame_23_1\
        );

    \I__14201\ : InMux
    port map (
            O => \N__60313\,
            I => \N__60305\
        );

    \I__14200\ : InMux
    port map (
            O => \N__60312\,
            I => \N__60305\
        );

    \I__14199\ : InMux
    port map (
            O => \N__60311\,
            I => \N__60302\
        );

    \I__14198\ : InMux
    port map (
            O => \N__60310\,
            I => \N__60299\
        );

    \I__14197\ : LocalMux
    port map (
            O => \N__60305\,
            I => \N__60296\
        );

    \I__14196\ : LocalMux
    port map (
            O => \N__60302\,
            I => \N__60293\
        );

    \I__14195\ : LocalMux
    port map (
            O => \N__60299\,
            I => \N__60290\
        );

    \I__14194\ : Span4Mux_v
    port map (
            O => \N__60296\,
            I => \N__60287\
        );

    \I__14193\ : Span4Mux_h
    port map (
            O => \N__60293\,
            I => \N__60284\
        );

    \I__14192\ : Odrv4
    port map (
            O => \N__60290\,
            I => data_in_frame_22_7
        );

    \I__14191\ : Odrv4
    port map (
            O => \N__60287\,
            I => data_in_frame_22_7
        );

    \I__14190\ : Odrv4
    port map (
            O => \N__60284\,
            I => data_in_frame_22_7
        );

    \I__14189\ : CascadeMux
    port map (
            O => \N__60277\,
            I => \N__60274\
        );

    \I__14188\ : InMux
    port map (
            O => \N__60274\,
            I => \N__60271\
        );

    \I__14187\ : LocalMux
    port map (
            O => \N__60271\,
            I => \N__60268\
        );

    \I__14186\ : Span4Mux_h
    port map (
            O => \N__60268\,
            I => \N__60265\
        );

    \I__14185\ : Span4Mux_v
    port map (
            O => \N__60265\,
            I => \N__60262\
        );

    \I__14184\ : Odrv4
    port map (
            O => \N__60262\,
            I => \c0.n21995\
        );

    \I__14183\ : CascadeMux
    port map (
            O => \N__60259\,
            I => \N__60256\
        );

    \I__14182\ : InMux
    port map (
            O => \N__60256\,
            I => \N__60250\
        );

    \I__14181\ : InMux
    port map (
            O => \N__60255\,
            I => \N__60245\
        );

    \I__14180\ : InMux
    port map (
            O => \N__60254\,
            I => \N__60245\
        );

    \I__14179\ : InMux
    port map (
            O => \N__60253\,
            I => \N__60242\
        );

    \I__14178\ : LocalMux
    port map (
            O => \N__60250\,
            I => \c0.data_in_frame_12_1\
        );

    \I__14177\ : LocalMux
    port map (
            O => \N__60245\,
            I => \c0.data_in_frame_12_1\
        );

    \I__14176\ : LocalMux
    port map (
            O => \N__60242\,
            I => \c0.data_in_frame_12_1\
        );

    \I__14175\ : InMux
    port map (
            O => \N__60235\,
            I => \N__60229\
        );

    \I__14174\ : InMux
    port map (
            O => \N__60234\,
            I => \N__60226\
        );

    \I__14173\ : InMux
    port map (
            O => \N__60233\,
            I => \N__60223\
        );

    \I__14172\ : InMux
    port map (
            O => \N__60232\,
            I => \N__60220\
        );

    \I__14171\ : LocalMux
    port map (
            O => \N__60229\,
            I => \c0.data_in_frame_12_2\
        );

    \I__14170\ : LocalMux
    port map (
            O => \N__60226\,
            I => \c0.data_in_frame_12_2\
        );

    \I__14169\ : LocalMux
    port map (
            O => \N__60223\,
            I => \c0.data_in_frame_12_2\
        );

    \I__14168\ : LocalMux
    port map (
            O => \N__60220\,
            I => \c0.data_in_frame_12_2\
        );

    \I__14167\ : CascadeMux
    port map (
            O => \N__60211\,
            I => \N__60208\
        );

    \I__14166\ : InMux
    port map (
            O => \N__60208\,
            I => \N__60204\
        );

    \I__14165\ : InMux
    port map (
            O => \N__60207\,
            I => \N__60201\
        );

    \I__14164\ : LocalMux
    port map (
            O => \N__60204\,
            I => \c0.data_in_frame_13_2\
        );

    \I__14163\ : LocalMux
    port map (
            O => \N__60201\,
            I => \c0.data_in_frame_13_2\
        );

    \I__14162\ : InMux
    port map (
            O => \N__60196\,
            I => \N__60192\
        );

    \I__14161\ : CascadeMux
    port map (
            O => \N__60195\,
            I => \N__60188\
        );

    \I__14160\ : LocalMux
    port map (
            O => \N__60192\,
            I => \N__60185\
        );

    \I__14159\ : InMux
    port map (
            O => \N__60191\,
            I => \N__60182\
        );

    \I__14158\ : InMux
    port map (
            O => \N__60188\,
            I => \N__60179\
        );

    \I__14157\ : Span4Mux_h
    port map (
            O => \N__60185\,
            I => \N__60176\
        );

    \I__14156\ : LocalMux
    port map (
            O => \N__60182\,
            I => \N__60173\
        );

    \I__14155\ : LocalMux
    port map (
            O => \N__60179\,
            I => \N__60169\
        );

    \I__14154\ : Span4Mux_v
    port map (
            O => \N__60176\,
            I => \N__60164\
        );

    \I__14153\ : Span4Mux_h
    port map (
            O => \N__60173\,
            I => \N__60164\
        );

    \I__14152\ : InMux
    port map (
            O => \N__60172\,
            I => \N__60161\
        );

    \I__14151\ : Odrv4
    port map (
            O => \N__60169\,
            I => \c0.data_in_frame_13_1\
        );

    \I__14150\ : Odrv4
    port map (
            O => \N__60164\,
            I => \c0.data_in_frame_13_1\
        );

    \I__14149\ : LocalMux
    port map (
            O => \N__60161\,
            I => \c0.data_in_frame_13_1\
        );

    \I__14148\ : CascadeMux
    port map (
            O => \N__60154\,
            I => \N__60151\
        );

    \I__14147\ : InMux
    port map (
            O => \N__60151\,
            I => \N__60147\
        );

    \I__14146\ : CascadeMux
    port map (
            O => \N__60150\,
            I => \N__60144\
        );

    \I__14145\ : LocalMux
    port map (
            O => \N__60147\,
            I => \N__60140\
        );

    \I__14144\ : InMux
    port map (
            O => \N__60144\,
            I => \N__60134\
        );

    \I__14143\ : InMux
    port map (
            O => \N__60143\,
            I => \N__60134\
        );

    \I__14142\ : Span4Mux_h
    port map (
            O => \N__60140\,
            I => \N__60131\
        );

    \I__14141\ : InMux
    port map (
            O => \N__60139\,
            I => \N__60128\
        );

    \I__14140\ : LocalMux
    port map (
            O => \N__60134\,
            I => \c0.data_in_frame_11_0\
        );

    \I__14139\ : Odrv4
    port map (
            O => \N__60131\,
            I => \c0.data_in_frame_11_0\
        );

    \I__14138\ : LocalMux
    port map (
            O => \N__60128\,
            I => \c0.data_in_frame_11_0\
        );

    \I__14137\ : InMux
    port map (
            O => \N__60121\,
            I => \N__60118\
        );

    \I__14136\ : LocalMux
    port map (
            O => \N__60118\,
            I => \N__60114\
        );

    \I__14135\ : InMux
    port map (
            O => \N__60117\,
            I => \N__60111\
        );

    \I__14134\ : Span4Mux_h
    port map (
            O => \N__60114\,
            I => \N__60108\
        );

    \I__14133\ : LocalMux
    port map (
            O => \N__60111\,
            I => \c0.n22274\
        );

    \I__14132\ : Odrv4
    port map (
            O => \N__60108\,
            I => \c0.n22274\
        );

    \I__14131\ : InMux
    port map (
            O => \N__60103\,
            I => \N__60098\
        );

    \I__14130\ : InMux
    port map (
            O => \N__60102\,
            I => \N__60095\
        );

    \I__14129\ : InMux
    port map (
            O => \N__60101\,
            I => \N__60091\
        );

    \I__14128\ : LocalMux
    port map (
            O => \N__60098\,
            I => \N__60088\
        );

    \I__14127\ : LocalMux
    port map (
            O => \N__60095\,
            I => \N__60085\
        );

    \I__14126\ : CascadeMux
    port map (
            O => \N__60094\,
            I => \N__60082\
        );

    \I__14125\ : LocalMux
    port map (
            O => \N__60091\,
            I => \N__60078\
        );

    \I__14124\ : Span4Mux_v
    port map (
            O => \N__60088\,
            I => \N__60073\
        );

    \I__14123\ : Span4Mux_h
    port map (
            O => \N__60085\,
            I => \N__60073\
        );

    \I__14122\ : InMux
    port map (
            O => \N__60082\,
            I => \N__60068\
        );

    \I__14121\ : InMux
    port map (
            O => \N__60081\,
            I => \N__60068\
        );

    \I__14120\ : Odrv12
    port map (
            O => \N__60078\,
            I => \c0.data_in_frame_10_6\
        );

    \I__14119\ : Odrv4
    port map (
            O => \N__60073\,
            I => \c0.data_in_frame_10_6\
        );

    \I__14118\ : LocalMux
    port map (
            O => \N__60068\,
            I => \c0.data_in_frame_10_6\
        );

    \I__14117\ : CascadeMux
    port map (
            O => \N__60061\,
            I => \c0.n13999_cascade_\
        );

    \I__14116\ : InMux
    port map (
            O => \N__60058\,
            I => \N__60055\
        );

    \I__14115\ : LocalMux
    port map (
            O => \N__60055\,
            I => \N__60051\
        );

    \I__14114\ : InMux
    port map (
            O => \N__60054\,
            I => \N__60048\
        );

    \I__14113\ : Span4Mux_h
    port map (
            O => \N__60051\,
            I => \N__60045\
        );

    \I__14112\ : LocalMux
    port map (
            O => \N__60048\,
            I => \N__60042\
        );

    \I__14111\ : Odrv4
    port map (
            O => \N__60045\,
            I => \c0.n21940\
        );

    \I__14110\ : Odrv4
    port map (
            O => \N__60042\,
            I => \c0.n21940\
        );

    \I__14109\ : CascadeMux
    port map (
            O => \N__60037\,
            I => \N__60034\
        );

    \I__14108\ : InMux
    port map (
            O => \N__60034\,
            I => \N__60031\
        );

    \I__14107\ : LocalMux
    port map (
            O => \N__60031\,
            I => \N__60027\
        );

    \I__14106\ : InMux
    port map (
            O => \N__60030\,
            I => \N__60024\
        );

    \I__14105\ : Span4Mux_h
    port map (
            O => \N__60027\,
            I => \N__60021\
        );

    \I__14104\ : LocalMux
    port map (
            O => \N__60024\,
            I => \N__60018\
        );

    \I__14103\ : Span4Mux_v
    port map (
            O => \N__60021\,
            I => \N__60015\
        );

    \I__14102\ : Span4Mux_h
    port map (
            O => \N__60018\,
            I => \N__60012\
        );

    \I__14101\ : Odrv4
    port map (
            O => \N__60015\,
            I => \c0.n13233\
        );

    \I__14100\ : Odrv4
    port map (
            O => \N__60012\,
            I => \c0.n13233\
        );

    \I__14099\ : InMux
    port map (
            O => \N__60007\,
            I => \N__60004\
        );

    \I__14098\ : LocalMux
    port map (
            O => \N__60004\,
            I => \N__59999\
        );

    \I__14097\ : InMux
    port map (
            O => \N__60003\,
            I => \N__59996\
        );

    \I__14096\ : InMux
    port map (
            O => \N__60002\,
            I => \N__59993\
        );

    \I__14095\ : Span4Mux_h
    port map (
            O => \N__59999\,
            I => \N__59990\
        );

    \I__14094\ : LocalMux
    port map (
            O => \N__59996\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14093\ : LocalMux
    port map (
            O => \N__59993\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14092\ : Odrv4
    port map (
            O => \N__59990\,
            I => \c0.data_in_frame_9_2\
        );

    \I__14091\ : InMux
    port map (
            O => \N__59983\,
            I => \N__59980\
        );

    \I__14090\ : LocalMux
    port map (
            O => \N__59980\,
            I => \N__59977\
        );

    \I__14089\ : Span4Mux_v
    port map (
            O => \N__59977\,
            I => \N__59973\
        );

    \I__14088\ : InMux
    port map (
            O => \N__59976\,
            I => \N__59970\
        );

    \I__14087\ : Odrv4
    port map (
            O => \N__59973\,
            I => \c0.n13993\
        );

    \I__14086\ : LocalMux
    port map (
            O => \N__59970\,
            I => \c0.n13993\
        );

    \I__14085\ : InMux
    port map (
            O => \N__59965\,
            I => \N__59962\
        );

    \I__14084\ : LocalMux
    port map (
            O => \N__59962\,
            I => \N__59959\
        );

    \I__14083\ : Span4Mux_h
    port map (
            O => \N__59959\,
            I => \N__59954\
        );

    \I__14082\ : InMux
    port map (
            O => \N__59958\,
            I => \N__59949\
        );

    \I__14081\ : InMux
    port map (
            O => \N__59957\,
            I => \N__59949\
        );

    \I__14080\ : Odrv4
    port map (
            O => \N__59954\,
            I => n91
        );

    \I__14079\ : LocalMux
    port map (
            O => \N__59949\,
            I => n91
        );

    \I__14078\ : InMux
    port map (
            O => \N__59944\,
            I => \N__59941\
        );

    \I__14077\ : LocalMux
    port map (
            O => \N__59941\,
            I => \N__59936\
        );

    \I__14076\ : InMux
    port map (
            O => \N__59940\,
            I => \N__59933\
        );

    \I__14075\ : InMux
    port map (
            O => \N__59939\,
            I => \N__59930\
        );

    \I__14074\ : Span4Mux_v
    port map (
            O => \N__59936\,
            I => \N__59925\
        );

    \I__14073\ : LocalMux
    port map (
            O => \N__59933\,
            I => \N__59925\
        );

    \I__14072\ : LocalMux
    port map (
            O => \N__59930\,
            I => \N__59922\
        );

    \I__14071\ : Span4Mux_h
    port map (
            O => \N__59925\,
            I => \N__59919\
        );

    \I__14070\ : Span4Mux_v
    port map (
            O => \N__59922\,
            I => \N__59914\
        );

    \I__14069\ : Span4Mux_v
    port map (
            O => \N__59919\,
            I => \N__59914\
        );

    \I__14068\ : Odrv4
    port map (
            O => \N__59914\,
            I => n12973
        );

    \I__14067\ : InMux
    port map (
            O => \N__59911\,
            I => \N__59907\
        );

    \I__14066\ : InMux
    port map (
            O => \N__59910\,
            I => \N__59904\
        );

    \I__14065\ : LocalMux
    port map (
            O => \N__59907\,
            I => n14917
        );

    \I__14064\ : LocalMux
    port map (
            O => \N__59904\,
            I => n14917
        );

    \I__14063\ : InMux
    port map (
            O => \N__59899\,
            I => \N__59894\
        );

    \I__14062\ : InMux
    port map (
            O => \N__59898\,
            I => \N__59889\
        );

    \I__14061\ : InMux
    port map (
            O => \N__59897\,
            I => \N__59889\
        );

    \I__14060\ : LocalMux
    port map (
            O => \N__59894\,
            I => n14436
        );

    \I__14059\ : LocalMux
    port map (
            O => \N__59889\,
            I => n14436
        );

    \I__14058\ : InMux
    port map (
            O => \N__59884\,
            I => \N__59880\
        );

    \I__14057\ : InMux
    port map (
            O => \N__59883\,
            I => \N__59877\
        );

    \I__14056\ : LocalMux
    port map (
            O => \N__59880\,
            I => \N__59874\
        );

    \I__14055\ : LocalMux
    port map (
            O => \N__59877\,
            I => \N__59869\
        );

    \I__14054\ : Span4Mux_v
    port map (
            O => \N__59874\,
            I => \N__59869\
        );

    \I__14053\ : Span4Mux_h
    port map (
            O => \N__59869\,
            I => \N__59865\
        );

    \I__14052\ : CascadeMux
    port map (
            O => \N__59868\,
            I => \N__59860\
        );

    \I__14051\ : Span4Mux_v
    port map (
            O => \N__59865\,
            I => \N__59856\
        );

    \I__14050\ : InMux
    port map (
            O => \N__59864\,
            I => \N__59853\
        );

    \I__14049\ : InMux
    port map (
            O => \N__59863\,
            I => \N__59850\
        );

    \I__14048\ : InMux
    port map (
            O => \N__59860\,
            I => \N__59845\
        );

    \I__14047\ : InMux
    port map (
            O => \N__59859\,
            I => \N__59845\
        );

    \I__14046\ : Span4Mux_h
    port map (
            O => \N__59856\,
            I => \N__59842\
        );

    \I__14045\ : LocalMux
    port map (
            O => \N__59853\,
            I => \r_Bit_Index_1\
        );

    \I__14044\ : LocalMux
    port map (
            O => \N__59850\,
            I => \r_Bit_Index_1\
        );

    \I__14043\ : LocalMux
    port map (
            O => \N__59845\,
            I => \r_Bit_Index_1\
        );

    \I__14042\ : Odrv4
    port map (
            O => \N__59842\,
            I => \r_Bit_Index_1\
        );

    \I__14041\ : InMux
    port map (
            O => \N__59833\,
            I => \N__59829\
        );

    \I__14040\ : CascadeMux
    port map (
            O => \N__59832\,
            I => \N__59826\
        );

    \I__14039\ : LocalMux
    port map (
            O => \N__59829\,
            I => \N__59823\
        );

    \I__14038\ : InMux
    port map (
            O => \N__59826\,
            I => \N__59820\
        );

    \I__14037\ : Span4Mux_v
    port map (
            O => \N__59823\,
            I => \N__59817\
        );

    \I__14036\ : LocalMux
    port map (
            O => \N__59820\,
            I => \N__59812\
        );

    \I__14035\ : Span4Mux_v
    port map (
            O => \N__59817\,
            I => \N__59812\
        );

    \I__14034\ : Span4Mux_v
    port map (
            O => \N__59812\,
            I => \N__59808\
        );

    \I__14033\ : InMux
    port map (
            O => \N__59811\,
            I => \N__59805\
        );

    \I__14032\ : Span4Mux_h
    port map (
            O => \N__59808\,
            I => \N__59802\
        );

    \I__14031\ : LocalMux
    port map (
            O => \N__59805\,
            I => data_in_frame_22_4
        );

    \I__14030\ : Odrv4
    port map (
            O => \N__59802\,
            I => data_in_frame_22_4
        );

    \I__14029\ : CascadeMux
    port map (
            O => \N__59797\,
            I => \N__59794\
        );

    \I__14028\ : InMux
    port map (
            O => \N__59794\,
            I => \N__59791\
        );

    \I__14027\ : LocalMux
    port map (
            O => \N__59791\,
            I => \N__59788\
        );

    \I__14026\ : Span4Mux_h
    port map (
            O => \N__59788\,
            I => \N__59784\
        );

    \I__14025\ : InMux
    port map (
            O => \N__59787\,
            I => \N__59781\
        );

    \I__14024\ : Span4Mux_v
    port map (
            O => \N__59784\,
            I => \N__59778\
        );

    \I__14023\ : LocalMux
    port map (
            O => \N__59781\,
            I => \N__59775\
        );

    \I__14022\ : Odrv4
    port map (
            O => \N__59778\,
            I => \c0.n22191\
        );

    \I__14021\ : Odrv12
    port map (
            O => \N__59775\,
            I => \c0.n22191\
        );

    \I__14020\ : InMux
    port map (
            O => \N__59770\,
            I => \N__59767\
        );

    \I__14019\ : LocalMux
    port map (
            O => \N__59767\,
            I => \N__59764\
        );

    \I__14018\ : Span4Mux_h
    port map (
            O => \N__59764\,
            I => \N__59761\
        );

    \I__14017\ : Odrv4
    port map (
            O => \N__59761\,
            I => \c0.n25\
        );

    \I__14016\ : CascadeMux
    port map (
            O => \N__59758\,
            I => \N__59753\
        );

    \I__14015\ : InMux
    port map (
            O => \N__59757\,
            I => \N__59740\
        );

    \I__14014\ : InMux
    port map (
            O => \N__59756\,
            I => \N__59740\
        );

    \I__14013\ : InMux
    port map (
            O => \N__59753\,
            I => \N__59740\
        );

    \I__14012\ : InMux
    port map (
            O => \N__59752\,
            I => \N__59733\
        );

    \I__14011\ : InMux
    port map (
            O => \N__59751\,
            I => \N__59733\
        );

    \I__14010\ : InMux
    port map (
            O => \N__59750\,
            I => \N__59733\
        );

    \I__14009\ : InMux
    port map (
            O => \N__59749\,
            I => \N__59728\
        );

    \I__14008\ : InMux
    port map (
            O => \N__59748\,
            I => \N__59728\
        );

    \I__14007\ : InMux
    port map (
            O => \N__59747\,
            I => \N__59725\
        );

    \I__14006\ : LocalMux
    port map (
            O => \N__59740\,
            I => \r_Bit_Index_0\
        );

    \I__14005\ : LocalMux
    port map (
            O => \N__59733\,
            I => \r_Bit_Index_0\
        );

    \I__14004\ : LocalMux
    port map (
            O => \N__59728\,
            I => \r_Bit_Index_0\
        );

    \I__14003\ : LocalMux
    port map (
            O => \N__59725\,
            I => \r_Bit_Index_0\
        );

    \I__14002\ : CascadeMux
    port map (
            O => \N__59716\,
            I => \N__59712\
        );

    \I__14001\ : CascadeMux
    port map (
            O => \N__59715\,
            I => \N__59705\
        );

    \I__14000\ : InMux
    port map (
            O => \N__59712\,
            I => \N__59700\
        );

    \I__13999\ : InMux
    port map (
            O => \N__59711\,
            I => \N__59700\
        );

    \I__13998\ : CascadeMux
    port map (
            O => \N__59710\,
            I => \N__59695\
        );

    \I__13997\ : CascadeMux
    port map (
            O => \N__59709\,
            I => \N__59691\
        );

    \I__13996\ : InMux
    port map (
            O => \N__59708\,
            I => \N__59685\
        );

    \I__13995\ : InMux
    port map (
            O => \N__59705\,
            I => \N__59685\
        );

    \I__13994\ : LocalMux
    port map (
            O => \N__59700\,
            I => \N__59682\
        );

    \I__13993\ : InMux
    port map (
            O => \N__59699\,
            I => \N__59677\
        );

    \I__13992\ : InMux
    port map (
            O => \N__59698\,
            I => \N__59677\
        );

    \I__13991\ : InMux
    port map (
            O => \N__59695\,
            I => \N__59672\
        );

    \I__13990\ : InMux
    port map (
            O => \N__59694\,
            I => \N__59672\
        );

    \I__13989\ : InMux
    port map (
            O => \N__59691\,
            I => \N__59669\
        );

    \I__13988\ : CascadeMux
    port map (
            O => \N__59690\,
            I => \N__59666\
        );

    \I__13987\ : LocalMux
    port map (
            O => \N__59685\,
            I => \N__59659\
        );

    \I__13986\ : Span4Mux_h
    port map (
            O => \N__59682\,
            I => \N__59659\
        );

    \I__13985\ : LocalMux
    port map (
            O => \N__59677\,
            I => \N__59659\
        );

    \I__13984\ : LocalMux
    port map (
            O => \N__59672\,
            I => \N__59656\
        );

    \I__13983\ : LocalMux
    port map (
            O => \N__59669\,
            I => \N__59650\
        );

    \I__13982\ : InMux
    port map (
            O => \N__59666\,
            I => \N__59647\
        );

    \I__13981\ : Span4Mux_h
    port map (
            O => \N__59659\,
            I => \N__59644\
        );

    \I__13980\ : Span4Mux_v
    port map (
            O => \N__59656\,
            I => \N__59641\
        );

    \I__13979\ : InMux
    port map (
            O => \N__59655\,
            I => \N__59634\
        );

    \I__13978\ : InMux
    port map (
            O => \N__59654\,
            I => \N__59634\
        );

    \I__13977\ : InMux
    port map (
            O => \N__59653\,
            I => \N__59634\
        );

    \I__13976\ : Span4Mux_v
    port map (
            O => \N__59650\,
            I => \N__59631\
        );

    \I__13975\ : LocalMux
    port map (
            O => \N__59647\,
            I => \N__59628\
        );

    \I__13974\ : Span4Mux_v
    port map (
            O => \N__59644\,
            I => \N__59625\
        );

    \I__13973\ : Sp12to4
    port map (
            O => \N__59641\,
            I => \N__59620\
        );

    \I__13972\ : LocalMux
    port map (
            O => \N__59634\,
            I => \N__59620\
        );

    \I__13971\ : Span4Mux_v
    port map (
            O => \N__59631\,
            I => \N__59617\
        );

    \I__13970\ : Span12Mux_h
    port map (
            O => \N__59628\,
            I => \N__59610\
        );

    \I__13969\ : Sp12to4
    port map (
            O => \N__59625\,
            I => \N__59610\
        );

    \I__13968\ : Span12Mux_v
    port map (
            O => \N__59620\,
            I => \N__59610\
        );

    \I__13967\ : Span4Mux_v
    port map (
            O => \N__59617\,
            I => \N__59607\
        );

    \I__13966\ : Span12Mux_h
    port map (
            O => \N__59610\,
            I => \N__59604\
        );

    \I__13965\ : Span4Mux_v
    port map (
            O => \N__59607\,
            I => \N__59601\
        );

    \I__13964\ : Span12Mux_v
    port map (
            O => \N__59604\,
            I => \N__59598\
        );

    \I__13963\ : Odrv4
    port map (
            O => \N__59601\,
            I => \r_Rx_Data\
        );

    \I__13962\ : Odrv12
    port map (
            O => \N__59598\,
            I => \r_Rx_Data\
        );

    \I__13961\ : CascadeMux
    port map (
            O => \N__59593\,
            I => \N__59589\
        );

    \I__13960\ : InMux
    port map (
            O => \N__59592\,
            I => \N__59584\
        );

    \I__13959\ : InMux
    port map (
            O => \N__59589\,
            I => \N__59584\
        );

    \I__13958\ : LocalMux
    port map (
            O => \N__59584\,
            I => n12970
        );

    \I__13957\ : InMux
    port map (
            O => \N__59581\,
            I => \N__59575\
        );

    \I__13956\ : InMux
    port map (
            O => \N__59580\,
            I => \N__59572\
        );

    \I__13955\ : InMux
    port map (
            O => \N__59579\,
            I => \N__59569\
        );

    \I__13954\ : CascadeMux
    port map (
            O => \N__59578\,
            I => \N__59566\
        );

    \I__13953\ : LocalMux
    port map (
            O => \N__59575\,
            I => \N__59563\
        );

    \I__13952\ : LocalMux
    port map (
            O => \N__59572\,
            I => \N__59558\
        );

    \I__13951\ : LocalMux
    port map (
            O => \N__59569\,
            I => \N__59558\
        );

    \I__13950\ : InMux
    port map (
            O => \N__59566\,
            I => \N__59555\
        );

    \I__13949\ : Span4Mux_h
    port map (
            O => \N__59563\,
            I => \N__59552\
        );

    \I__13948\ : Span4Mux_h
    port map (
            O => \N__59558\,
            I => \N__59549\
        );

    \I__13947\ : LocalMux
    port map (
            O => \N__59555\,
            I => \c0.data_in_frame_12_0\
        );

    \I__13946\ : Odrv4
    port map (
            O => \N__59552\,
            I => \c0.data_in_frame_12_0\
        );

    \I__13945\ : Odrv4
    port map (
            O => \N__59549\,
            I => \c0.data_in_frame_12_0\
        );

    \I__13944\ : InMux
    port map (
            O => \N__59542\,
            I => \N__59538\
        );

    \I__13943\ : InMux
    port map (
            O => \N__59541\,
            I => \N__59535\
        );

    \I__13942\ : LocalMux
    port map (
            O => \N__59538\,
            I => \N__59528\
        );

    \I__13941\ : LocalMux
    port map (
            O => \N__59535\,
            I => \N__59528\
        );

    \I__13940\ : InMux
    port map (
            O => \N__59534\,
            I => \N__59523\
        );

    \I__13939\ : InMux
    port map (
            O => \N__59533\,
            I => \N__59523\
        );

    \I__13938\ : Span4Mux_v
    port map (
            O => \N__59528\,
            I => \N__59517\
        );

    \I__13937\ : LocalMux
    port map (
            O => \N__59523\,
            I => \N__59517\
        );

    \I__13936\ : CascadeMux
    port map (
            O => \N__59522\,
            I => \N__59514\
        );

    \I__13935\ : Span4Mux_v
    port map (
            O => \N__59517\,
            I => \N__59511\
        );

    \I__13934\ : InMux
    port map (
            O => \N__59514\,
            I => \N__59508\
        );

    \I__13933\ : Span4Mux_v
    port map (
            O => \N__59511\,
            I => \N__59505\
        );

    \I__13932\ : LocalMux
    port map (
            O => \N__59508\,
            I => \c0.data_in_frame_24_7\
        );

    \I__13931\ : Odrv4
    port map (
            O => \N__59505\,
            I => \c0.data_in_frame_24_7\
        );

    \I__13930\ : InMux
    port map (
            O => \N__59500\,
            I => \N__59496\
        );

    \I__13929\ : CascadeMux
    port map (
            O => \N__59499\,
            I => \N__59493\
        );

    \I__13928\ : LocalMux
    port map (
            O => \N__59496\,
            I => \N__59490\
        );

    \I__13927\ : InMux
    port map (
            O => \N__59493\,
            I => \N__59485\
        );

    \I__13926\ : Span4Mux_v
    port map (
            O => \N__59490\,
            I => \N__59482\
        );

    \I__13925\ : InMux
    port map (
            O => \N__59489\,
            I => \N__59477\
        );

    \I__13924\ : InMux
    port map (
            O => \N__59488\,
            I => \N__59477\
        );

    \I__13923\ : LocalMux
    port map (
            O => \N__59485\,
            I => \c0.data_in_frame_26_4\
        );

    \I__13922\ : Odrv4
    port map (
            O => \N__59482\,
            I => \c0.data_in_frame_26_4\
        );

    \I__13921\ : LocalMux
    port map (
            O => \N__59477\,
            I => \c0.data_in_frame_26_4\
        );

    \I__13920\ : InMux
    port map (
            O => \N__59470\,
            I => \N__59467\
        );

    \I__13919\ : LocalMux
    port map (
            O => \N__59467\,
            I => \c0.n22337\
        );

    \I__13918\ : CascadeMux
    port map (
            O => \N__59464\,
            I => \c0.n10_adj_4285_cascade_\
        );

    \I__13917\ : InMux
    port map (
            O => \N__59461\,
            I => \N__59458\
        );

    \I__13916\ : LocalMux
    port map (
            O => \N__59458\,
            I => \N__59455\
        );

    \I__13915\ : Span4Mux_h
    port map (
            O => \N__59455\,
            I => \N__59452\
        );

    \I__13914\ : Span4Mux_h
    port map (
            O => \N__59452\,
            I => \N__59449\
        );

    \I__13913\ : Odrv4
    port map (
            O => \N__59449\,
            I => \c0.n22995\
        );

    \I__13912\ : InMux
    port map (
            O => \N__59446\,
            I => \N__59440\
        );

    \I__13911\ : InMux
    port map (
            O => \N__59445\,
            I => \N__59440\
        );

    \I__13910\ : LocalMux
    port map (
            O => \N__59440\,
            I => \N__59436\
        );

    \I__13909\ : CascadeMux
    port map (
            O => \N__59439\,
            I => \N__59433\
        );

    \I__13908\ : Span4Mux_h
    port map (
            O => \N__59436\,
            I => \N__59430\
        );

    \I__13907\ : InMux
    port map (
            O => \N__59433\,
            I => \N__59427\
        );

    \I__13906\ : Span4Mux_v
    port map (
            O => \N__59430\,
            I => \N__59424\
        );

    \I__13905\ : LocalMux
    port map (
            O => \N__59427\,
            I => \c0.data_in_frame_26_6\
        );

    \I__13904\ : Odrv4
    port map (
            O => \N__59424\,
            I => \c0.data_in_frame_26_6\
        );

    \I__13903\ : InMux
    port map (
            O => \N__59419\,
            I => \N__59416\
        );

    \I__13902\ : LocalMux
    port map (
            O => \N__59416\,
            I => \N__59413\
        );

    \I__13901\ : Odrv4
    port map (
            O => \N__59413\,
            I => \c0.n22054\
        );

    \I__13900\ : InMux
    port map (
            O => \N__59410\,
            I => \N__59402\
        );

    \I__13899\ : InMux
    port map (
            O => \N__59409\,
            I => \N__59402\
        );

    \I__13898\ : CascadeMux
    port map (
            O => \N__59408\,
            I => \N__59397\
        );

    \I__13897\ : CascadeMux
    port map (
            O => \N__59407\,
            I => \N__59394\
        );

    \I__13896\ : LocalMux
    port map (
            O => \N__59402\,
            I => \N__59390\
        );

    \I__13895\ : InMux
    port map (
            O => \N__59401\,
            I => \N__59385\
        );

    \I__13894\ : InMux
    port map (
            O => \N__59400\,
            I => \N__59385\
        );

    \I__13893\ : InMux
    port map (
            O => \N__59397\,
            I => \N__59382\
        );

    \I__13892\ : InMux
    port map (
            O => \N__59394\,
            I => \N__59377\
        );

    \I__13891\ : InMux
    port map (
            O => \N__59393\,
            I => \N__59377\
        );

    \I__13890\ : Span4Mux_v
    port map (
            O => \N__59390\,
            I => \N__59372\
        );

    \I__13889\ : LocalMux
    port map (
            O => \N__59385\,
            I => \N__59372\
        );

    \I__13888\ : LocalMux
    port map (
            O => \N__59382\,
            I => \c0.data_in_frame_24_6\
        );

    \I__13887\ : LocalMux
    port map (
            O => \N__59377\,
            I => \c0.data_in_frame_24_6\
        );

    \I__13886\ : Odrv4
    port map (
            O => \N__59372\,
            I => \c0.data_in_frame_24_6\
        );

    \I__13885\ : CascadeMux
    port map (
            O => \N__59365\,
            I => \N__59362\
        );

    \I__13884\ : InMux
    port map (
            O => \N__59362\,
            I => \N__59359\
        );

    \I__13883\ : LocalMux
    port map (
            O => \N__59359\,
            I => \N__59356\
        );

    \I__13882\ : Odrv12
    port map (
            O => \N__59356\,
            I => \c0.n22434\
        );

    \I__13881\ : InMux
    port map (
            O => \N__59353\,
            I => \N__59349\
        );

    \I__13880\ : InMux
    port map (
            O => \N__59352\,
            I => \N__59346\
        );

    \I__13879\ : LocalMux
    port map (
            O => \N__59349\,
            I => \N__59343\
        );

    \I__13878\ : LocalMux
    port map (
            O => \N__59346\,
            I => \N__59340\
        );

    \I__13877\ : Span4Mux_v
    port map (
            O => \N__59343\,
            I => \N__59337\
        );

    \I__13876\ : Span4Mux_v
    port map (
            O => \N__59340\,
            I => \N__59332\
        );

    \I__13875\ : Sp12to4
    port map (
            O => \N__59337\,
            I => \N__59329\
        );

    \I__13874\ : InMux
    port map (
            O => \N__59336\,
            I => \N__59324\
        );

    \I__13873\ : InMux
    port map (
            O => \N__59335\,
            I => \N__59324\
        );

    \I__13872\ : Odrv4
    port map (
            O => \N__59332\,
            I => \c0.data_in_frame_20_0\
        );

    \I__13871\ : Odrv12
    port map (
            O => \N__59329\,
            I => \c0.data_in_frame_20_0\
        );

    \I__13870\ : LocalMux
    port map (
            O => \N__59324\,
            I => \c0.data_in_frame_20_0\
        );

    \I__13869\ : CascadeMux
    port map (
            O => \N__59317\,
            I => \N__59314\
        );

    \I__13868\ : InMux
    port map (
            O => \N__59314\,
            I => \N__59311\
        );

    \I__13867\ : LocalMux
    port map (
            O => \N__59311\,
            I => \N__59307\
        );

    \I__13866\ : InMux
    port map (
            O => \N__59310\,
            I => \N__59303\
        );

    \I__13865\ : Span12Mux_h
    port map (
            O => \N__59307\,
            I => \N__59300\
        );

    \I__13864\ : InMux
    port map (
            O => \N__59306\,
            I => \N__59297\
        );

    \I__13863\ : LocalMux
    port map (
            O => \N__59303\,
            I => data_in_frame_22_2
        );

    \I__13862\ : Odrv12
    port map (
            O => \N__59300\,
            I => data_in_frame_22_2
        );

    \I__13861\ : LocalMux
    port map (
            O => \N__59297\,
            I => data_in_frame_22_2
        );

    \I__13860\ : InMux
    port map (
            O => \N__59290\,
            I => \N__59286\
        );

    \I__13859\ : InMux
    port map (
            O => \N__59289\,
            I => \N__59283\
        );

    \I__13858\ : LocalMux
    port map (
            O => \N__59286\,
            I => \N__59280\
        );

    \I__13857\ : LocalMux
    port map (
            O => \N__59283\,
            I => \N__59275\
        );

    \I__13856\ : Span4Mux_v
    port map (
            O => \N__59280\,
            I => \N__59272\
        );

    \I__13855\ : InMux
    port map (
            O => \N__59279\,
            I => \N__59269\
        );

    \I__13854\ : InMux
    port map (
            O => \N__59278\,
            I => \N__59266\
        );

    \I__13853\ : Odrv4
    port map (
            O => \N__59275\,
            I => \c0.n12594\
        );

    \I__13852\ : Odrv4
    port map (
            O => \N__59272\,
            I => \c0.n12594\
        );

    \I__13851\ : LocalMux
    port map (
            O => \N__59269\,
            I => \c0.n12594\
        );

    \I__13850\ : LocalMux
    port map (
            O => \N__59266\,
            I => \c0.n12594\
        );

    \I__13849\ : InMux
    port map (
            O => \N__59257\,
            I => \N__59253\
        );

    \I__13848\ : InMux
    port map (
            O => \N__59256\,
            I => \N__59250\
        );

    \I__13847\ : LocalMux
    port map (
            O => \N__59253\,
            I => \c0.n20596\
        );

    \I__13846\ : LocalMux
    port map (
            O => \N__59250\,
            I => \c0.n20596\
        );

    \I__13845\ : InMux
    port map (
            O => \N__59245\,
            I => \N__59241\
        );

    \I__13844\ : InMux
    port map (
            O => \N__59244\,
            I => \N__59238\
        );

    \I__13843\ : LocalMux
    port map (
            O => \N__59241\,
            I => \N__59235\
        );

    \I__13842\ : LocalMux
    port map (
            O => \N__59238\,
            I => \N__59232\
        );

    \I__13841\ : Span4Mux_v
    port map (
            O => \N__59235\,
            I => \N__59227\
        );

    \I__13840\ : Span4Mux_h
    port map (
            O => \N__59232\,
            I => \N__59227\
        );

    \I__13839\ : Span4Mux_v
    port map (
            O => \N__59227\,
            I => \N__59223\
        );

    \I__13838\ : InMux
    port map (
            O => \N__59226\,
            I => \N__59220\
        );

    \I__13837\ : Span4Mux_v
    port map (
            O => \N__59223\,
            I => \N__59217\
        );

    \I__13836\ : LocalMux
    port map (
            O => \N__59220\,
            I => \c0.data_in_frame_11_7\
        );

    \I__13835\ : Odrv4
    port map (
            O => \N__59217\,
            I => \c0.data_in_frame_11_7\
        );

    \I__13834\ : InMux
    port map (
            O => \N__59212\,
            I => \N__59207\
        );

    \I__13833\ : InMux
    port map (
            O => \N__59211\,
            I => \N__59204\
        );

    \I__13832\ : InMux
    port map (
            O => \N__59210\,
            I => \N__59201\
        );

    \I__13831\ : LocalMux
    port map (
            O => \N__59207\,
            I => \N__59195\
        );

    \I__13830\ : LocalMux
    port map (
            O => \N__59204\,
            I => \N__59190\
        );

    \I__13829\ : LocalMux
    port map (
            O => \N__59201\,
            I => \N__59190\
        );

    \I__13828\ : InMux
    port map (
            O => \N__59200\,
            I => \N__59187\
        );

    \I__13827\ : InMux
    port map (
            O => \N__59199\,
            I => \N__59184\
        );

    \I__13826\ : InMux
    port map (
            O => \N__59198\,
            I => \N__59181\
        );

    \I__13825\ : Span4Mux_v
    port map (
            O => \N__59195\,
            I => \N__59178\
        );

    \I__13824\ : Span4Mux_v
    port map (
            O => \N__59190\,
            I => \N__59173\
        );

    \I__13823\ : LocalMux
    port map (
            O => \N__59187\,
            I => \N__59173\
        );

    \I__13822\ : LocalMux
    port map (
            O => \N__59184\,
            I => \N__59170\
        );

    \I__13821\ : LocalMux
    port map (
            O => \N__59181\,
            I => \N__59165\
        );

    \I__13820\ : Span4Mux_v
    port map (
            O => \N__59178\,
            I => \N__59162\
        );

    \I__13819\ : Span4Mux_v
    port map (
            O => \N__59173\,
            I => \N__59157\
        );

    \I__13818\ : Span4Mux_v
    port map (
            O => \N__59170\,
            I => \N__59157\
        );

    \I__13817\ : InMux
    port map (
            O => \N__59169\,
            I => \N__59154\
        );

    \I__13816\ : InMux
    port map (
            O => \N__59168\,
            I => \N__59151\
        );

    \I__13815\ : Span4Mux_v
    port map (
            O => \N__59165\,
            I => \N__59148\
        );

    \I__13814\ : Sp12to4
    port map (
            O => \N__59162\,
            I => \N__59141\
        );

    \I__13813\ : Sp12to4
    port map (
            O => \N__59157\,
            I => \N__59141\
        );

    \I__13812\ : LocalMux
    port map (
            O => \N__59154\,
            I => \N__59141\
        );

    \I__13811\ : LocalMux
    port map (
            O => \N__59151\,
            I => \N__59138\
        );

    \I__13810\ : Sp12to4
    port map (
            O => \N__59148\,
            I => \N__59135\
        );

    \I__13809\ : Span12Mux_h
    port map (
            O => \N__59141\,
            I => \N__59130\
        );

    \I__13808\ : Span12Mux_h
    port map (
            O => \N__59138\,
            I => \N__59130\
        );

    \I__13807\ : Odrv12
    port map (
            O => \N__59135\,
            I => n21760
        );

    \I__13806\ : Odrv12
    port map (
            O => \N__59130\,
            I => n21760
        );

    \I__13805\ : CascadeMux
    port map (
            O => \N__59125\,
            I => \N__59122\
        );

    \I__13804\ : InMux
    port map (
            O => \N__59122\,
            I => \N__59119\
        );

    \I__13803\ : LocalMux
    port map (
            O => \N__59119\,
            I => \N__59114\
        );

    \I__13802\ : InMux
    port map (
            O => \N__59118\,
            I => \N__59109\
        );

    \I__13801\ : InMux
    port map (
            O => \N__59117\,
            I => \N__59109\
        );

    \I__13800\ : Odrv12
    port map (
            O => \N__59114\,
            I => \c0.data_in_frame_26_2\
        );

    \I__13799\ : LocalMux
    port map (
            O => \N__59109\,
            I => \c0.data_in_frame_26_2\
        );

    \I__13798\ : InMux
    port map (
            O => \N__59104\,
            I => \N__59101\
        );

    \I__13797\ : LocalMux
    port map (
            O => \N__59101\,
            I => \N__59098\
        );

    \I__13796\ : Odrv4
    port map (
            O => \N__59098\,
            I => \c0.n10_adj_4483\
        );

    \I__13795\ : CascadeMux
    port map (
            O => \N__59095\,
            I => \c0.n20537_cascade_\
        );

    \I__13794\ : InMux
    port map (
            O => \N__59092\,
            I => \N__59089\
        );

    \I__13793\ : LocalMux
    port map (
            O => \N__59089\,
            I => \N__59086\
        );

    \I__13792\ : Span4Mux_v
    port map (
            O => \N__59086\,
            I => \N__59083\
        );

    \I__13791\ : Odrv4
    port map (
            O => \N__59083\,
            I => \c0.n14_adj_4484\
        );

    \I__13790\ : InMux
    port map (
            O => \N__59080\,
            I => \N__59074\
        );

    \I__13789\ : InMux
    port map (
            O => \N__59079\,
            I => \N__59074\
        );

    \I__13788\ : LocalMux
    port map (
            O => \N__59074\,
            I => \c0.n21890\
        );

    \I__13787\ : InMux
    port map (
            O => \N__59071\,
            I => \N__59068\
        );

    \I__13786\ : LocalMux
    port map (
            O => \N__59068\,
            I => \N__59062\
        );

    \I__13785\ : InMux
    port map (
            O => \N__59067\,
            I => \N__59059\
        );

    \I__13784\ : InMux
    port map (
            O => \N__59066\,
            I => \N__59054\
        );

    \I__13783\ : InMux
    port map (
            O => \N__59065\,
            I => \N__59054\
        );

    \I__13782\ : Odrv4
    port map (
            O => \N__59062\,
            I => \c0.n21087\
        );

    \I__13781\ : LocalMux
    port map (
            O => \N__59059\,
            I => \c0.n21087\
        );

    \I__13780\ : LocalMux
    port map (
            O => \N__59054\,
            I => \c0.n21087\
        );

    \I__13779\ : CascadeMux
    port map (
            O => \N__59047\,
            I => \c0.n13320_cascade_\
        );

    \I__13778\ : InMux
    port map (
            O => \N__59044\,
            I => \N__59038\
        );

    \I__13777\ : InMux
    port map (
            O => \N__59043\,
            I => \N__59038\
        );

    \I__13776\ : LocalMux
    port map (
            O => \N__59038\,
            I => \c0.n22468\
        );

    \I__13775\ : CascadeMux
    port map (
            O => \N__59035\,
            I => \c0.n10_cascade_\
        );

    \I__13774\ : InMux
    port map (
            O => \N__59032\,
            I => \N__59026\
        );

    \I__13773\ : InMux
    port map (
            O => \N__59031\,
            I => \N__59026\
        );

    \I__13772\ : LocalMux
    port map (
            O => \N__59026\,
            I => \c0.n20537\
        );

    \I__13771\ : InMux
    port map (
            O => \N__59023\,
            I => \N__59020\
        );

    \I__13770\ : LocalMux
    port map (
            O => \N__59020\,
            I => \N__59016\
        );

    \I__13769\ : InMux
    port map (
            O => \N__59019\,
            I => \N__59013\
        );

    \I__13768\ : Odrv4
    port map (
            O => \N__59016\,
            I => \c0.n22314\
        );

    \I__13767\ : LocalMux
    port map (
            O => \N__59013\,
            I => \c0.n22314\
        );

    \I__13766\ : InMux
    port map (
            O => \N__59008\,
            I => \N__59003\
        );

    \I__13765\ : InMux
    port map (
            O => \N__59007\,
            I => \N__59000\
        );

    \I__13764\ : CascadeMux
    port map (
            O => \N__59006\,
            I => \N__58997\
        );

    \I__13763\ : LocalMux
    port map (
            O => \N__59003\,
            I => \N__58993\
        );

    \I__13762\ : LocalMux
    port map (
            O => \N__59000\,
            I => \N__58990\
        );

    \I__13761\ : InMux
    port map (
            O => \N__58997\,
            I => \N__58987\
        );

    \I__13760\ : InMux
    port map (
            O => \N__58996\,
            I => \N__58984\
        );

    \I__13759\ : Span4Mux_v
    port map (
            O => \N__58993\,
            I => \N__58979\
        );

    \I__13758\ : Span4Mux_v
    port map (
            O => \N__58990\,
            I => \N__58979\
        );

    \I__13757\ : LocalMux
    port map (
            O => \N__58987\,
            I => \c0.data_in_frame_24_3\
        );

    \I__13756\ : LocalMux
    port map (
            O => \N__58984\,
            I => \c0.data_in_frame_24_3\
        );

    \I__13755\ : Odrv4
    port map (
            O => \N__58979\,
            I => \c0.data_in_frame_24_3\
        );

    \I__13754\ : InMux
    port map (
            O => \N__58972\,
            I => \N__58969\
        );

    \I__13753\ : LocalMux
    port map (
            O => \N__58969\,
            I => \N__58966\
        );

    \I__13752\ : Span4Mux_v
    port map (
            O => \N__58966\,
            I => \N__58963\
        );

    \I__13751\ : Odrv4
    port map (
            O => \N__58963\,
            I => \c0.n22142\
        );

    \I__13750\ : InMux
    port map (
            O => \N__58960\,
            I => \N__58957\
        );

    \I__13749\ : LocalMux
    port map (
            O => \N__58957\,
            I => \N__58954\
        );

    \I__13748\ : Span4Mux_v
    port map (
            O => \N__58954\,
            I => \N__58949\
        );

    \I__13747\ : InMux
    port map (
            O => \N__58953\,
            I => \N__58944\
        );

    \I__13746\ : InMux
    port map (
            O => \N__58952\,
            I => \N__58944\
        );

    \I__13745\ : Span4Mux_h
    port map (
            O => \N__58949\,
            I => \N__58939\
        );

    \I__13744\ : LocalMux
    port map (
            O => \N__58944\,
            I => \N__58939\
        );

    \I__13743\ : Span4Mux_v
    port map (
            O => \N__58939\,
            I => \N__58935\
        );

    \I__13742\ : CascadeMux
    port map (
            O => \N__58938\,
            I => \N__58932\
        );

    \I__13741\ : Span4Mux_h
    port map (
            O => \N__58935\,
            I => \N__58929\
        );

    \I__13740\ : InMux
    port map (
            O => \N__58932\,
            I => \N__58926\
        );

    \I__13739\ : Span4Mux_h
    port map (
            O => \N__58929\,
            I => \N__58923\
        );

    \I__13738\ : LocalMux
    port map (
            O => \N__58926\,
            I => \c0.data_in_frame_24_4\
        );

    \I__13737\ : Odrv4
    port map (
            O => \N__58923\,
            I => \c0.data_in_frame_24_4\
        );

    \I__13736\ : InMux
    port map (
            O => \N__58918\,
            I => \N__58915\
        );

    \I__13735\ : LocalMux
    port map (
            O => \N__58915\,
            I => \N__58912\
        );

    \I__13734\ : Span4Mux_h
    port map (
            O => \N__58912\,
            I => \N__58909\
        );

    \I__13733\ : Odrv4
    port map (
            O => \N__58909\,
            I => \c0.n22028\
        );

    \I__13732\ : CascadeMux
    port map (
            O => \N__58906\,
            I => \c0.n22337_cascade_\
        );

    \I__13731\ : InMux
    port map (
            O => \N__58903\,
            I => \N__58900\
        );

    \I__13730\ : LocalMux
    port map (
            O => \N__58900\,
            I => \N__58893\
        );

    \I__13729\ : InMux
    port map (
            O => \N__58899\,
            I => \N__58890\
        );

    \I__13728\ : InMux
    port map (
            O => \N__58898\,
            I => \N__58885\
        );

    \I__13727\ : InMux
    port map (
            O => \N__58897\,
            I => \N__58885\
        );

    \I__13726\ : InMux
    port map (
            O => \N__58896\,
            I => \N__58882\
        );

    \I__13725\ : Span4Mux_h
    port map (
            O => \N__58893\,
            I => \N__58873\
        );

    \I__13724\ : LocalMux
    port map (
            O => \N__58890\,
            I => \N__58873\
        );

    \I__13723\ : LocalMux
    port map (
            O => \N__58885\,
            I => \N__58873\
        );

    \I__13722\ : LocalMux
    port map (
            O => \N__58882\,
            I => \N__58873\
        );

    \I__13721\ : Span4Mux_v
    port map (
            O => \N__58873\,
            I => \N__58870\
        );

    \I__13720\ : Odrv4
    port map (
            O => \N__58870\,
            I => \c0.n22020\
        );

    \I__13719\ : InMux
    port map (
            O => \N__58867\,
            I => \N__58861\
        );

    \I__13718\ : InMux
    port map (
            O => \N__58866\,
            I => \N__58861\
        );

    \I__13717\ : LocalMux
    port map (
            O => \N__58861\,
            I => \N__58858\
        );

    \I__13716\ : Span12Mux_v
    port map (
            O => \N__58858\,
            I => \N__58855\
        );

    \I__13715\ : Odrv12
    port map (
            O => \N__58855\,
            I => \c0.n21095\
        );

    \I__13714\ : InMux
    port map (
            O => \N__58852\,
            I => \N__58849\
        );

    \I__13713\ : LocalMux
    port map (
            O => \N__58849\,
            I => \c0.n6_adj_4418\
        );

    \I__13712\ : CascadeMux
    port map (
            O => \N__58846\,
            I => \N__58842\
        );

    \I__13711\ : CascadeMux
    port map (
            O => \N__58845\,
            I => \N__58839\
        );

    \I__13710\ : InMux
    port map (
            O => \N__58842\,
            I => \N__58832\
        );

    \I__13709\ : InMux
    port map (
            O => \N__58839\,
            I => \N__58829\
        );

    \I__13708\ : InMux
    port map (
            O => \N__58838\,
            I => \N__58826\
        );

    \I__13707\ : InMux
    port map (
            O => \N__58837\,
            I => \N__58823\
        );

    \I__13706\ : CascadeMux
    port map (
            O => \N__58836\,
            I => \N__58819\
        );

    \I__13705\ : CascadeMux
    port map (
            O => \N__58835\,
            I => \N__58816\
        );

    \I__13704\ : LocalMux
    port map (
            O => \N__58832\,
            I => \N__58813\
        );

    \I__13703\ : LocalMux
    port map (
            O => \N__58829\,
            I => \N__58810\
        );

    \I__13702\ : LocalMux
    port map (
            O => \N__58826\,
            I => \N__58807\
        );

    \I__13701\ : LocalMux
    port map (
            O => \N__58823\,
            I => \N__58804\
        );

    \I__13700\ : InMux
    port map (
            O => \N__58822\,
            I => \N__58799\
        );

    \I__13699\ : InMux
    port map (
            O => \N__58819\,
            I => \N__58799\
        );

    \I__13698\ : InMux
    port map (
            O => \N__58816\,
            I => \N__58796\
        );

    \I__13697\ : Span4Mux_h
    port map (
            O => \N__58813\,
            I => \N__58793\
        );

    \I__13696\ : Span4Mux_h
    port map (
            O => \N__58810\,
            I => \N__58788\
        );

    \I__13695\ : Span4Mux_v
    port map (
            O => \N__58807\,
            I => \N__58788\
        );

    \I__13694\ : Span4Mux_v
    port map (
            O => \N__58804\,
            I => \N__58783\
        );

    \I__13693\ : LocalMux
    port map (
            O => \N__58799\,
            I => \N__58783\
        );

    \I__13692\ : LocalMux
    port map (
            O => \N__58796\,
            I => \c0.data_in_frame_19_5\
        );

    \I__13691\ : Odrv4
    port map (
            O => \N__58793\,
            I => \c0.data_in_frame_19_5\
        );

    \I__13690\ : Odrv4
    port map (
            O => \N__58788\,
            I => \c0.data_in_frame_19_5\
        );

    \I__13689\ : Odrv4
    port map (
            O => \N__58783\,
            I => \c0.data_in_frame_19_5\
        );

    \I__13688\ : InMux
    port map (
            O => \N__58774\,
            I => \N__58771\
        );

    \I__13687\ : LocalMux
    port map (
            O => \N__58771\,
            I => \N__58767\
        );

    \I__13686\ : InMux
    port map (
            O => \N__58770\,
            I => \N__58763\
        );

    \I__13685\ : Span4Mux_h
    port map (
            O => \N__58767\,
            I => \N__58760\
        );

    \I__13684\ : InMux
    port map (
            O => \N__58766\,
            I => \N__58757\
        );

    \I__13683\ : LocalMux
    port map (
            O => \N__58763\,
            I => \N__58754\
        );

    \I__13682\ : Span4Mux_h
    port map (
            O => \N__58760\,
            I => \N__58751\
        );

    \I__13681\ : LocalMux
    port map (
            O => \N__58757\,
            I => \N__58746\
        );

    \I__13680\ : Span4Mux_v
    port map (
            O => \N__58754\,
            I => \N__58746\
        );

    \I__13679\ : Odrv4
    port map (
            O => \N__58751\,
            I => \c0.data_in_frame_26_1\
        );

    \I__13678\ : Odrv4
    port map (
            O => \N__58746\,
            I => \c0.data_in_frame_26_1\
        );

    \I__13677\ : InMux
    port map (
            O => \N__58741\,
            I => \N__58737\
        );

    \I__13676\ : InMux
    port map (
            O => \N__58740\,
            I => \N__58734\
        );

    \I__13675\ : LocalMux
    port map (
            O => \N__58737\,
            I => \c0.n21039\
        );

    \I__13674\ : LocalMux
    port map (
            O => \N__58734\,
            I => \c0.n21039\
        );

    \I__13673\ : CascadeMux
    port map (
            O => \N__58729\,
            I => \c0.n24_adj_4282_cascade_\
        );

    \I__13672\ : InMux
    port map (
            O => \N__58726\,
            I => \N__58723\
        );

    \I__13671\ : LocalMux
    port map (
            O => \N__58723\,
            I => \c0.n22711\
        );

    \I__13670\ : CascadeMux
    port map (
            O => \N__58720\,
            I => \c0.n22711_cascade_\
        );

    \I__13669\ : InMux
    port map (
            O => \N__58717\,
            I => \N__58714\
        );

    \I__13668\ : LocalMux
    port map (
            O => \N__58714\,
            I => \N__58709\
        );

    \I__13667\ : InMux
    port map (
            O => \N__58713\,
            I => \N__58706\
        );

    \I__13666\ : InMux
    port map (
            O => \N__58712\,
            I => \N__58703\
        );

    \I__13665\ : Odrv4
    port map (
            O => \N__58709\,
            I => \c0.n21200\
        );

    \I__13664\ : LocalMux
    port map (
            O => \N__58706\,
            I => \c0.n21200\
        );

    \I__13663\ : LocalMux
    port map (
            O => \N__58703\,
            I => \c0.n21200\
        );

    \I__13662\ : InMux
    port map (
            O => \N__58696\,
            I => \N__58693\
        );

    \I__13661\ : LocalMux
    port map (
            O => \N__58693\,
            I => \N__58688\
        );

    \I__13660\ : InMux
    port map (
            O => \N__58692\,
            I => \N__58685\
        );

    \I__13659\ : InMux
    port map (
            O => \N__58691\,
            I => \N__58682\
        );

    \I__13658\ : Odrv4
    port map (
            O => \N__58688\,
            I => \c0.n12596\
        );

    \I__13657\ : LocalMux
    port map (
            O => \N__58685\,
            I => \c0.n12596\
        );

    \I__13656\ : LocalMux
    port map (
            O => \N__58682\,
            I => \c0.n12596\
        );

    \I__13655\ : CascadeMux
    port map (
            O => \N__58675\,
            I => \N__58672\
        );

    \I__13654\ : InMux
    port map (
            O => \N__58672\,
            I => \N__58669\
        );

    \I__13653\ : LocalMux
    port map (
            O => \N__58669\,
            I => \N__58666\
        );

    \I__13652\ : Span12Mux_s10_h
    port map (
            O => \N__58666\,
            I => \N__58663\
        );

    \I__13651\ : Odrv12
    port map (
            O => \N__58663\,
            I => \c0.n6707\
        );

    \I__13650\ : CascadeMux
    port map (
            O => \N__58660\,
            I => \c0.n15_adj_4284_cascade_\
        );

    \I__13649\ : InMux
    port map (
            O => \N__58657\,
            I => \N__58654\
        );

    \I__13648\ : LocalMux
    port map (
            O => \N__58654\,
            I => \c0.n14_adj_4283\
        );

    \I__13647\ : InMux
    port map (
            O => \N__58651\,
            I => \N__58648\
        );

    \I__13646\ : LocalMux
    port map (
            O => \N__58648\,
            I => \c0.n22437\
        );

    \I__13645\ : InMux
    port map (
            O => \N__58645\,
            I => \N__58638\
        );

    \I__13644\ : InMux
    port map (
            O => \N__58644\,
            I => \N__58638\
        );

    \I__13643\ : InMux
    port map (
            O => \N__58643\,
            I => \N__58634\
        );

    \I__13642\ : LocalMux
    port map (
            O => \N__58638\,
            I => \N__58631\
        );

    \I__13641\ : InMux
    port map (
            O => \N__58637\,
            I => \N__58628\
        );

    \I__13640\ : LocalMux
    port map (
            O => \N__58634\,
            I => \N__58623\
        );

    \I__13639\ : Sp12to4
    port map (
            O => \N__58631\,
            I => \N__58623\
        );

    \I__13638\ : LocalMux
    port map (
            O => \N__58628\,
            I => \c0.data_in_frame_25_0\
        );

    \I__13637\ : Odrv12
    port map (
            O => \N__58623\,
            I => \c0.data_in_frame_25_0\
        );

    \I__13636\ : InMux
    port map (
            O => \N__58618\,
            I => \N__58615\
        );

    \I__13635\ : LocalMux
    port map (
            O => \N__58615\,
            I => \N__58611\
        );

    \I__13634\ : InMux
    port map (
            O => \N__58614\,
            I => \N__58606\
        );

    \I__13633\ : Span4Mux_v
    port map (
            O => \N__58611\,
            I => \N__58603\
        );

    \I__13632\ : CascadeMux
    port map (
            O => \N__58610\,
            I => \N__58600\
        );

    \I__13631\ : InMux
    port map (
            O => \N__58609\,
            I => \N__58597\
        );

    \I__13630\ : LocalMux
    port map (
            O => \N__58606\,
            I => \N__58594\
        );

    \I__13629\ : Span4Mux_h
    port map (
            O => \N__58603\,
            I => \N__58591\
        );

    \I__13628\ : InMux
    port map (
            O => \N__58600\,
            I => \N__58588\
        );

    \I__13627\ : LocalMux
    port map (
            O => \N__58597\,
            I => \N__58583\
        );

    \I__13626\ : Span4Mux_v
    port map (
            O => \N__58594\,
            I => \N__58583\
        );

    \I__13625\ : Span4Mux_v
    port map (
            O => \N__58591\,
            I => \N__58580\
        );

    \I__13624\ : LocalMux
    port map (
            O => \N__58588\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13623\ : Odrv4
    port map (
            O => \N__58583\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13622\ : Odrv4
    port map (
            O => \N__58580\,
            I => \c0.data_in_frame_25_6\
        );

    \I__13621\ : CascadeMux
    port map (
            O => \N__58573\,
            I => \c0.n22437_cascade_\
        );

    \I__13620\ : CascadeMux
    port map (
            O => \N__58570\,
            I => \N__58567\
        );

    \I__13619\ : InMux
    port map (
            O => \N__58567\,
            I => \N__58564\
        );

    \I__13618\ : LocalMux
    port map (
            O => \N__58564\,
            I => \c0.n50_adj_4487\
        );

    \I__13617\ : InMux
    port map (
            O => \N__58561\,
            I => \N__58557\
        );

    \I__13616\ : InMux
    port map (
            O => \N__58560\,
            I => \N__58554\
        );

    \I__13615\ : LocalMux
    port map (
            O => \N__58557\,
            I => \N__58551\
        );

    \I__13614\ : LocalMux
    port map (
            O => \N__58554\,
            I => \N__58548\
        );

    \I__13613\ : Odrv12
    port map (
            O => \N__58551\,
            I => \c0.n22323\
        );

    \I__13612\ : Odrv4
    port map (
            O => \N__58548\,
            I => \c0.n22323\
        );

    \I__13611\ : InMux
    port map (
            O => \N__58543\,
            I => \N__58536\
        );

    \I__13610\ : InMux
    port map (
            O => \N__58542\,
            I => \N__58536\
        );

    \I__13609\ : InMux
    port map (
            O => \N__58541\,
            I => \N__58533\
        );

    \I__13608\ : LocalMux
    port map (
            O => \N__58536\,
            I => \c0.n20203\
        );

    \I__13607\ : LocalMux
    port map (
            O => \N__58533\,
            I => \c0.n20203\
        );

    \I__13606\ : InMux
    port map (
            O => \N__58528\,
            I => \N__58525\
        );

    \I__13605\ : LocalMux
    port map (
            O => \N__58525\,
            I => \N__58522\
        );

    \I__13604\ : Span4Mux_v
    port map (
            O => \N__58522\,
            I => \N__58519\
        );

    \I__13603\ : Odrv4
    port map (
            O => \N__58519\,
            I => \c0.n21870\
        );

    \I__13602\ : CascadeMux
    port map (
            O => \N__58516\,
            I => \c0.n18_adj_4249_cascade_\
        );

    \I__13601\ : InMux
    port map (
            O => \N__58513\,
            I => \N__58510\
        );

    \I__13600\ : LocalMux
    port map (
            O => \N__58510\,
            I => \N__58507\
        );

    \I__13599\ : Odrv4
    port map (
            O => \N__58507\,
            I => \c0.n24_adj_4248\
        );

    \I__13598\ : InMux
    port map (
            O => \N__58504\,
            I => \N__58501\
        );

    \I__13597\ : LocalMux
    port map (
            O => \N__58501\,
            I => \c0.n26_adj_4250\
        );

    \I__13596\ : CascadeMux
    port map (
            O => \N__58498\,
            I => \N__58494\
        );

    \I__13595\ : InMux
    port map (
            O => \N__58497\,
            I => \N__58491\
        );

    \I__13594\ : InMux
    port map (
            O => \N__58494\,
            I => \N__58487\
        );

    \I__13593\ : LocalMux
    port map (
            O => \N__58491\,
            I => \N__58484\
        );

    \I__13592\ : InMux
    port map (
            O => \N__58490\,
            I => \N__58480\
        );

    \I__13591\ : LocalMux
    port map (
            O => \N__58487\,
            I => \N__58475\
        );

    \I__13590\ : Span4Mux_h
    port map (
            O => \N__58484\,
            I => \N__58475\
        );

    \I__13589\ : InMux
    port map (
            O => \N__58483\,
            I => \N__58472\
        );

    \I__13588\ : LocalMux
    port map (
            O => \N__58480\,
            I => \N__58469\
        );

    \I__13587\ : Span4Mux_v
    port map (
            O => \N__58475\,
            I => \N__58466\
        );

    \I__13586\ : LocalMux
    port map (
            O => \N__58472\,
            I => \c0.data_in_frame_15_4\
        );

    \I__13585\ : Odrv4
    port map (
            O => \N__58469\,
            I => \c0.data_in_frame_15_4\
        );

    \I__13584\ : Odrv4
    port map (
            O => \N__58466\,
            I => \c0.data_in_frame_15_4\
        );

    \I__13583\ : InMux
    port map (
            O => \N__58459\,
            I => \N__58455\
        );

    \I__13582\ : InMux
    port map (
            O => \N__58458\,
            I => \N__58452\
        );

    \I__13581\ : LocalMux
    port map (
            O => \N__58455\,
            I => \c0.n23072\
        );

    \I__13580\ : LocalMux
    port map (
            O => \N__58452\,
            I => \c0.n23072\
        );

    \I__13579\ : InMux
    port map (
            O => \N__58447\,
            I => \N__58441\
        );

    \I__13578\ : InMux
    port map (
            O => \N__58446\,
            I => \N__58441\
        );

    \I__13577\ : LocalMux
    port map (
            O => \N__58441\,
            I => \N__58438\
        );

    \I__13576\ : Span4Mux_h
    port map (
            O => \N__58438\,
            I => \N__58435\
        );

    \I__13575\ : Odrv4
    port map (
            O => \N__58435\,
            I => \c0.n13457\
        );

    \I__13574\ : CascadeMux
    port map (
            O => \N__58432\,
            I => \c0.n23072_cascade_\
        );

    \I__13573\ : InMux
    port map (
            O => \N__58429\,
            I => \N__58423\
        );

    \I__13572\ : InMux
    port map (
            O => \N__58428\,
            I => \N__58420\
        );

    \I__13571\ : InMux
    port map (
            O => \N__58427\,
            I => \N__58417\
        );

    \I__13570\ : InMux
    port map (
            O => \N__58426\,
            I => \N__58414\
        );

    \I__13569\ : LocalMux
    port map (
            O => \N__58423\,
            I => \N__58409\
        );

    \I__13568\ : LocalMux
    port map (
            O => \N__58420\,
            I => \N__58409\
        );

    \I__13567\ : LocalMux
    port map (
            O => \N__58417\,
            I => \N__58404\
        );

    \I__13566\ : LocalMux
    port map (
            O => \N__58414\,
            I => \N__58404\
        );

    \I__13565\ : Span4Mux_v
    port map (
            O => \N__58409\,
            I => \N__58401\
        );

    \I__13564\ : Odrv12
    port map (
            O => \N__58404\,
            I => \c0.n21067\
        );

    \I__13563\ : Odrv4
    port map (
            O => \N__58401\,
            I => \c0.n21067\
        );

    \I__13562\ : InMux
    port map (
            O => \N__58396\,
            I => \N__58393\
        );

    \I__13561\ : LocalMux
    port map (
            O => \N__58393\,
            I => \c0.n14_adj_4251\
        );

    \I__13560\ : InMux
    port map (
            O => \N__58390\,
            I => \N__58387\
        );

    \I__13559\ : LocalMux
    port map (
            O => \N__58387\,
            I => \c0.n21054\
        );

    \I__13558\ : CascadeMux
    port map (
            O => \N__58384\,
            I => \c0.n6_adj_4292_cascade_\
        );

    \I__13557\ : InMux
    port map (
            O => \N__58381\,
            I => \N__58378\
        );

    \I__13556\ : LocalMux
    port map (
            O => \N__58378\,
            I => \N__58374\
        );

    \I__13555\ : CascadeMux
    port map (
            O => \N__58377\,
            I => \N__58371\
        );

    \I__13554\ : Span4Mux_v
    port map (
            O => \N__58374\,
            I => \N__58368\
        );

    \I__13553\ : InMux
    port map (
            O => \N__58371\,
            I => \N__58365\
        );

    \I__13552\ : Span4Mux_h
    port map (
            O => \N__58368\,
            I => \N__58362\
        );

    \I__13551\ : LocalMux
    port map (
            O => \N__58365\,
            I => \c0.data_in_frame_28_5\
        );

    \I__13550\ : Odrv4
    port map (
            O => \N__58362\,
            I => \c0.data_in_frame_28_5\
        );

    \I__13549\ : InMux
    port map (
            O => \N__58357\,
            I => \N__58354\
        );

    \I__13548\ : LocalMux
    port map (
            O => \N__58354\,
            I => \N__58351\
        );

    \I__13547\ : Span4Mux_v
    port map (
            O => \N__58351\,
            I => \N__58348\
        );

    \I__13546\ : Span4Mux_h
    port map (
            O => \N__58348\,
            I => \N__58345\
        );

    \I__13545\ : Odrv4
    port map (
            O => \N__58345\,
            I => \c0.n23073\
        );

    \I__13544\ : InMux
    port map (
            O => \N__58342\,
            I => \N__58338\
        );

    \I__13543\ : InMux
    port map (
            O => \N__58341\,
            I => \N__58334\
        );

    \I__13542\ : LocalMux
    port map (
            O => \N__58338\,
            I => \N__58331\
        );

    \I__13541\ : CascadeMux
    port map (
            O => \N__58337\,
            I => \N__58328\
        );

    \I__13540\ : LocalMux
    port map (
            O => \N__58334\,
            I => \N__58324\
        );

    \I__13539\ : Span4Mux_h
    port map (
            O => \N__58331\,
            I => \N__58321\
        );

    \I__13538\ : InMux
    port map (
            O => \N__58328\,
            I => \N__58318\
        );

    \I__13537\ : InMux
    port map (
            O => \N__58327\,
            I => \N__58315\
        );

    \I__13536\ : Span4Mux_h
    port map (
            O => \N__58324\,
            I => \N__58312\
        );

    \I__13535\ : Span4Mux_v
    port map (
            O => \N__58321\,
            I => \N__58309\
        );

    \I__13534\ : LocalMux
    port map (
            O => \N__58318\,
            I => \c0.data_in_frame_21_4\
        );

    \I__13533\ : LocalMux
    port map (
            O => \N__58315\,
            I => \c0.data_in_frame_21_4\
        );

    \I__13532\ : Odrv4
    port map (
            O => \N__58312\,
            I => \c0.data_in_frame_21_4\
        );

    \I__13531\ : Odrv4
    port map (
            O => \N__58309\,
            I => \c0.data_in_frame_21_4\
        );

    \I__13530\ : InMux
    port map (
            O => \N__58300\,
            I => \N__58297\
        );

    \I__13529\ : LocalMux
    port map (
            O => \N__58297\,
            I => \c0.n21905\
        );

    \I__13528\ : CascadeMux
    port map (
            O => \N__58294\,
            I => \c0.n21905_cascade_\
        );

    \I__13527\ : InMux
    port map (
            O => \N__58291\,
            I => \N__58288\
        );

    \I__13526\ : LocalMux
    port map (
            O => \N__58288\,
            I => \N__58285\
        );

    \I__13525\ : Span12Mux_v
    port map (
            O => \N__58285\,
            I => \N__58282\
        );

    \I__13524\ : Odrv12
    port map (
            O => \N__58282\,
            I => \c0.n21069\
        );

    \I__13523\ : InMux
    port map (
            O => \N__58279\,
            I => \N__58275\
        );

    \I__13522\ : InMux
    port map (
            O => \N__58278\,
            I => \N__58272\
        );

    \I__13521\ : LocalMux
    port map (
            O => \N__58275\,
            I => \N__58269\
        );

    \I__13520\ : LocalMux
    port map (
            O => \N__58272\,
            I => \N__58266\
        );

    \I__13519\ : Odrv4
    port map (
            O => \N__58269\,
            I => \c0.n22113\
        );

    \I__13518\ : Odrv4
    port map (
            O => \N__58266\,
            I => \c0.n22113\
        );

    \I__13517\ : CascadeMux
    port map (
            O => \N__58261\,
            I => \N__58258\
        );

    \I__13516\ : InMux
    port map (
            O => \N__58258\,
            I => \N__58253\
        );

    \I__13515\ : InMux
    port map (
            O => \N__58257\,
            I => \N__58248\
        );

    \I__13514\ : InMux
    port map (
            O => \N__58256\,
            I => \N__58248\
        );

    \I__13513\ : LocalMux
    port map (
            O => \N__58253\,
            I => \c0.data_in_frame_20_3\
        );

    \I__13512\ : LocalMux
    port map (
            O => \N__58248\,
            I => \c0.data_in_frame_20_3\
        );

    \I__13511\ : InMux
    port map (
            O => \N__58243\,
            I => \N__58240\
        );

    \I__13510\ : LocalMux
    port map (
            O => \N__58240\,
            I => \c0.n22352\
        );

    \I__13509\ : CascadeMux
    port map (
            O => \N__58237\,
            I => \N__58233\
        );

    \I__13508\ : CascadeMux
    port map (
            O => \N__58236\,
            I => \N__58230\
        );

    \I__13507\ : InMux
    port map (
            O => \N__58233\,
            I => \N__58227\
        );

    \I__13506\ : InMux
    port map (
            O => \N__58230\,
            I => \N__58224\
        );

    \I__13505\ : LocalMux
    port map (
            O => \N__58227\,
            I => \N__58221\
        );

    \I__13504\ : LocalMux
    port map (
            O => \N__58224\,
            I => \c0.data_in_frame_18_4\
        );

    \I__13503\ : Odrv4
    port map (
            O => \N__58221\,
            I => \c0.data_in_frame_18_4\
        );

    \I__13502\ : InMux
    port map (
            O => \N__58216\,
            I => \N__58213\
        );

    \I__13501\ : LocalMux
    port map (
            O => \N__58213\,
            I => \N__58209\
        );

    \I__13500\ : InMux
    port map (
            O => \N__58212\,
            I => \N__58206\
        );

    \I__13499\ : Span4Mux_h
    port map (
            O => \N__58209\,
            I => \N__58200\
        );

    \I__13498\ : LocalMux
    port map (
            O => \N__58206\,
            I => \N__58200\
        );

    \I__13497\ : InMux
    port map (
            O => \N__58205\,
            I => \N__58197\
        );

    \I__13496\ : Span4Mux_v
    port map (
            O => \N__58200\,
            I => \N__58194\
        );

    \I__13495\ : LocalMux
    port map (
            O => \N__58197\,
            I => \c0.n13598\
        );

    \I__13494\ : Odrv4
    port map (
            O => \N__58194\,
            I => \c0.n13598\
        );

    \I__13493\ : InMux
    port map (
            O => \N__58189\,
            I => \N__58186\
        );

    \I__13492\ : LocalMux
    port map (
            O => \N__58186\,
            I => \N__58182\
        );

    \I__13491\ : InMux
    port map (
            O => \N__58185\,
            I => \N__58179\
        );

    \I__13490\ : Odrv12
    port map (
            O => \N__58182\,
            I => \c0.n20374\
        );

    \I__13489\ : LocalMux
    port map (
            O => \N__58179\,
            I => \c0.n20374\
        );

    \I__13488\ : CascadeMux
    port map (
            O => \N__58174\,
            I => \N__58169\
        );

    \I__13487\ : CascadeMux
    port map (
            O => \N__58173\,
            I => \N__58166\
        );

    \I__13486\ : InMux
    port map (
            O => \N__58172\,
            I => \N__58163\
        );

    \I__13485\ : InMux
    port map (
            O => \N__58169\,
            I => \N__58159\
        );

    \I__13484\ : InMux
    port map (
            O => \N__58166\,
            I => \N__58156\
        );

    \I__13483\ : LocalMux
    port map (
            O => \N__58163\,
            I => \N__58153\
        );

    \I__13482\ : InMux
    port map (
            O => \N__58162\,
            I => \N__58150\
        );

    \I__13481\ : LocalMux
    port map (
            O => \N__58159\,
            I => \c0.data_in_frame_16_5\
        );

    \I__13480\ : LocalMux
    port map (
            O => \N__58156\,
            I => \c0.data_in_frame_16_5\
        );

    \I__13479\ : Odrv4
    port map (
            O => \N__58153\,
            I => \c0.data_in_frame_16_5\
        );

    \I__13478\ : LocalMux
    port map (
            O => \N__58150\,
            I => \c0.data_in_frame_16_5\
        );

    \I__13477\ : InMux
    port map (
            O => \N__58141\,
            I => \N__58138\
        );

    \I__13476\ : LocalMux
    port map (
            O => \N__58138\,
            I => \N__58134\
        );

    \I__13475\ : InMux
    port map (
            O => \N__58137\,
            I => \N__58131\
        );

    \I__13474\ : Span4Mux_v
    port map (
            O => \N__58134\,
            I => \N__58127\
        );

    \I__13473\ : LocalMux
    port map (
            O => \N__58131\,
            I => \N__58124\
        );

    \I__13472\ : CascadeMux
    port map (
            O => \N__58130\,
            I => \N__58121\
        );

    \I__13471\ : Span4Mux_v
    port map (
            O => \N__58127\,
            I => \N__58118\
        );

    \I__13470\ : Span4Mux_h
    port map (
            O => \N__58124\,
            I => \N__58115\
        );

    \I__13469\ : InMux
    port map (
            O => \N__58121\,
            I => \N__58112\
        );

    \I__13468\ : Span4Mux_h
    port map (
            O => \N__58118\,
            I => \N__58109\
        );

    \I__13467\ : Span4Mux_h
    port map (
            O => \N__58115\,
            I => \N__58106\
        );

    \I__13466\ : LocalMux
    port map (
            O => \N__58112\,
            I => \c0.data_in_frame_16_3\
        );

    \I__13465\ : Odrv4
    port map (
            O => \N__58109\,
            I => \c0.data_in_frame_16_3\
        );

    \I__13464\ : Odrv4
    port map (
            O => \N__58106\,
            I => \c0.data_in_frame_16_3\
        );

    \I__13463\ : CascadeMux
    port map (
            O => \N__58099\,
            I => \N__58095\
        );

    \I__13462\ : InMux
    port map (
            O => \N__58098\,
            I => \N__58091\
        );

    \I__13461\ : InMux
    port map (
            O => \N__58095\,
            I => \N__58088\
        );

    \I__13460\ : InMux
    port map (
            O => \N__58094\,
            I => \N__58085\
        );

    \I__13459\ : LocalMux
    port map (
            O => \N__58091\,
            I => \N__58082\
        );

    \I__13458\ : LocalMux
    port map (
            O => \N__58088\,
            I => \c0.data_in_frame_16_2\
        );

    \I__13457\ : LocalMux
    port map (
            O => \N__58085\,
            I => \c0.data_in_frame_16_2\
        );

    \I__13456\ : Odrv4
    port map (
            O => \N__58082\,
            I => \c0.data_in_frame_16_2\
        );

    \I__13455\ : InMux
    port map (
            O => \N__58075\,
            I => \N__58072\
        );

    \I__13454\ : LocalMux
    port map (
            O => \N__58072\,
            I => \c0.n10_adj_4230\
        );

    \I__13453\ : CascadeMux
    port map (
            O => \N__58069\,
            I => \N__58064\
        );

    \I__13452\ : InMux
    port map (
            O => \N__58068\,
            I => \N__58056\
        );

    \I__13451\ : InMux
    port map (
            O => \N__58067\,
            I => \N__58056\
        );

    \I__13450\ : InMux
    port map (
            O => \N__58064\,
            I => \N__58051\
        );

    \I__13449\ : InMux
    port map (
            O => \N__58063\,
            I => \N__58051\
        );

    \I__13448\ : InMux
    port map (
            O => \N__58062\,
            I => \N__58046\
        );

    \I__13447\ : InMux
    port map (
            O => \N__58061\,
            I => \N__58046\
        );

    \I__13446\ : LocalMux
    port map (
            O => \N__58056\,
            I => \N__58043\
        );

    \I__13445\ : LocalMux
    port map (
            O => \N__58051\,
            I => \c0.data_in_frame_13_4\
        );

    \I__13444\ : LocalMux
    port map (
            O => \N__58046\,
            I => \c0.data_in_frame_13_4\
        );

    \I__13443\ : Odrv12
    port map (
            O => \N__58043\,
            I => \c0.data_in_frame_13_4\
        );

    \I__13442\ : CascadeMux
    port map (
            O => \N__58036\,
            I => \N__58033\
        );

    \I__13441\ : InMux
    port map (
            O => \N__58033\,
            I => \N__58030\
        );

    \I__13440\ : LocalMux
    port map (
            O => \N__58030\,
            I => \N__58025\
        );

    \I__13439\ : InMux
    port map (
            O => \N__58029\,
            I => \N__58022\
        );

    \I__13438\ : CascadeMux
    port map (
            O => \N__58028\,
            I => \N__58019\
        );

    \I__13437\ : Span4Mux_v
    port map (
            O => \N__58025\,
            I => \N__58013\
        );

    \I__13436\ : LocalMux
    port map (
            O => \N__58022\,
            I => \N__58013\
        );

    \I__13435\ : InMux
    port map (
            O => \N__58019\,
            I => \N__58010\
        );

    \I__13434\ : InMux
    port map (
            O => \N__58018\,
            I => \N__58007\
        );

    \I__13433\ : Span4Mux_h
    port map (
            O => \N__58013\,
            I => \N__58004\
        );

    \I__13432\ : LocalMux
    port map (
            O => \N__58010\,
            I => \c0.data_in_frame_15_5\
        );

    \I__13431\ : LocalMux
    port map (
            O => \N__58007\,
            I => \c0.data_in_frame_15_5\
        );

    \I__13430\ : Odrv4
    port map (
            O => \N__58004\,
            I => \c0.data_in_frame_15_5\
        );

    \I__13429\ : CascadeMux
    port map (
            O => \N__57997\,
            I => \N__57994\
        );

    \I__13428\ : InMux
    port map (
            O => \N__57994\,
            I => \N__57991\
        );

    \I__13427\ : LocalMux
    port map (
            O => \N__57991\,
            I => \N__57988\
        );

    \I__13426\ : Span4Mux_v
    port map (
            O => \N__57988\,
            I => \N__57984\
        );

    \I__13425\ : InMux
    port map (
            O => \N__57987\,
            I => \N__57981\
        );

    \I__13424\ : Span4Mux_h
    port map (
            O => \N__57984\,
            I => \N__57978\
        );

    \I__13423\ : LocalMux
    port map (
            O => \N__57981\,
            I => \c0.data_in_frame_26_3\
        );

    \I__13422\ : Odrv4
    port map (
            O => \N__57978\,
            I => \c0.data_in_frame_26_3\
        );

    \I__13421\ : InMux
    port map (
            O => \N__57973\,
            I => \N__57969\
        );

    \I__13420\ : CascadeMux
    port map (
            O => \N__57972\,
            I => \N__57966\
        );

    \I__13419\ : LocalMux
    port map (
            O => \N__57969\,
            I => \N__57963\
        );

    \I__13418\ : InMux
    port map (
            O => \N__57966\,
            I => \N__57960\
        );

    \I__13417\ : Odrv4
    port map (
            O => \N__57963\,
            I => \c0.n20266\
        );

    \I__13416\ : LocalMux
    port map (
            O => \N__57960\,
            I => \c0.n20266\
        );

    \I__13415\ : CascadeMux
    port map (
            O => \N__57955\,
            I => \c0.n22402_cascade_\
        );

    \I__13414\ : InMux
    port map (
            O => \N__57952\,
            I => \N__57949\
        );

    \I__13413\ : LocalMux
    port map (
            O => \N__57949\,
            I => \N__57946\
        );

    \I__13412\ : Span4Mux_v
    port map (
            O => \N__57946\,
            I => \N__57943\
        );

    \I__13411\ : Odrv4
    port map (
            O => \N__57943\,
            I => \c0.n33\
        );

    \I__13410\ : InMux
    port map (
            O => \N__57940\,
            I => \N__57937\
        );

    \I__13409\ : LocalMux
    port map (
            O => \N__57937\,
            I => \N__57933\
        );

    \I__13408\ : InMux
    port map (
            O => \N__57936\,
            I => \N__57930\
        );

    \I__13407\ : Odrv4
    port map (
            O => \N__57933\,
            I => \c0.n21982\
        );

    \I__13406\ : LocalMux
    port map (
            O => \N__57930\,
            I => \c0.n21982\
        );

    \I__13405\ : InMux
    port map (
            O => \N__57925\,
            I => \N__57921\
        );

    \I__13404\ : InMux
    port map (
            O => \N__57924\,
            I => \N__57918\
        );

    \I__13403\ : LocalMux
    port map (
            O => \N__57921\,
            I => \N__57915\
        );

    \I__13402\ : LocalMux
    port map (
            O => \N__57918\,
            I => data_in_frame_14_0
        );

    \I__13401\ : Odrv12
    port map (
            O => \N__57915\,
            I => data_in_frame_14_0
        );

    \I__13400\ : InMux
    port map (
            O => \N__57910\,
            I => \N__57905\
        );

    \I__13399\ : InMux
    port map (
            O => \N__57909\,
            I => \N__57902\
        );

    \I__13398\ : InMux
    port map (
            O => \N__57908\,
            I => \N__57899\
        );

    \I__13397\ : LocalMux
    port map (
            O => \N__57905\,
            I => \N__57896\
        );

    \I__13396\ : LocalMux
    port map (
            O => \N__57902\,
            I => \N__57893\
        );

    \I__13395\ : LocalMux
    port map (
            O => \N__57899\,
            I => \N__57890\
        );

    \I__13394\ : Span4Mux_h
    port map (
            O => \N__57896\,
            I => \N__57882\
        );

    \I__13393\ : Span4Mux_v
    port map (
            O => \N__57893\,
            I => \N__57882\
        );

    \I__13392\ : Span4Mux_v
    port map (
            O => \N__57890\,
            I => \N__57882\
        );

    \I__13391\ : InMux
    port map (
            O => \N__57889\,
            I => \N__57879\
        );

    \I__13390\ : Odrv4
    port map (
            O => \N__57882\,
            I => \c0.n13865\
        );

    \I__13389\ : LocalMux
    port map (
            O => \N__57879\,
            I => \c0.n13865\
        );

    \I__13388\ : InMux
    port map (
            O => \N__57874\,
            I => \N__57871\
        );

    \I__13387\ : LocalMux
    port map (
            O => \N__57871\,
            I => \N__57866\
        );

    \I__13386\ : InMux
    port map (
            O => \N__57870\,
            I => \N__57863\
        );

    \I__13385\ : InMux
    port map (
            O => \N__57869\,
            I => \N__57860\
        );

    \I__13384\ : Span4Mux_v
    port map (
            O => \N__57866\,
            I => \N__57857\
        );

    \I__13383\ : LocalMux
    port map (
            O => \N__57863\,
            I => \c0.data_in_frame_15_6\
        );

    \I__13382\ : LocalMux
    port map (
            O => \N__57860\,
            I => \c0.data_in_frame_15_6\
        );

    \I__13381\ : Odrv4
    port map (
            O => \N__57857\,
            I => \c0.data_in_frame_15_6\
        );

    \I__13380\ : InMux
    port map (
            O => \N__57850\,
            I => \N__57844\
        );

    \I__13379\ : InMux
    port map (
            O => \N__57849\,
            I => \N__57844\
        );

    \I__13378\ : LocalMux
    port map (
            O => \N__57844\,
            I => \N__57839\
        );

    \I__13377\ : InMux
    port map (
            O => \N__57843\,
            I => \N__57834\
        );

    \I__13376\ : InMux
    port map (
            O => \N__57842\,
            I => \N__57834\
        );

    \I__13375\ : Odrv4
    port map (
            O => \N__57839\,
            I => \c0.n4_adj_4240\
        );

    \I__13374\ : LocalMux
    port map (
            O => \N__57834\,
            I => \c0.n4_adj_4240\
        );

    \I__13373\ : CascadeMux
    port map (
            O => \N__57829\,
            I => \c0.n22352_cascade_\
        );

    \I__13372\ : CascadeMux
    port map (
            O => \N__57826\,
            I => \c0.n22000_cascade_\
        );

    \I__13371\ : InMux
    port map (
            O => \N__57823\,
            I => \N__57820\
        );

    \I__13370\ : LocalMux
    port map (
            O => \N__57820\,
            I => \c0.n31\
        );

    \I__13369\ : InMux
    port map (
            O => \N__57817\,
            I => \N__57814\
        );

    \I__13368\ : LocalMux
    port map (
            O => \N__57814\,
            I => \N__57811\
        );

    \I__13367\ : Span4Mux_h
    port map (
            O => \N__57811\,
            I => \N__57806\
        );

    \I__13366\ : InMux
    port map (
            O => \N__57810\,
            I => \N__57801\
        );

    \I__13365\ : InMux
    port map (
            O => \N__57809\,
            I => \N__57801\
        );

    \I__13364\ : Odrv4
    port map (
            O => \N__57806\,
            I => \c0.data_in_frame_15_7\
        );

    \I__13363\ : LocalMux
    port map (
            O => \N__57801\,
            I => \c0.data_in_frame_15_7\
        );

    \I__13362\ : CascadeMux
    port map (
            O => \N__57796\,
            I => \N__57792\
        );

    \I__13361\ : CascadeMux
    port map (
            O => \N__57795\,
            I => \N__57789\
        );

    \I__13360\ : InMux
    port map (
            O => \N__57792\,
            I => \N__57786\
        );

    \I__13359\ : InMux
    port map (
            O => \N__57789\,
            I => \N__57783\
        );

    \I__13358\ : LocalMux
    port map (
            O => \N__57786\,
            I => \c0.data_in_frame_18_2\
        );

    \I__13357\ : LocalMux
    port map (
            O => \N__57783\,
            I => \c0.data_in_frame_18_2\
        );

    \I__13356\ : InMux
    port map (
            O => \N__57778\,
            I => \N__57775\
        );

    \I__13355\ : LocalMux
    port map (
            O => \N__57775\,
            I => \N__57772\
        );

    \I__13354\ : Odrv4
    port map (
            O => \N__57772\,
            I => \c0.n22000\
        );

    \I__13353\ : CascadeMux
    port map (
            O => \N__57769\,
            I => \c0.n12_cascade_\
        );

    \I__13352\ : InMux
    port map (
            O => \N__57766\,
            I => \N__57763\
        );

    \I__13351\ : LocalMux
    port map (
            O => \N__57763\,
            I => \N__57760\
        );

    \I__13350\ : Odrv12
    port map (
            O => \N__57760\,
            I => \c0.n10_adj_4239\
        );

    \I__13349\ : CascadeMux
    port map (
            O => \N__57757\,
            I => \N__57753\
        );

    \I__13348\ : InMux
    port map (
            O => \N__57756\,
            I => \N__57750\
        );

    \I__13347\ : InMux
    port map (
            O => \N__57753\,
            I => \N__57747\
        );

    \I__13346\ : LocalMux
    port map (
            O => \N__57750\,
            I => \c0.data_in_frame_18_0\
        );

    \I__13345\ : LocalMux
    port map (
            O => \N__57747\,
            I => \c0.data_in_frame_18_0\
        );

    \I__13344\ : InMux
    port map (
            O => \N__57742\,
            I => \N__57739\
        );

    \I__13343\ : LocalMux
    port map (
            O => \N__57739\,
            I => \c0.n14_adj_4238\
        );

    \I__13342\ : CascadeMux
    port map (
            O => \N__57736\,
            I => \c0.n13210_cascade_\
        );

    \I__13341\ : InMux
    port map (
            O => \N__57733\,
            I => \N__57727\
        );

    \I__13340\ : InMux
    port map (
            O => \N__57732\,
            I => \N__57724\
        );

    \I__13339\ : CascadeMux
    port map (
            O => \N__57731\,
            I => \N__57721\
        );

    \I__13338\ : InMux
    port map (
            O => \N__57730\,
            I => \N__57718\
        );

    \I__13337\ : LocalMux
    port map (
            O => \N__57727\,
            I => \N__57713\
        );

    \I__13336\ : LocalMux
    port map (
            O => \N__57724\,
            I => \N__57713\
        );

    \I__13335\ : InMux
    port map (
            O => \N__57721\,
            I => \N__57709\
        );

    \I__13334\ : LocalMux
    port map (
            O => \N__57718\,
            I => \N__57706\
        );

    \I__13333\ : Span4Mux_h
    port map (
            O => \N__57713\,
            I => \N__57703\
        );

    \I__13332\ : InMux
    port map (
            O => \N__57712\,
            I => \N__57700\
        );

    \I__13331\ : LocalMux
    port map (
            O => \N__57709\,
            I => \c0.data_in_frame_8_7\
        );

    \I__13330\ : Odrv12
    port map (
            O => \N__57706\,
            I => \c0.data_in_frame_8_7\
        );

    \I__13329\ : Odrv4
    port map (
            O => \N__57703\,
            I => \c0.data_in_frame_8_7\
        );

    \I__13328\ : LocalMux
    port map (
            O => \N__57700\,
            I => \c0.data_in_frame_8_7\
        );

    \I__13327\ : InMux
    port map (
            O => \N__57691\,
            I => \N__57688\
        );

    \I__13326\ : LocalMux
    port map (
            O => \N__57688\,
            I => \N__57685\
        );

    \I__13325\ : Odrv4
    port map (
            O => \N__57685\,
            I => \c0.n21822\
        );

    \I__13324\ : CascadeMux
    port map (
            O => \N__57682\,
            I => \c0.n7_adj_4277_cascade_\
        );

    \I__13323\ : CascadeMux
    port map (
            O => \N__57679\,
            I => \N__57676\
        );

    \I__13322\ : InMux
    port map (
            O => \N__57676\,
            I => \N__57671\
        );

    \I__13321\ : InMux
    port map (
            O => \N__57675\,
            I => \N__57668\
        );

    \I__13320\ : InMux
    port map (
            O => \N__57674\,
            I => \N__57665\
        );

    \I__13319\ : LocalMux
    port map (
            O => \N__57671\,
            I => \c0.data_in_frame_11_5\
        );

    \I__13318\ : LocalMux
    port map (
            O => \N__57668\,
            I => \c0.data_in_frame_11_5\
        );

    \I__13317\ : LocalMux
    port map (
            O => \N__57665\,
            I => \c0.data_in_frame_11_5\
        );

    \I__13316\ : CascadeMux
    port map (
            O => \N__57658\,
            I => \c0.n10_adj_4264_cascade_\
        );

    \I__13315\ : InMux
    port map (
            O => \N__57655\,
            I => \N__57652\
        );

    \I__13314\ : LocalMux
    port map (
            O => \N__57652\,
            I => \N__57649\
        );

    \I__13313\ : Span4Mux_h
    port map (
            O => \N__57649\,
            I => \N__57646\
        );

    \I__13312\ : Odrv4
    port map (
            O => \N__57646\,
            I => \c0.n16_adj_4265\
        );

    \I__13311\ : InMux
    port map (
            O => \N__57643\,
            I => \N__57640\
        );

    \I__13310\ : LocalMux
    port map (
            O => \N__57640\,
            I => \N__57636\
        );

    \I__13309\ : CascadeMux
    port map (
            O => \N__57639\,
            I => \N__57633\
        );

    \I__13308\ : Span4Mux_h
    port map (
            O => \N__57636\,
            I => \N__57629\
        );

    \I__13307\ : InMux
    port map (
            O => \N__57633\,
            I => \N__57624\
        );

    \I__13306\ : InMux
    port map (
            O => \N__57632\,
            I => \N__57624\
        );

    \I__13305\ : Odrv4
    port map (
            O => \N__57629\,
            I => \c0.data_in_frame_11_6\
        );

    \I__13304\ : LocalMux
    port map (
            O => \N__57624\,
            I => \c0.data_in_frame_11_6\
        );

    \I__13303\ : CascadeMux
    port map (
            O => \N__57619\,
            I => \N__57616\
        );

    \I__13302\ : InMux
    port map (
            O => \N__57616\,
            I => \N__57609\
        );

    \I__13301\ : InMux
    port map (
            O => \N__57615\,
            I => \N__57609\
        );

    \I__13300\ : CascadeMux
    port map (
            O => \N__57614\,
            I => \N__57606\
        );

    \I__13299\ : LocalMux
    port map (
            O => \N__57609\,
            I => \N__57602\
        );

    \I__13298\ : InMux
    port map (
            O => \N__57606\,
            I => \N__57597\
        );

    \I__13297\ : InMux
    port map (
            O => \N__57605\,
            I => \N__57597\
        );

    \I__13296\ : Odrv12
    port map (
            O => \N__57602\,
            I => \c0.data_in_frame_11_2\
        );

    \I__13295\ : LocalMux
    port map (
            O => \N__57597\,
            I => \c0.data_in_frame_11_2\
        );

    \I__13294\ : InMux
    port map (
            O => \N__57592\,
            I => \N__57589\
        );

    \I__13293\ : LocalMux
    port map (
            O => \N__57589\,
            I => \N__57586\
        );

    \I__13292\ : Span4Mux_h
    port map (
            O => \N__57586\,
            I => \N__57578\
        );

    \I__13291\ : InMux
    port map (
            O => \N__57585\,
            I => \N__57573\
        );

    \I__13290\ : InMux
    port map (
            O => \N__57584\,
            I => \N__57573\
        );

    \I__13289\ : InMux
    port map (
            O => \N__57583\,
            I => \N__57570\
        );

    \I__13288\ : InMux
    port map (
            O => \N__57582\,
            I => \N__57567\
        );

    \I__13287\ : InMux
    port map (
            O => \N__57581\,
            I => \N__57564\
        );

    \I__13286\ : Odrv4
    port map (
            O => \N__57578\,
            I => \c0.n20135\
        );

    \I__13285\ : LocalMux
    port map (
            O => \N__57573\,
            I => \c0.n20135\
        );

    \I__13284\ : LocalMux
    port map (
            O => \N__57570\,
            I => \c0.n20135\
        );

    \I__13283\ : LocalMux
    port map (
            O => \N__57567\,
            I => \c0.n20135\
        );

    \I__13282\ : LocalMux
    port map (
            O => \N__57564\,
            I => \c0.n20135\
        );

    \I__13281\ : CascadeMux
    port map (
            O => \N__57553\,
            I => \N__57550\
        );

    \I__13280\ : InMux
    port map (
            O => \N__57550\,
            I => \N__57547\
        );

    \I__13279\ : LocalMux
    port map (
            O => \N__57547\,
            I => \N__57544\
        );

    \I__13278\ : Odrv4
    port map (
            O => \N__57544\,
            I => \c0.n22464\
        );

    \I__13277\ : InMux
    port map (
            O => \N__57541\,
            I => \N__57537\
        );

    \I__13276\ : InMux
    port map (
            O => \N__57540\,
            I => \N__57534\
        );

    \I__13275\ : LocalMux
    port map (
            O => \N__57537\,
            I => \c0.n21867\
        );

    \I__13274\ : LocalMux
    port map (
            O => \N__57534\,
            I => \c0.n21867\
        );

    \I__13273\ : InMux
    port map (
            O => \N__57529\,
            I => \N__57526\
        );

    \I__13272\ : LocalMux
    port map (
            O => \N__57526\,
            I => \c0.n6_adj_4225\
        );

    \I__13271\ : InMux
    port map (
            O => \N__57523\,
            I => \N__57520\
        );

    \I__13270\ : LocalMux
    port map (
            O => \N__57520\,
            I => \N__57517\
        );

    \I__13269\ : Odrv4
    port map (
            O => \N__57517\,
            I => \c0.n15_adj_4269\
        );

    \I__13268\ : CascadeMux
    port map (
            O => \N__57514\,
            I => \c0.n22464_cascade_\
        );

    \I__13267\ : InMux
    port map (
            O => \N__57511\,
            I => \N__57508\
        );

    \I__13266\ : LocalMux
    port map (
            O => \N__57508\,
            I => \N__57505\
        );

    \I__13265\ : Span4Mux_h
    port map (
            O => \N__57505\,
            I => \N__57502\
        );

    \I__13264\ : Odrv4
    port map (
            O => \N__57502\,
            I => \c0.n22415\
        );

    \I__13263\ : InMux
    port map (
            O => \N__57499\,
            I => \N__57493\
        );

    \I__13262\ : InMux
    port map (
            O => \N__57498\,
            I => \N__57493\
        );

    \I__13261\ : LocalMux
    port map (
            O => \N__57493\,
            I => \c0.n13728\
        );

    \I__13260\ : InMux
    port map (
            O => \N__57490\,
            I => \N__57486\
        );

    \I__13259\ : InMux
    port map (
            O => \N__57489\,
            I => \N__57483\
        );

    \I__13258\ : LocalMux
    port map (
            O => \N__57486\,
            I => \N__57480\
        );

    \I__13257\ : LocalMux
    port map (
            O => \N__57483\,
            I => \N__57477\
        );

    \I__13256\ : Span4Mux_h
    port map (
            O => \N__57480\,
            I => \N__57472\
        );

    \I__13255\ : Span4Mux_v
    port map (
            O => \N__57477\,
            I => \N__57472\
        );

    \I__13254\ : Odrv4
    port map (
            O => \N__57472\,
            I => \c0.n14053\
        );

    \I__13253\ : CascadeMux
    port map (
            O => \N__57469\,
            I => \N__57465\
        );

    \I__13252\ : InMux
    port map (
            O => \N__57468\,
            I => \N__57462\
        );

    \I__13251\ : InMux
    port map (
            O => \N__57465\,
            I => \N__57459\
        );

    \I__13250\ : LocalMux
    port map (
            O => \N__57462\,
            I => \N__57456\
        );

    \I__13249\ : LocalMux
    port map (
            O => \N__57459\,
            I => \c0.data_in_frame_18_1\
        );

    \I__13248\ : Odrv4
    port map (
            O => \N__57456\,
            I => \c0.data_in_frame_18_1\
        );

    \I__13247\ : CascadeMux
    port map (
            O => \N__57451\,
            I => \c0.n14053_cascade_\
        );

    \I__13246\ : InMux
    port map (
            O => \N__57448\,
            I => \N__57441\
        );

    \I__13245\ : InMux
    port map (
            O => \N__57447\,
            I => \N__57438\
        );

    \I__13244\ : InMux
    port map (
            O => \N__57446\,
            I => \N__57433\
        );

    \I__13243\ : InMux
    port map (
            O => \N__57445\,
            I => \N__57433\
        );

    \I__13242\ : CascadeMux
    port map (
            O => \N__57444\,
            I => \N__57430\
        );

    \I__13241\ : LocalMux
    port map (
            O => \N__57441\,
            I => \N__57425\
        );

    \I__13240\ : LocalMux
    port map (
            O => \N__57438\,
            I => \N__57425\
        );

    \I__13239\ : LocalMux
    port map (
            O => \N__57433\,
            I => \N__57422\
        );

    \I__13238\ : InMux
    port map (
            O => \N__57430\,
            I => \N__57419\
        );

    \I__13237\ : Span12Mux_v
    port map (
            O => \N__57425\,
            I => \N__57416\
        );

    \I__13236\ : Span4Mux_h
    port map (
            O => \N__57422\,
            I => \N__57413\
        );

    \I__13235\ : LocalMux
    port map (
            O => \N__57419\,
            I => \c0.data_in_frame_17_7\
        );

    \I__13234\ : Odrv12
    port map (
            O => \N__57416\,
            I => \c0.data_in_frame_17_7\
        );

    \I__13233\ : Odrv4
    port map (
            O => \N__57413\,
            I => \c0.data_in_frame_17_7\
        );

    \I__13232\ : CascadeMux
    port map (
            O => \N__57406\,
            I => \c0.n23586_cascade_\
        );

    \I__13231\ : InMux
    port map (
            O => \N__57403\,
            I => \N__57400\
        );

    \I__13230\ : LocalMux
    port map (
            O => \N__57400\,
            I => \N__57397\
        );

    \I__13229\ : Span4Mux_h
    port map (
            O => \N__57397\,
            I => \N__57392\
        );

    \I__13228\ : InMux
    port map (
            O => \N__57396\,
            I => \N__57387\
        );

    \I__13227\ : InMux
    port map (
            O => \N__57395\,
            I => \N__57387\
        );

    \I__13226\ : Odrv4
    port map (
            O => \N__57392\,
            I => \c0.data_in_frame_9_3\
        );

    \I__13225\ : LocalMux
    port map (
            O => \N__57387\,
            I => \c0.data_in_frame_9_3\
        );

    \I__13224\ : InMux
    port map (
            O => \N__57382\,
            I => \N__57379\
        );

    \I__13223\ : LocalMux
    port map (
            O => \N__57379\,
            I => \N__57376\
        );

    \I__13222\ : Span4Mux_h
    port map (
            O => \N__57376\,
            I => \N__57373\
        );

    \I__13221\ : Odrv4
    port map (
            O => \N__57373\,
            I => \c0.n22043\
        );

    \I__13220\ : CascadeMux
    port map (
            O => \N__57370\,
            I => \N__57366\
        );

    \I__13219\ : InMux
    port map (
            O => \N__57369\,
            I => \N__57362\
        );

    \I__13218\ : InMux
    port map (
            O => \N__57366\,
            I => \N__57359\
        );

    \I__13217\ : InMux
    port map (
            O => \N__57365\,
            I => \N__57356\
        );

    \I__13216\ : LocalMux
    port map (
            O => \N__57362\,
            I => \N__57353\
        );

    \I__13215\ : LocalMux
    port map (
            O => \N__57359\,
            I => \c0.data_in_frame_9_7\
        );

    \I__13214\ : LocalMux
    port map (
            O => \N__57356\,
            I => \c0.data_in_frame_9_7\
        );

    \I__13213\ : Odrv4
    port map (
            O => \N__57353\,
            I => \c0.data_in_frame_9_7\
        );

    \I__13212\ : InMux
    port map (
            O => \N__57346\,
            I => \N__57342\
        );

    \I__13211\ : InMux
    port map (
            O => \N__57345\,
            I => \N__57339\
        );

    \I__13210\ : LocalMux
    port map (
            O => \N__57342\,
            I => \N__57336\
        );

    \I__13209\ : LocalMux
    port map (
            O => \N__57339\,
            I => \N__57333\
        );

    \I__13208\ : Span4Mux_v
    port map (
            O => \N__57336\,
            I => \N__57330\
        );

    \I__13207\ : Odrv4
    port map (
            O => \N__57333\,
            I => \c0.n22471\
        );

    \I__13206\ : Odrv4
    port map (
            O => \N__57330\,
            I => \c0.n22471\
        );

    \I__13205\ : InMux
    port map (
            O => \N__57325\,
            I => \N__57321\
        );

    \I__13204\ : CascadeMux
    port map (
            O => \N__57324\,
            I => \N__57318\
        );

    \I__13203\ : LocalMux
    port map (
            O => \N__57321\,
            I => \N__57315\
        );

    \I__13202\ : InMux
    port map (
            O => \N__57318\,
            I => \N__57310\
        );

    \I__13201\ : Span12Mux_v
    port map (
            O => \N__57315\,
            I => \N__57307\
        );

    \I__13200\ : InMux
    port map (
            O => \N__57314\,
            I => \N__57304\
        );

    \I__13199\ : InMux
    port map (
            O => \N__57313\,
            I => \N__57301\
        );

    \I__13198\ : LocalMux
    port map (
            O => \N__57310\,
            I => \c0.data_in_frame_16_4\
        );

    \I__13197\ : Odrv12
    port map (
            O => \N__57307\,
            I => \c0.data_in_frame_16_4\
        );

    \I__13196\ : LocalMux
    port map (
            O => \N__57304\,
            I => \c0.data_in_frame_16_4\
        );

    \I__13195\ : LocalMux
    port map (
            O => \N__57301\,
            I => \c0.data_in_frame_16_4\
        );

    \I__13194\ : InMux
    port map (
            O => \N__57292\,
            I => \N__57286\
        );

    \I__13193\ : InMux
    port map (
            O => \N__57291\,
            I => \N__57286\
        );

    \I__13192\ : LocalMux
    port map (
            O => \N__57286\,
            I => \N__57280\
        );

    \I__13191\ : InMux
    port map (
            O => \N__57285\,
            I => \N__57277\
        );

    \I__13190\ : InMux
    port map (
            O => \N__57284\,
            I => \N__57274\
        );

    \I__13189\ : InMux
    port map (
            O => \N__57283\,
            I => \N__57271\
        );

    \I__13188\ : Span4Mux_v
    port map (
            O => \N__57280\,
            I => \N__57266\
        );

    \I__13187\ : LocalMux
    port map (
            O => \N__57277\,
            I => \N__57266\
        );

    \I__13186\ : LocalMux
    port map (
            O => \N__57274\,
            I => \N__57263\
        );

    \I__13185\ : LocalMux
    port map (
            O => \N__57271\,
            I => \N__57258\
        );

    \I__13184\ : Span4Mux_v
    port map (
            O => \N__57266\,
            I => \N__57258\
        );

    \I__13183\ : Odrv12
    port map (
            O => \N__57263\,
            I => \c0.n20240\
        );

    \I__13182\ : Odrv4
    port map (
            O => \N__57258\,
            I => \c0.n20240\
        );

    \I__13181\ : CascadeMux
    port map (
            O => \N__57253\,
            I => \N__57250\
        );

    \I__13180\ : InMux
    port map (
            O => \N__57250\,
            I => \N__57247\
        );

    \I__13179\ : LocalMux
    port map (
            O => \N__57247\,
            I => \c0.n22446\
        );

    \I__13178\ : CascadeMux
    port map (
            O => \N__57244\,
            I => \N__57241\
        );

    \I__13177\ : InMux
    port map (
            O => \N__57241\,
            I => \N__57238\
        );

    \I__13176\ : LocalMux
    port map (
            O => \N__57238\,
            I => \N__57235\
        );

    \I__13175\ : Span4Mux_h
    port map (
            O => \N__57235\,
            I => \N__57231\
        );

    \I__13174\ : InMux
    port map (
            O => \N__57234\,
            I => \N__57228\
        );

    \I__13173\ : Span4Mux_v
    port map (
            O => \N__57231\,
            I => \N__57225\
        );

    \I__13172\ : LocalMux
    port map (
            O => \N__57228\,
            I => \c0.n22328\
        );

    \I__13171\ : Odrv4
    port map (
            O => \N__57225\,
            I => \c0.n22328\
        );

    \I__13170\ : CascadeMux
    port map (
            O => \N__57220\,
            I => \c0.n22446_cascade_\
        );

    \I__13169\ : InMux
    port map (
            O => \N__57217\,
            I => \N__57213\
        );

    \I__13168\ : InMux
    port map (
            O => \N__57216\,
            I => \N__57210\
        );

    \I__13167\ : LocalMux
    port map (
            O => \N__57213\,
            I => \N__57207\
        );

    \I__13166\ : LocalMux
    port map (
            O => \N__57210\,
            I => \N__57204\
        );

    \I__13165\ : Odrv4
    port map (
            O => \N__57207\,
            I => \c0.n22424\
        );

    \I__13164\ : Odrv4
    port map (
            O => \N__57204\,
            I => \c0.n22424\
        );

    \I__13163\ : InMux
    port map (
            O => \N__57199\,
            I => \N__57196\
        );

    \I__13162\ : LocalMux
    port map (
            O => \N__57196\,
            I => \N__57193\
        );

    \I__13161\ : Span4Mux_v
    port map (
            O => \N__57193\,
            I => \N__57190\
        );

    \I__13160\ : Odrv4
    port map (
            O => \N__57190\,
            I => \c0.n30_adj_4233\
        );

    \I__13159\ : CascadeMux
    port map (
            O => \N__57187\,
            I => \N__57183\
        );

    \I__13158\ : InMux
    port map (
            O => \N__57186\,
            I => \N__57178\
        );

    \I__13157\ : InMux
    port map (
            O => \N__57183\,
            I => \N__57178\
        );

    \I__13156\ : LocalMux
    port map (
            O => \N__57178\,
            I => data_in_frame_14_2
        );

    \I__13155\ : InMux
    port map (
            O => \N__57175\,
            I => \N__57172\
        );

    \I__13154\ : LocalMux
    port map (
            O => \N__57172\,
            I => \N__57169\
        );

    \I__13153\ : Odrv4
    port map (
            O => \N__57169\,
            I => \c0.n22340\
        );

    \I__13152\ : InMux
    port map (
            O => \N__57166\,
            I => \N__57163\
        );

    \I__13151\ : LocalMux
    port map (
            O => \N__57163\,
            I => \N__57160\
        );

    \I__13150\ : Span4Mux_v
    port map (
            O => \N__57160\,
            I => \N__57151\
        );

    \I__13149\ : InMux
    port map (
            O => \N__57159\,
            I => \N__57146\
        );

    \I__13148\ : InMux
    port map (
            O => \N__57158\,
            I => \N__57146\
        );

    \I__13147\ : InMux
    port map (
            O => \N__57157\,
            I => \N__57143\
        );

    \I__13146\ : InMux
    port map (
            O => \N__57156\,
            I => \N__57136\
        );

    \I__13145\ : InMux
    port map (
            O => \N__57155\,
            I => \N__57136\
        );

    \I__13144\ : InMux
    port map (
            O => \N__57154\,
            I => \N__57136\
        );

    \I__13143\ : Odrv4
    port map (
            O => \N__57151\,
            I => n21755
        );

    \I__13142\ : LocalMux
    port map (
            O => \N__57146\,
            I => n21755
        );

    \I__13141\ : LocalMux
    port map (
            O => \N__57143\,
            I => n21755
        );

    \I__13140\ : LocalMux
    port map (
            O => \N__57136\,
            I => n21755
        );

    \I__13139\ : InMux
    port map (
            O => \N__57127\,
            I => \N__57123\
        );

    \I__13138\ : InMux
    port map (
            O => \N__57126\,
            I => \N__57120\
        );

    \I__13137\ : LocalMux
    port map (
            O => \N__57123\,
            I => data_in_frame_14_4
        );

    \I__13136\ : LocalMux
    port map (
            O => \N__57120\,
            I => data_in_frame_14_4
        );

    \I__13135\ : InMux
    port map (
            O => \N__57115\,
            I => \N__57112\
        );

    \I__13134\ : LocalMux
    port map (
            O => \N__57112\,
            I => n19619
        );

    \I__13133\ : InMux
    port map (
            O => \N__57109\,
            I => \N__57106\
        );

    \I__13132\ : LocalMux
    port map (
            O => \N__57106\,
            I => \N__57102\
        );

    \I__13131\ : InMux
    port map (
            O => \N__57105\,
            I => \N__57098\
        );

    \I__13130\ : Span4Mux_h
    port map (
            O => \N__57102\,
            I => \N__57095\
        );

    \I__13129\ : CascadeMux
    port map (
            O => \N__57101\,
            I => \N__57092\
        );

    \I__13128\ : LocalMux
    port map (
            O => \N__57098\,
            I => \N__57085\
        );

    \I__13127\ : Sp12to4
    port map (
            O => \N__57095\,
            I => \N__57085\
        );

    \I__13126\ : InMux
    port map (
            O => \N__57092\,
            I => \N__57082\
        );

    \I__13125\ : InMux
    port map (
            O => \N__57091\,
            I => \N__57079\
        );

    \I__13124\ : InMux
    port map (
            O => \N__57090\,
            I => \N__57076\
        );

    \I__13123\ : Span12Mux_v
    port map (
            O => \N__57085\,
            I => \N__57073\
        );

    \I__13122\ : LocalMux
    port map (
            O => \N__57082\,
            I => \r_Bit_Index_2\
        );

    \I__13121\ : LocalMux
    port map (
            O => \N__57079\,
            I => \r_Bit_Index_2\
        );

    \I__13120\ : LocalMux
    port map (
            O => \N__57076\,
            I => \r_Bit_Index_2\
        );

    \I__13119\ : Odrv12
    port map (
            O => \N__57073\,
            I => \r_Bit_Index_2\
        );

    \I__13118\ : CascadeMux
    port map (
            O => \N__57064\,
            I => \n91_cascade_\
        );

    \I__13117\ : InMux
    port map (
            O => \N__57061\,
            I => \N__57055\
        );

    \I__13116\ : InMux
    port map (
            O => \N__57060\,
            I => \N__57051\
        );

    \I__13115\ : InMux
    port map (
            O => \N__57059\,
            I => \N__57048\
        );

    \I__13114\ : InMux
    port map (
            O => \N__57058\,
            I => \N__57045\
        );

    \I__13113\ : LocalMux
    port map (
            O => \N__57055\,
            I => \N__57042\
        );

    \I__13112\ : InMux
    port map (
            O => \N__57054\,
            I => \N__57039\
        );

    \I__13111\ : LocalMux
    port map (
            O => \N__57051\,
            I => \r_SM_Main_2_N_3681_2\
        );

    \I__13110\ : LocalMux
    port map (
            O => \N__57048\,
            I => \r_SM_Main_2_N_3681_2\
        );

    \I__13109\ : LocalMux
    port map (
            O => \N__57045\,
            I => \r_SM_Main_2_N_3681_2\
        );

    \I__13108\ : Odrv4
    port map (
            O => \N__57042\,
            I => \r_SM_Main_2_N_3681_2\
        );

    \I__13107\ : LocalMux
    port map (
            O => \N__57039\,
            I => \r_SM_Main_2_N_3681_2\
        );

    \I__13106\ : InMux
    port map (
            O => \N__57028\,
            I => \N__57024\
        );

    \I__13105\ : InMux
    port map (
            O => \N__57027\,
            I => \N__57021\
        );

    \I__13104\ : LocalMux
    port map (
            O => \N__57024\,
            I => \N__57018\
        );

    \I__13103\ : LocalMux
    port map (
            O => \N__57021\,
            I => \N__57015\
        );

    \I__13102\ : Span4Mux_v
    port map (
            O => \N__57018\,
            I => \N__57012\
        );

    \I__13101\ : Span4Mux_h
    port map (
            O => \N__57015\,
            I => \N__57009\
        );

    \I__13100\ : Sp12to4
    port map (
            O => \N__57012\,
            I => \N__57004\
        );

    \I__13099\ : Span4Mux_v
    port map (
            O => \N__57009\,
            I => \N__56999\
        );

    \I__13098\ : InMux
    port map (
            O => \N__57008\,
            I => \N__56994\
        );

    \I__13097\ : InMux
    port map (
            O => \N__57007\,
            I => \N__56994\
        );

    \I__13096\ : Span12Mux_v
    port map (
            O => \N__57004\,
            I => \N__56988\
        );

    \I__13095\ : InMux
    port map (
            O => \N__57003\,
            I => \N__56985\
        );

    \I__13094\ : InMux
    port map (
            O => \N__57002\,
            I => \N__56982\
        );

    \I__13093\ : Span4Mux_h
    port map (
            O => \N__56999\,
            I => \N__56979\
        );

    \I__13092\ : LocalMux
    port map (
            O => \N__56994\,
            I => \N__56976\
        );

    \I__13091\ : InMux
    port map (
            O => \N__56993\,
            I => \N__56973\
        );

    \I__13090\ : InMux
    port map (
            O => \N__56992\,
            I => \N__56970\
        );

    \I__13089\ : InMux
    port map (
            O => \N__56991\,
            I => \N__56967\
        );

    \I__13088\ : Odrv12
    port map (
            O => \N__56988\,
            I => \r_SM_Main_2\
        );

    \I__13087\ : LocalMux
    port map (
            O => \N__56985\,
            I => \r_SM_Main_2\
        );

    \I__13086\ : LocalMux
    port map (
            O => \N__56982\,
            I => \r_SM_Main_2\
        );

    \I__13085\ : Odrv4
    port map (
            O => \N__56979\,
            I => \r_SM_Main_2\
        );

    \I__13084\ : Odrv4
    port map (
            O => \N__56976\,
            I => \r_SM_Main_2\
        );

    \I__13083\ : LocalMux
    port map (
            O => \N__56973\,
            I => \r_SM_Main_2\
        );

    \I__13082\ : LocalMux
    port map (
            O => \N__56970\,
            I => \r_SM_Main_2\
        );

    \I__13081\ : LocalMux
    port map (
            O => \N__56967\,
            I => \r_SM_Main_2\
        );

    \I__13080\ : InMux
    port map (
            O => \N__56950\,
            I => \N__56947\
        );

    \I__13079\ : LocalMux
    port map (
            O => \N__56947\,
            I => \N__56943\
        );

    \I__13078\ : CascadeMux
    port map (
            O => \N__56946\,
            I => \N__56940\
        );

    \I__13077\ : Span4Mux_v
    port map (
            O => \N__56943\,
            I => \N__56935\
        );

    \I__13076\ : InMux
    port map (
            O => \N__56940\,
            I => \N__56929\
        );

    \I__13075\ : InMux
    port map (
            O => \N__56939\,
            I => \N__56929\
        );

    \I__13074\ : CascadeMux
    port map (
            O => \N__56938\,
            I => \N__56924\
        );

    \I__13073\ : Span4Mux_v
    port map (
            O => \N__56935\,
            I => \N__56921\
        );

    \I__13072\ : InMux
    port map (
            O => \N__56934\,
            I => \N__56918\
        );

    \I__13071\ : LocalMux
    port map (
            O => \N__56929\,
            I => \N__56915\
        );

    \I__13070\ : CascadeMux
    port map (
            O => \N__56928\,
            I => \N__56911\
        );

    \I__13069\ : InMux
    port map (
            O => \N__56927\,
            I => \N__56905\
        );

    \I__13068\ : InMux
    port map (
            O => \N__56924\,
            I => \N__56905\
        );

    \I__13067\ : Span4Mux_v
    port map (
            O => \N__56921\,
            I => \N__56902\
        );

    \I__13066\ : LocalMux
    port map (
            O => \N__56918\,
            I => \N__56899\
        );

    \I__13065\ : Span4Mux_v
    port map (
            O => \N__56915\,
            I => \N__56895\
        );

    \I__13064\ : InMux
    port map (
            O => \N__56914\,
            I => \N__56890\
        );

    \I__13063\ : InMux
    port map (
            O => \N__56911\,
            I => \N__56890\
        );

    \I__13062\ : CascadeMux
    port map (
            O => \N__56910\,
            I => \N__56886\
        );

    \I__13061\ : LocalMux
    port map (
            O => \N__56905\,
            I => \N__56883\
        );

    \I__13060\ : Span4Mux_h
    port map (
            O => \N__56902\,
            I => \N__56878\
        );

    \I__13059\ : Span4Mux_v
    port map (
            O => \N__56899\,
            I => \N__56878\
        );

    \I__13058\ : InMux
    port map (
            O => \N__56898\,
            I => \N__56875\
        );

    \I__13057\ : Span4Mux_h
    port map (
            O => \N__56895\,
            I => \N__56870\
        );

    \I__13056\ : LocalMux
    port map (
            O => \N__56890\,
            I => \N__56870\
        );

    \I__13055\ : InMux
    port map (
            O => \N__56889\,
            I => \N__56867\
        );

    \I__13054\ : InMux
    port map (
            O => \N__56886\,
            I => \N__56864\
        );

    \I__13053\ : Span4Mux_h
    port map (
            O => \N__56883\,
            I => \N__56861\
        );

    \I__13052\ : Span4Mux_h
    port map (
            O => \N__56878\,
            I => \N__56858\
        );

    \I__13051\ : LocalMux
    port map (
            O => \N__56875\,
            I => \r_SM_Main_1\
        );

    \I__13050\ : Odrv4
    port map (
            O => \N__56870\,
            I => \r_SM_Main_1\
        );

    \I__13049\ : LocalMux
    port map (
            O => \N__56867\,
            I => \r_SM_Main_1\
        );

    \I__13048\ : LocalMux
    port map (
            O => \N__56864\,
            I => \r_SM_Main_1\
        );

    \I__13047\ : Odrv4
    port map (
            O => \N__56861\,
            I => \r_SM_Main_1\
        );

    \I__13046\ : Odrv4
    port map (
            O => \N__56858\,
            I => \r_SM_Main_1\
        );

    \I__13045\ : CascadeMux
    port map (
            O => \N__56845\,
            I => \c0.rx.n14_cascade_\
        );

    \I__13044\ : InMux
    port map (
            O => \N__56842\,
            I => \N__56839\
        );

    \I__13043\ : LocalMux
    port map (
            O => \N__56839\,
            I => \c0.rx.n36\
        );

    \I__13042\ : InMux
    port map (
            O => \N__56836\,
            I => \N__56832\
        );

    \I__13041\ : InMux
    port map (
            O => \N__56835\,
            I => \N__56829\
        );

    \I__13040\ : LocalMux
    port map (
            O => \N__56832\,
            I => \N__56823\
        );

    \I__13039\ : LocalMux
    port map (
            O => \N__56829\,
            I => \N__56819\
        );

    \I__13038\ : InMux
    port map (
            O => \N__56828\,
            I => \N__56811\
        );

    \I__13037\ : InMux
    port map (
            O => \N__56827\,
            I => \N__56811\
        );

    \I__13036\ : InMux
    port map (
            O => \N__56826\,
            I => \N__56811\
        );

    \I__13035\ : Span12Mux_h
    port map (
            O => \N__56823\,
            I => \N__56805\
        );

    \I__13034\ : InMux
    port map (
            O => \N__56822\,
            I => \N__56802\
        );

    \I__13033\ : Span4Mux_h
    port map (
            O => \N__56819\,
            I => \N__56799\
        );

    \I__13032\ : InMux
    port map (
            O => \N__56818\,
            I => \N__56796\
        );

    \I__13031\ : LocalMux
    port map (
            O => \N__56811\,
            I => \N__56793\
        );

    \I__13030\ : InMux
    port map (
            O => \N__56810\,
            I => \N__56788\
        );

    \I__13029\ : InMux
    port map (
            O => \N__56809\,
            I => \N__56788\
        );

    \I__13028\ : InMux
    port map (
            O => \N__56808\,
            I => \N__56785\
        );

    \I__13027\ : Odrv12
    port map (
            O => \N__56805\,
            I => \r_SM_Main_0\
        );

    \I__13026\ : LocalMux
    port map (
            O => \N__56802\,
            I => \r_SM_Main_0\
        );

    \I__13025\ : Odrv4
    port map (
            O => \N__56799\,
            I => \r_SM_Main_0\
        );

    \I__13024\ : LocalMux
    port map (
            O => \N__56796\,
            I => \r_SM_Main_0\
        );

    \I__13023\ : Odrv12
    port map (
            O => \N__56793\,
            I => \r_SM_Main_0\
        );

    \I__13022\ : LocalMux
    port map (
            O => \N__56788\,
            I => \r_SM_Main_0\
        );

    \I__13021\ : LocalMux
    port map (
            O => \N__56785\,
            I => \r_SM_Main_0\
        );

    \I__13020\ : CascadeMux
    port map (
            O => \N__56770\,
            I => \n21755_cascade_\
        );

    \I__13019\ : CascadeMux
    port map (
            O => \N__56767\,
            I => \N__56764\
        );

    \I__13018\ : InMux
    port map (
            O => \N__56764\,
            I => \N__56760\
        );

    \I__13017\ : InMux
    port map (
            O => \N__56763\,
            I => \N__56757\
        );

    \I__13016\ : LocalMux
    port map (
            O => \N__56760\,
            I => \N__56754\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__56757\,
            I => data_in_frame_14_1
        );

    \I__13014\ : Odrv4
    port map (
            O => \N__56754\,
            I => data_in_frame_14_1
        );

    \I__13013\ : CascadeMux
    port map (
            O => \N__56749\,
            I => \N__56745\
        );

    \I__13012\ : CascadeMux
    port map (
            O => \N__56748\,
            I => \N__56739\
        );

    \I__13011\ : InMux
    port map (
            O => \N__56745\,
            I => \N__56736\
        );

    \I__13010\ : CascadeMux
    port map (
            O => \N__56744\,
            I => \N__56733\
        );

    \I__13009\ : CascadeMux
    port map (
            O => \N__56743\,
            I => \N__56730\
        );

    \I__13008\ : CascadeMux
    port map (
            O => \N__56742\,
            I => \N__56726\
        );

    \I__13007\ : InMux
    port map (
            O => \N__56739\,
            I => \N__56723\
        );

    \I__13006\ : LocalMux
    port map (
            O => \N__56736\,
            I => \N__56720\
        );

    \I__13005\ : InMux
    port map (
            O => \N__56733\,
            I => \N__56715\
        );

    \I__13004\ : InMux
    port map (
            O => \N__56730\,
            I => \N__56712\
        );

    \I__13003\ : InMux
    port map (
            O => \N__56729\,
            I => \N__56709\
        );

    \I__13002\ : InMux
    port map (
            O => \N__56726\,
            I => \N__56705\
        );

    \I__13001\ : LocalMux
    port map (
            O => \N__56723\,
            I => \N__56700\
        );

    \I__13000\ : Span4Mux_v
    port map (
            O => \N__56720\,
            I => \N__56700\
        );

    \I__12999\ : CascadeMux
    port map (
            O => \N__56719\,
            I => \N__56696\
        );

    \I__12998\ : InMux
    port map (
            O => \N__56718\,
            I => \N__56693\
        );

    \I__12997\ : LocalMux
    port map (
            O => \N__56715\,
            I => \N__56688\
        );

    \I__12996\ : LocalMux
    port map (
            O => \N__56712\,
            I => \N__56683\
        );

    \I__12995\ : LocalMux
    port map (
            O => \N__56709\,
            I => \N__56683\
        );

    \I__12994\ : InMux
    port map (
            O => \N__56708\,
            I => \N__56680\
        );

    \I__12993\ : LocalMux
    port map (
            O => \N__56705\,
            I => \N__56675\
        );

    \I__12992\ : Span4Mux_v
    port map (
            O => \N__56700\,
            I => \N__56675\
        );

    \I__12991\ : InMux
    port map (
            O => \N__56699\,
            I => \N__56672\
        );

    \I__12990\ : InMux
    port map (
            O => \N__56696\,
            I => \N__56669\
        );

    \I__12989\ : LocalMux
    port map (
            O => \N__56693\,
            I => \N__56666\
        );

    \I__12988\ : InMux
    port map (
            O => \N__56692\,
            I => \N__56661\
        );

    \I__12987\ : InMux
    port map (
            O => \N__56691\,
            I => \N__56661\
        );

    \I__12986\ : Span4Mux_v
    port map (
            O => \N__56688\,
            I => \N__56658\
        );

    \I__12985\ : Span4Mux_v
    port map (
            O => \N__56683\,
            I => \N__56653\
        );

    \I__12984\ : LocalMux
    port map (
            O => \N__56680\,
            I => \N__56653\
        );

    \I__12983\ : Span4Mux_v
    port map (
            O => \N__56675\,
            I => \N__56648\
        );

    \I__12982\ : LocalMux
    port map (
            O => \N__56672\,
            I => \N__56648\
        );

    \I__12981\ : LocalMux
    port map (
            O => \N__56669\,
            I => \N__56645\
        );

    \I__12980\ : Span4Mux_v
    port map (
            O => \N__56666\,
            I => \N__56642\
        );

    \I__12979\ : LocalMux
    port map (
            O => \N__56661\,
            I => \N__56639\
        );

    \I__12978\ : Sp12to4
    port map (
            O => \N__56658\,
            I => \N__56636\
        );

    \I__12977\ : Span4Mux_h
    port map (
            O => \N__56653\,
            I => \N__56631\
        );

    \I__12976\ : Span4Mux_v
    port map (
            O => \N__56648\,
            I => \N__56631\
        );

    \I__12975\ : Span4Mux_v
    port map (
            O => \N__56645\,
            I => \N__56625\
        );

    \I__12974\ : Span4Mux_v
    port map (
            O => \N__56642\,
            I => \N__56625\
        );

    \I__12973\ : Span12Mux_h
    port map (
            O => \N__56639\,
            I => \N__56620\
        );

    \I__12972\ : Span12Mux_v
    port map (
            O => \N__56636\,
            I => \N__56620\
        );

    \I__12971\ : Span4Mux_v
    port map (
            O => \N__56631\,
            I => \N__56617\
        );

    \I__12970\ : InMux
    port map (
            O => \N__56630\,
            I => \N__56614\
        );

    \I__12969\ : Odrv4
    port map (
            O => \N__56625\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__12968\ : Odrv12
    port map (
            O => \N__56620\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__12967\ : Odrv4
    port map (
            O => \N__56617\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__12966\ : LocalMux
    port map (
            O => \N__56614\,
            I => \c0.FRAME_MATCHER_i_0\
        );

    \I__12965\ : InMux
    port map (
            O => \N__56605\,
            I => \N__56602\
        );

    \I__12964\ : LocalMux
    port map (
            O => \N__56602\,
            I => \N__56593\
        );

    \I__12963\ : InMux
    port map (
            O => \N__56601\,
            I => \N__56590\
        );

    \I__12962\ : InMux
    port map (
            O => \N__56600\,
            I => \N__56586\
        );

    \I__12961\ : InMux
    port map (
            O => \N__56599\,
            I => \N__56583\
        );

    \I__12960\ : InMux
    port map (
            O => \N__56598\,
            I => \N__56579\
        );

    \I__12959\ : InMux
    port map (
            O => \N__56597\,
            I => \N__56574\
        );

    \I__12958\ : InMux
    port map (
            O => \N__56596\,
            I => \N__56574\
        );

    \I__12957\ : Span4Mux_h
    port map (
            O => \N__56593\,
            I => \N__56570\
        );

    \I__12956\ : LocalMux
    port map (
            O => \N__56590\,
            I => \N__56565\
        );

    \I__12955\ : InMux
    port map (
            O => \N__56589\,
            I => \N__56562\
        );

    \I__12954\ : LocalMux
    port map (
            O => \N__56586\,
            I => \N__56557\
        );

    \I__12953\ : LocalMux
    port map (
            O => \N__56583\,
            I => \N__56557\
        );

    \I__12952\ : InMux
    port map (
            O => \N__56582\,
            I => \N__56554\
        );

    \I__12951\ : LocalMux
    port map (
            O => \N__56579\,
            I => \N__56551\
        );

    \I__12950\ : LocalMux
    port map (
            O => \N__56574\,
            I => \N__56548\
        );

    \I__12949\ : InMux
    port map (
            O => \N__56573\,
            I => \N__56545\
        );

    \I__12948\ : Span4Mux_v
    port map (
            O => \N__56570\,
            I => \N__56541\
        );

    \I__12947\ : InMux
    port map (
            O => \N__56569\,
            I => \N__56538\
        );

    \I__12946\ : InMux
    port map (
            O => \N__56568\,
            I => \N__56535\
        );

    \I__12945\ : Span4Mux_v
    port map (
            O => \N__56565\,
            I => \N__56530\
        );

    \I__12944\ : LocalMux
    port map (
            O => \N__56562\,
            I => \N__56530\
        );

    \I__12943\ : Span4Mux_h
    port map (
            O => \N__56557\,
            I => \N__56527\
        );

    \I__12942\ : LocalMux
    port map (
            O => \N__56554\,
            I => \N__56520\
        );

    \I__12941\ : Span4Mux_h
    port map (
            O => \N__56551\,
            I => \N__56520\
        );

    \I__12940\ : Span4Mux_v
    port map (
            O => \N__56548\,
            I => \N__56520\
        );

    \I__12939\ : LocalMux
    port map (
            O => \N__56545\,
            I => \N__56517\
        );

    \I__12938\ : CascadeMux
    port map (
            O => \N__56544\,
            I => \N__56514\
        );

    \I__12937\ : Span4Mux_v
    port map (
            O => \N__56541\,
            I => \N__56507\
        );

    \I__12936\ : LocalMux
    port map (
            O => \N__56538\,
            I => \N__56507\
        );

    \I__12935\ : LocalMux
    port map (
            O => \N__56535\,
            I => \N__56507\
        );

    \I__12934\ : Span4Mux_v
    port map (
            O => \N__56530\,
            I => \N__56504\
        );

    \I__12933\ : Sp12to4
    port map (
            O => \N__56527\,
            I => \N__56501\
        );

    \I__12932\ : Span4Mux_h
    port map (
            O => \N__56520\,
            I => \N__56496\
        );

    \I__12931\ : Span4Mux_h
    port map (
            O => \N__56517\,
            I => \N__56496\
        );

    \I__12930\ : InMux
    port map (
            O => \N__56514\,
            I => \N__56492\
        );

    \I__12929\ : Span4Mux_v
    port map (
            O => \N__56507\,
            I => \N__56487\
        );

    \I__12928\ : Span4Mux_v
    port map (
            O => \N__56504\,
            I => \N__56487\
        );

    \I__12927\ : Span12Mux_v
    port map (
            O => \N__56501\,
            I => \N__56484\
        );

    \I__12926\ : Span4Mux_v
    port map (
            O => \N__56496\,
            I => \N__56481\
        );

    \I__12925\ : InMux
    port map (
            O => \N__56495\,
            I => \N__56478\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__56492\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__12923\ : Odrv4
    port map (
            O => \N__56487\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__12922\ : Odrv12
    port map (
            O => \N__56484\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__12921\ : Odrv4
    port map (
            O => \N__56481\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__12920\ : LocalMux
    port map (
            O => \N__56478\,
            I => \c0.FRAME_MATCHER_i_1\
        );

    \I__12919\ : InMux
    port map (
            O => \N__56467\,
            I => \N__56462\
        );

    \I__12918\ : InMux
    port map (
            O => \N__56466\,
            I => \N__56459\
        );

    \I__12917\ : InMux
    port map (
            O => \N__56465\,
            I => \N__56452\
        );

    \I__12916\ : LocalMux
    port map (
            O => \N__56462\,
            I => \N__56449\
        );

    \I__12915\ : LocalMux
    port map (
            O => \N__56459\,
            I => \N__56446\
        );

    \I__12914\ : CascadeMux
    port map (
            O => \N__56458\,
            I => \N__56443\
        );

    \I__12913\ : InMux
    port map (
            O => \N__56457\,
            I => \N__56440\
        );

    \I__12912\ : InMux
    port map (
            O => \N__56456\,
            I => \N__56436\
        );

    \I__12911\ : InMux
    port map (
            O => \N__56455\,
            I => \N__56431\
        );

    \I__12910\ : LocalMux
    port map (
            O => \N__56452\,
            I => \N__56428\
        );

    \I__12909\ : Span4Mux_v
    port map (
            O => \N__56449\,
            I => \N__56423\
        );

    \I__12908\ : Span4Mux_v
    port map (
            O => \N__56446\,
            I => \N__56423\
        );

    \I__12907\ : InMux
    port map (
            O => \N__56443\,
            I => \N__56420\
        );

    \I__12906\ : LocalMux
    port map (
            O => \N__56440\,
            I => \N__56416\
        );

    \I__12905\ : InMux
    port map (
            O => \N__56439\,
            I => \N__56413\
        );

    \I__12904\ : LocalMux
    port map (
            O => \N__56436\,
            I => \N__56410\
        );

    \I__12903\ : InMux
    port map (
            O => \N__56435\,
            I => \N__56407\
        );

    \I__12902\ : InMux
    port map (
            O => \N__56434\,
            I => \N__56404\
        );

    \I__12901\ : LocalMux
    port map (
            O => \N__56431\,
            I => \N__56400\
        );

    \I__12900\ : Span4Mux_v
    port map (
            O => \N__56428\,
            I => \N__56395\
        );

    \I__12899\ : Span4Mux_v
    port map (
            O => \N__56423\,
            I => \N__56395\
        );

    \I__12898\ : LocalMux
    port map (
            O => \N__56420\,
            I => \N__56391\
        );

    \I__12897\ : InMux
    port map (
            O => \N__56419\,
            I => \N__56388\
        );

    \I__12896\ : Span4Mux_v
    port map (
            O => \N__56416\,
            I => \N__56383\
        );

    \I__12895\ : LocalMux
    port map (
            O => \N__56413\,
            I => \N__56383\
        );

    \I__12894\ : Span4Mux_v
    port map (
            O => \N__56410\,
            I => \N__56376\
        );

    \I__12893\ : LocalMux
    port map (
            O => \N__56407\,
            I => \N__56376\
        );

    \I__12892\ : LocalMux
    port map (
            O => \N__56404\,
            I => \N__56376\
        );

    \I__12891\ : CascadeMux
    port map (
            O => \N__56403\,
            I => \N__56373\
        );

    \I__12890\ : Span4Mux_v
    port map (
            O => \N__56400\,
            I => \N__56370\
        );

    \I__12889\ : Span4Mux_v
    port map (
            O => \N__56395\,
            I => \N__56367\
        );

    \I__12888\ : InMux
    port map (
            O => \N__56394\,
            I => \N__56364\
        );

    \I__12887\ : Span4Mux_h
    port map (
            O => \N__56391\,
            I => \N__56357\
        );

    \I__12886\ : LocalMux
    port map (
            O => \N__56388\,
            I => \N__56357\
        );

    \I__12885\ : Span4Mux_h
    port map (
            O => \N__56383\,
            I => \N__56357\
        );

    \I__12884\ : Span4Mux_v
    port map (
            O => \N__56376\,
            I => \N__56354\
        );

    \I__12883\ : InMux
    port map (
            O => \N__56373\,
            I => \N__56350\
        );

    \I__12882\ : Span4Mux_v
    port map (
            O => \N__56370\,
            I => \N__56345\
        );

    \I__12881\ : Span4Mux_v
    port map (
            O => \N__56367\,
            I => \N__56345\
        );

    \I__12880\ : LocalMux
    port map (
            O => \N__56364\,
            I => \N__56338\
        );

    \I__12879\ : Span4Mux_v
    port map (
            O => \N__56357\,
            I => \N__56338\
        );

    \I__12878\ : Span4Mux_h
    port map (
            O => \N__56354\,
            I => \N__56338\
        );

    \I__12877\ : InMux
    port map (
            O => \N__56353\,
            I => \N__56335\
        );

    \I__12876\ : LocalMux
    port map (
            O => \N__56350\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__12875\ : Odrv4
    port map (
            O => \N__56345\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__12874\ : Odrv4
    port map (
            O => \N__56338\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__12873\ : LocalMux
    port map (
            O => \N__56335\,
            I => \c0.FRAME_MATCHER_i_2\
        );

    \I__12872\ : InMux
    port map (
            O => \N__56326\,
            I => \N__56323\
        );

    \I__12871\ : LocalMux
    port map (
            O => \N__56323\,
            I => \N__56319\
        );

    \I__12870\ : InMux
    port map (
            O => \N__56322\,
            I => \N__56316\
        );

    \I__12869\ : Span4Mux_h
    port map (
            O => \N__56319\,
            I => \N__56311\
        );

    \I__12868\ : LocalMux
    port map (
            O => \N__56316\,
            I => \N__56311\
        );

    \I__12867\ : Odrv4
    port map (
            O => \N__56311\,
            I => \c0.n20370\
        );

    \I__12866\ : CascadeMux
    port map (
            O => \N__56308\,
            I => \N__56305\
        );

    \I__12865\ : InMux
    port map (
            O => \N__56305\,
            I => \N__56301\
        );

    \I__12864\ : InMux
    port map (
            O => \N__56304\,
            I => \N__56298\
        );

    \I__12863\ : LocalMux
    port map (
            O => \N__56301\,
            I => \c0.data_in_frame_29_5\
        );

    \I__12862\ : LocalMux
    port map (
            O => \N__56298\,
            I => \c0.data_in_frame_29_5\
        );

    \I__12861\ : InMux
    port map (
            O => \N__56293\,
            I => \N__56290\
        );

    \I__12860\ : LocalMux
    port map (
            O => \N__56290\,
            I => \N__56287\
        );

    \I__12859\ : Odrv4
    port map (
            O => \N__56287\,
            I => \c0.n22157\
        );

    \I__12858\ : CascadeMux
    port map (
            O => \N__56284\,
            I => \N__56280\
        );

    \I__12857\ : CascadeMux
    port map (
            O => \N__56283\,
            I => \N__56275\
        );

    \I__12856\ : InMux
    port map (
            O => \N__56280\,
            I => \N__56272\
        );

    \I__12855\ : InMux
    port map (
            O => \N__56279\,
            I => \N__56269\
        );

    \I__12854\ : InMux
    port map (
            O => \N__56278\,
            I => \N__56266\
        );

    \I__12853\ : InMux
    port map (
            O => \N__56275\,
            I => \N__56263\
        );

    \I__12852\ : LocalMux
    port map (
            O => \N__56272\,
            I => \N__56258\
        );

    \I__12851\ : LocalMux
    port map (
            O => \N__56269\,
            I => \N__56258\
        );

    \I__12850\ : LocalMux
    port map (
            O => \N__56266\,
            I => \N__56253\
        );

    \I__12849\ : LocalMux
    port map (
            O => \N__56263\,
            I => \N__56253\
        );

    \I__12848\ : Odrv4
    port map (
            O => \N__56258\,
            I => \c0.data_in_frame_27_3\
        );

    \I__12847\ : Odrv12
    port map (
            O => \N__56253\,
            I => \c0.data_in_frame_27_3\
        );

    \I__12846\ : InMux
    port map (
            O => \N__56248\,
            I => \N__56245\
        );

    \I__12845\ : LocalMux
    port map (
            O => \N__56245\,
            I => \c0.n22719\
        );

    \I__12844\ : CascadeMux
    port map (
            O => \N__56242\,
            I => \c0.n8_adj_4291_cascade_\
        );

    \I__12843\ : InMux
    port map (
            O => \N__56239\,
            I => \N__56236\
        );

    \I__12842\ : LocalMux
    port map (
            O => \N__56236\,
            I => \c0.n22148\
        );

    \I__12841\ : InMux
    port map (
            O => \N__56233\,
            I => \N__56230\
        );

    \I__12840\ : LocalMux
    port map (
            O => \N__56230\,
            I => \N__56227\
        );

    \I__12839\ : Span4Mux_h
    port map (
            O => \N__56227\,
            I => \N__56224\
        );

    \I__12838\ : Odrv4
    port map (
            O => \N__56224\,
            I => \c0.n23811\
        );

    \I__12837\ : InMux
    port map (
            O => \N__56221\,
            I => \N__56217\
        );

    \I__12836\ : CascadeMux
    port map (
            O => \N__56220\,
            I => \N__56214\
        );

    \I__12835\ : LocalMux
    port map (
            O => \N__56217\,
            I => \N__56211\
        );

    \I__12834\ : InMux
    port map (
            O => \N__56214\,
            I => \N__56208\
        );

    \I__12833\ : Span4Mux_h
    port map (
            O => \N__56211\,
            I => \N__56204\
        );

    \I__12832\ : LocalMux
    port map (
            O => \N__56208\,
            I => \N__56201\
        );

    \I__12831\ : InMux
    port map (
            O => \N__56207\,
            I => \N__56198\
        );

    \I__12830\ : Span4Mux_v
    port map (
            O => \N__56204\,
            I => \N__56195\
        );

    \I__12829\ : Odrv4
    port map (
            O => \N__56201\,
            I => n12977
        );

    \I__12828\ : LocalMux
    port map (
            O => \N__56198\,
            I => n12977
        );

    \I__12827\ : Odrv4
    port map (
            O => \N__56195\,
            I => n12977
        );

    \I__12826\ : InMux
    port map (
            O => \N__56188\,
            I => \N__56181\
        );

    \I__12825\ : InMux
    port map (
            O => \N__56187\,
            I => \N__56181\
        );

    \I__12824\ : InMux
    port map (
            O => \N__56186\,
            I => \N__56178\
        );

    \I__12823\ : LocalMux
    port map (
            O => \N__56181\,
            I => \N__56175\
        );

    \I__12822\ : LocalMux
    port map (
            O => \N__56178\,
            I => \N__56172\
        );

    \I__12821\ : Span4Mux_v
    port map (
            O => \N__56175\,
            I => \N__56169\
        );

    \I__12820\ : Odrv4
    port map (
            O => \N__56172\,
            I => \c0.rx.n21704\
        );

    \I__12819\ : Odrv4
    port map (
            O => \N__56169\,
            I => \c0.rx.n21704\
        );

    \I__12818\ : CascadeMux
    port map (
            O => \N__56164\,
            I => \n14436_cascade_\
        );

    \I__12817\ : InMux
    port map (
            O => \N__56161\,
            I => \N__56157\
        );

    \I__12816\ : InMux
    port map (
            O => \N__56160\,
            I => \N__56154\
        );

    \I__12815\ : LocalMux
    port map (
            O => \N__56157\,
            I => \c0.rx.n12862\
        );

    \I__12814\ : LocalMux
    port map (
            O => \N__56154\,
            I => \c0.rx.n12862\
        );

    \I__12813\ : CascadeMux
    port map (
            O => \N__56149\,
            I => \N__56146\
        );

    \I__12812\ : InMux
    port map (
            O => \N__56146\,
            I => \N__56143\
        );

    \I__12811\ : LocalMux
    port map (
            O => \N__56143\,
            I => \N__56139\
        );

    \I__12810\ : InMux
    port map (
            O => \N__56142\,
            I => \N__56135\
        );

    \I__12809\ : Span4Mux_v
    port map (
            O => \N__56139\,
            I => \N__56132\
        );

    \I__12808\ : CascadeMux
    port map (
            O => \N__56138\,
            I => \N__56129\
        );

    \I__12807\ : LocalMux
    port map (
            O => \N__56135\,
            I => \N__56126\
        );

    \I__12806\ : Span4Mux_v
    port map (
            O => \N__56132\,
            I => \N__56123\
        );

    \I__12805\ : InMux
    port map (
            O => \N__56129\,
            I => \N__56120\
        );

    \I__12804\ : Span12Mux_v
    port map (
            O => \N__56126\,
            I => \N__56117\
        );

    \I__12803\ : Span4Mux_h
    port map (
            O => \N__56123\,
            I => \N__56114\
        );

    \I__12802\ : LocalMux
    port map (
            O => \N__56120\,
            I => \c0.data_in_frame_25_1\
        );

    \I__12801\ : Odrv12
    port map (
            O => \N__56117\,
            I => \c0.data_in_frame_25_1\
        );

    \I__12800\ : Odrv4
    port map (
            O => \N__56114\,
            I => \c0.data_in_frame_25_1\
        );

    \I__12799\ : InMux
    port map (
            O => \N__56107\,
            I => \N__56104\
        );

    \I__12798\ : LocalMux
    port map (
            O => \N__56104\,
            I => \N__56101\
        );

    \I__12797\ : Span4Mux_v
    port map (
            O => \N__56101\,
            I => \N__56098\
        );

    \I__12796\ : Span4Mux_h
    port map (
            O => \N__56098\,
            I => \N__56095\
        );

    \I__12795\ : Odrv4
    port map (
            O => \N__56095\,
            I => \c0.n49_adj_4488\
        );

    \I__12794\ : InMux
    port map (
            O => \N__56092\,
            I => \N__56089\
        );

    \I__12793\ : LocalMux
    port map (
            O => \N__56089\,
            I => \c0.n55\
        );

    \I__12792\ : InMux
    port map (
            O => \N__56086\,
            I => \N__56083\
        );

    \I__12791\ : LocalMux
    port map (
            O => \N__56083\,
            I => \c0.n53\
        );

    \I__12790\ : InMux
    port map (
            O => \N__56080\,
            I => \N__56077\
        );

    \I__12789\ : LocalMux
    port map (
            O => \N__56077\,
            I => \N__56074\
        );

    \I__12788\ : Span4Mux_h
    port map (
            O => \N__56074\,
            I => \N__56071\
        );

    \I__12787\ : Odrv4
    port map (
            O => \N__56071\,
            I => \c0.n23416\
        );

    \I__12786\ : CascadeMux
    port map (
            O => \N__56068\,
            I => \c0.n23416_cascade_\
        );

    \I__12785\ : InMux
    port map (
            O => \N__56065\,
            I => \N__56062\
        );

    \I__12784\ : LocalMux
    port map (
            O => \N__56062\,
            I => \c0.n12_adj_4296\
        );

    \I__12783\ : InMux
    port map (
            O => \N__56059\,
            I => \N__56054\
        );

    \I__12782\ : CascadeMux
    port map (
            O => \N__56058\,
            I => \N__56050\
        );

    \I__12781\ : InMux
    port map (
            O => \N__56057\,
            I => \N__56047\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__56054\,
            I => \N__56044\
        );

    \I__12779\ : InMux
    port map (
            O => \N__56053\,
            I => \N__56041\
        );

    \I__12778\ : InMux
    port map (
            O => \N__56050\,
            I => \N__56038\
        );

    \I__12777\ : LocalMux
    port map (
            O => \N__56047\,
            I => \N__56035\
        );

    \I__12776\ : Span4Mux_h
    port map (
            O => \N__56044\,
            I => \N__56032\
        );

    \I__12775\ : LocalMux
    port map (
            O => \N__56041\,
            I => \N__56029\
        );

    \I__12774\ : LocalMux
    port map (
            O => \N__56038\,
            I => \c0.data_in_frame_27_2\
        );

    \I__12773\ : Odrv4
    port map (
            O => \N__56035\,
            I => \c0.data_in_frame_27_2\
        );

    \I__12772\ : Odrv4
    port map (
            O => \N__56032\,
            I => \c0.data_in_frame_27_2\
        );

    \I__12771\ : Odrv12
    port map (
            O => \N__56029\,
            I => \c0.data_in_frame_27_2\
        );

    \I__12770\ : InMux
    port map (
            O => \N__56020\,
            I => \N__56017\
        );

    \I__12769\ : LocalMux
    port map (
            O => \N__56017\,
            I => \c0.n36_adj_4489\
        );

    \I__12768\ : CascadeMux
    port map (
            O => \N__56014\,
            I => \N__56011\
        );

    \I__12767\ : InMux
    port map (
            O => \N__56011\,
            I => \N__56007\
        );

    \I__12766\ : InMux
    port map (
            O => \N__56010\,
            I => \N__56003\
        );

    \I__12765\ : LocalMux
    port map (
            O => \N__56007\,
            I => \N__56000\
        );

    \I__12764\ : CascadeMux
    port map (
            O => \N__56006\,
            I => \N__55996\
        );

    \I__12763\ : LocalMux
    port map (
            O => \N__56003\,
            I => \N__55993\
        );

    \I__12762\ : Span4Mux_h
    port map (
            O => \N__56000\,
            I => \N__55990\
        );

    \I__12761\ : InMux
    port map (
            O => \N__55999\,
            I => \N__55987\
        );

    \I__12760\ : InMux
    port map (
            O => \N__55996\,
            I => \N__55984\
        );

    \I__12759\ : Span4Mux_h
    port map (
            O => \N__55993\,
            I => \N__55981\
        );

    \I__12758\ : Span4Mux_v
    port map (
            O => \N__55990\,
            I => \N__55978\
        );

    \I__12757\ : LocalMux
    port map (
            O => \N__55987\,
            I => \N__55975\
        );

    \I__12756\ : LocalMux
    port map (
            O => \N__55984\,
            I => \c0.data_in_frame_19_2\
        );

    \I__12755\ : Odrv4
    port map (
            O => \N__55981\,
            I => \c0.data_in_frame_19_2\
        );

    \I__12754\ : Odrv4
    port map (
            O => \N__55978\,
            I => \c0.data_in_frame_19_2\
        );

    \I__12753\ : Odrv4
    port map (
            O => \N__55975\,
            I => \c0.data_in_frame_19_2\
        );

    \I__12752\ : InMux
    port map (
            O => \N__55966\,
            I => \N__55959\
        );

    \I__12751\ : InMux
    port map (
            O => \N__55965\,
            I => \N__55959\
        );

    \I__12750\ : InMux
    port map (
            O => \N__55964\,
            I => \N__55956\
        );

    \I__12749\ : LocalMux
    port map (
            O => \N__55959\,
            I => \N__55953\
        );

    \I__12748\ : LocalMux
    port map (
            O => \N__55956\,
            I => \N__55948\
        );

    \I__12747\ : Span4Mux_v
    port map (
            O => \N__55953\,
            I => \N__55948\
        );

    \I__12746\ : Odrv4
    port map (
            O => \N__55948\,
            I => \c0.n6221\
        );

    \I__12745\ : CascadeMux
    port map (
            O => \N__55945\,
            I => \N__55942\
        );

    \I__12744\ : InMux
    port map (
            O => \N__55942\,
            I => \N__55939\
        );

    \I__12743\ : LocalMux
    port map (
            O => \N__55939\,
            I => \N__55935\
        );

    \I__12742\ : InMux
    port map (
            O => \N__55938\,
            I => \N__55932\
        );

    \I__12741\ : Span4Mux_h
    port map (
            O => \N__55935\,
            I => \N__55929\
        );

    \I__12740\ : LocalMux
    port map (
            O => \N__55932\,
            I => \c0.n21037\
        );

    \I__12739\ : Odrv4
    port map (
            O => \N__55929\,
            I => \c0.n21037\
        );

    \I__12738\ : InMux
    port map (
            O => \N__55924\,
            I => \N__55921\
        );

    \I__12737\ : LocalMux
    port map (
            O => \N__55921\,
            I => \N__55916\
        );

    \I__12736\ : InMux
    port map (
            O => \N__55920\,
            I => \N__55911\
        );

    \I__12735\ : InMux
    port map (
            O => \N__55919\,
            I => \N__55911\
        );

    \I__12734\ : Span4Mux_h
    port map (
            O => \N__55916\,
            I => \N__55908\
        );

    \I__12733\ : LocalMux
    port map (
            O => \N__55911\,
            I => \N__55905\
        );

    \I__12732\ : Odrv4
    port map (
            O => \N__55908\,
            I => \c0.data_in_frame_23_6\
        );

    \I__12731\ : Odrv4
    port map (
            O => \N__55905\,
            I => \c0.data_in_frame_23_6\
        );

    \I__12730\ : CascadeMux
    port map (
            O => \N__55900\,
            I => \c0.n21037_cascade_\
        );

    \I__12729\ : CascadeMux
    port map (
            O => \N__55897\,
            I => \N__55891\
        );

    \I__12728\ : InMux
    port map (
            O => \N__55896\,
            I => \N__55887\
        );

    \I__12727\ : InMux
    port map (
            O => \N__55895\,
            I => \N__55884\
        );

    \I__12726\ : InMux
    port map (
            O => \N__55894\,
            I => \N__55877\
        );

    \I__12725\ : InMux
    port map (
            O => \N__55891\,
            I => \N__55877\
        );

    \I__12724\ : InMux
    port map (
            O => \N__55890\,
            I => \N__55877\
        );

    \I__12723\ : LocalMux
    port map (
            O => \N__55887\,
            I => \N__55873\
        );

    \I__12722\ : LocalMux
    port map (
            O => \N__55884\,
            I => \N__55870\
        );

    \I__12721\ : LocalMux
    port map (
            O => \N__55877\,
            I => \N__55867\
        );

    \I__12720\ : InMux
    port map (
            O => \N__55876\,
            I => \N__55864\
        );

    \I__12719\ : Span4Mux_v
    port map (
            O => \N__55873\,
            I => \N__55861\
        );

    \I__12718\ : Span4Mux_h
    port map (
            O => \N__55870\,
            I => \N__55858\
        );

    \I__12717\ : Span4Mux_h
    port map (
            O => \N__55867\,
            I => \N__55855\
        );

    \I__12716\ : LocalMux
    port map (
            O => \N__55864\,
            I => \c0.data_in_frame_19_4\
        );

    \I__12715\ : Odrv4
    port map (
            O => \N__55861\,
            I => \c0.data_in_frame_19_4\
        );

    \I__12714\ : Odrv4
    port map (
            O => \N__55858\,
            I => \c0.data_in_frame_19_4\
        );

    \I__12713\ : Odrv4
    port map (
            O => \N__55855\,
            I => \c0.data_in_frame_19_4\
        );

    \I__12712\ : InMux
    port map (
            O => \N__55846\,
            I => \N__55843\
        );

    \I__12711\ : LocalMux
    port map (
            O => \N__55843\,
            I => \c0.n13282\
        );

    \I__12710\ : CascadeMux
    port map (
            O => \N__55840\,
            I => \N__55836\
        );

    \I__12709\ : CascadeMux
    port map (
            O => \N__55839\,
            I => \N__55833\
        );

    \I__12708\ : InMux
    port map (
            O => \N__55836\,
            I => \N__55830\
        );

    \I__12707\ : InMux
    port map (
            O => \N__55833\,
            I => \N__55826\
        );

    \I__12706\ : LocalMux
    port map (
            O => \N__55830\,
            I => \N__55823\
        );

    \I__12705\ : InMux
    port map (
            O => \N__55829\,
            I => \N__55820\
        );

    \I__12704\ : LocalMux
    port map (
            O => \N__55826\,
            I => \N__55815\
        );

    \I__12703\ : Span4Mux_h
    port map (
            O => \N__55823\,
            I => \N__55815\
        );

    \I__12702\ : LocalMux
    port map (
            O => \N__55820\,
            I => \c0.data_in_frame_27_4\
        );

    \I__12701\ : Odrv4
    port map (
            O => \N__55815\,
            I => \c0.data_in_frame_27_4\
        );

    \I__12700\ : CascadeMux
    port map (
            O => \N__55810\,
            I => \c0.n52_cascade_\
        );

    \I__12699\ : InMux
    port map (
            O => \N__55807\,
            I => \N__55804\
        );

    \I__12698\ : LocalMux
    port map (
            O => \N__55804\,
            I => \N__55801\
        );

    \I__12697\ : Odrv4
    port map (
            O => \N__55801\,
            I => \c0.n13872\
        );

    \I__12696\ : InMux
    port map (
            O => \N__55798\,
            I => \N__55795\
        );

    \I__12695\ : LocalMux
    port map (
            O => \N__55795\,
            I => \N__55791\
        );

    \I__12694\ : InMux
    port map (
            O => \N__55794\,
            I => \N__55788\
        );

    \I__12693\ : Odrv12
    port map (
            O => \N__55791\,
            I => \c0.n12420\
        );

    \I__12692\ : LocalMux
    port map (
            O => \N__55788\,
            I => \c0.n12420\
        );

    \I__12691\ : InMux
    port map (
            O => \N__55783\,
            I => \N__55780\
        );

    \I__12690\ : LocalMux
    port map (
            O => \N__55780\,
            I => \N__55777\
        );

    \I__12689\ : Odrv4
    port map (
            O => \N__55777\,
            I => \c0.n23615\
        );

    \I__12688\ : InMux
    port map (
            O => \N__55774\,
            I => \N__55771\
        );

    \I__12687\ : LocalMux
    port map (
            O => \N__55771\,
            I => \c0.n44_adj_4490\
        );

    \I__12686\ : CascadeMux
    port map (
            O => \N__55768\,
            I => \c0.n48_adj_4485_cascade_\
        );

    \I__12685\ : InMux
    port map (
            O => \N__55765\,
            I => \N__55762\
        );

    \I__12684\ : LocalMux
    port map (
            O => \N__55762\,
            I => \N__55759\
        );

    \I__12683\ : Span4Mux_h
    port map (
            O => \N__55759\,
            I => \N__55756\
        );

    \I__12682\ : Odrv4
    port map (
            O => \N__55756\,
            I => \c0.n12_adj_4290\
        );

    \I__12681\ : InMux
    port map (
            O => \N__55753\,
            I => \N__55750\
        );

    \I__12680\ : LocalMux
    port map (
            O => \N__55750\,
            I => \N__55746\
        );

    \I__12679\ : InMux
    port map (
            O => \N__55749\,
            I => \N__55743\
        );

    \I__12678\ : Span4Mux_v
    port map (
            O => \N__55746\,
            I => \N__55738\
        );

    \I__12677\ : LocalMux
    port map (
            O => \N__55743\,
            I => \N__55738\
        );

    \I__12676\ : Span4Mux_v
    port map (
            O => \N__55738\,
            I => \N__55735\
        );

    \I__12675\ : Odrv4
    port map (
            O => \N__55735\,
            I => \c0.n22355\
        );

    \I__12674\ : CascadeMux
    port map (
            O => \N__55732\,
            I => \c0.n23062_cascade_\
        );

    \I__12673\ : CascadeMux
    port map (
            O => \N__55729\,
            I => \N__55725\
        );

    \I__12672\ : CascadeMux
    port map (
            O => \N__55728\,
            I => \N__55721\
        );

    \I__12671\ : InMux
    port map (
            O => \N__55725\,
            I => \N__55718\
        );

    \I__12670\ : InMux
    port map (
            O => \N__55724\,
            I => \N__55715\
        );

    \I__12669\ : InMux
    port map (
            O => \N__55721\,
            I => \N__55712\
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__55718\,
            I => \N__55709\
        );

    \I__12667\ : LocalMux
    port map (
            O => \N__55715\,
            I => \N__55706\
        );

    \I__12666\ : LocalMux
    port map (
            O => \N__55712\,
            I => \N__55703\
        );

    \I__12665\ : Span4Mux_v
    port map (
            O => \N__55709\,
            I => \N__55700\
        );

    \I__12664\ : Span4Mux_v
    port map (
            O => \N__55706\,
            I => \N__55697\
        );

    \I__12663\ : Odrv4
    port map (
            O => \N__55703\,
            I => \c0.data_in_frame_21_0\
        );

    \I__12662\ : Odrv4
    port map (
            O => \N__55700\,
            I => \c0.data_in_frame_21_0\
        );

    \I__12661\ : Odrv4
    port map (
            O => \N__55697\,
            I => \c0.data_in_frame_21_0\
        );

    \I__12660\ : InMux
    port map (
            O => \N__55690\,
            I => \N__55687\
        );

    \I__12659\ : LocalMux
    port map (
            O => \N__55687\,
            I => \c0.n23062\
        );

    \I__12658\ : InMux
    port map (
            O => \N__55684\,
            I => \N__55681\
        );

    \I__12657\ : LocalMux
    port map (
            O => \N__55681\,
            I => \c0.n8\
        );

    \I__12656\ : InMux
    port map (
            O => \N__55678\,
            I => \N__55675\
        );

    \I__12655\ : LocalMux
    port map (
            O => \N__55675\,
            I => \c0.n27\
        );

    \I__12654\ : InMux
    port map (
            O => \N__55672\,
            I => \N__55669\
        );

    \I__12653\ : LocalMux
    port map (
            O => \N__55669\,
            I => \N__55665\
        );

    \I__12652\ : InMux
    port map (
            O => \N__55668\,
            I => \N__55662\
        );

    \I__12651\ : Span4Mux_v
    port map (
            O => \N__55665\,
            I => \N__55659\
        );

    \I__12650\ : LocalMux
    port map (
            O => \N__55662\,
            I => \N__55656\
        );

    \I__12649\ : Span4Mux_v
    port map (
            O => \N__55659\,
            I => \N__55653\
        );

    \I__12648\ : Span4Mux_v
    port map (
            O => \N__55656\,
            I => \N__55650\
        );

    \I__12647\ : Odrv4
    port map (
            O => \N__55653\,
            I => \c0.n22296\
        );

    \I__12646\ : Odrv4
    port map (
            O => \N__55650\,
            I => \c0.n22296\
        );

    \I__12645\ : InMux
    port map (
            O => \N__55645\,
            I => \N__55642\
        );

    \I__12644\ : LocalMux
    port map (
            O => \N__55642\,
            I => \N__55638\
        );

    \I__12643\ : InMux
    port map (
            O => \N__55641\,
            I => \N__55635\
        );

    \I__12642\ : Span4Mux_v
    port map (
            O => \N__55638\,
            I => \N__55630\
        );

    \I__12641\ : LocalMux
    port map (
            O => \N__55635\,
            I => \N__55630\
        );

    \I__12640\ : Odrv4
    port map (
            O => \N__55630\,
            I => \c0.n21831\
        );

    \I__12639\ : CascadeMux
    port map (
            O => \N__55627\,
            I => \N__55620\
        );

    \I__12638\ : InMux
    port map (
            O => \N__55626\,
            I => \N__55617\
        );

    \I__12637\ : InMux
    port map (
            O => \N__55625\,
            I => \N__55614\
        );

    \I__12636\ : InMux
    port map (
            O => \N__55624\,
            I => \N__55609\
        );

    \I__12635\ : InMux
    port map (
            O => \N__55623\,
            I => \N__55609\
        );

    \I__12634\ : InMux
    port map (
            O => \N__55620\,
            I => \N__55606\
        );

    \I__12633\ : LocalMux
    port map (
            O => \N__55617\,
            I => \N__55603\
        );

    \I__12632\ : LocalMux
    port map (
            O => \N__55614\,
            I => \N__55600\
        );

    \I__12631\ : LocalMux
    port map (
            O => \N__55609\,
            I => \N__55597\
        );

    \I__12630\ : LocalMux
    port map (
            O => \N__55606\,
            I => \N__55594\
        );

    \I__12629\ : Span4Mux_h
    port map (
            O => \N__55603\,
            I => \N__55591\
        );

    \I__12628\ : Span4Mux_h
    port map (
            O => \N__55600\,
            I => \N__55588\
        );

    \I__12627\ : Span4Mux_h
    port map (
            O => \N__55597\,
            I => \N__55585\
        );

    \I__12626\ : Odrv4
    port map (
            O => \N__55594\,
            I => \c0.data_in_frame_17_0\
        );

    \I__12625\ : Odrv4
    port map (
            O => \N__55591\,
            I => \c0.data_in_frame_17_0\
        );

    \I__12624\ : Odrv4
    port map (
            O => \N__55588\,
            I => \c0.data_in_frame_17_0\
        );

    \I__12623\ : Odrv4
    port map (
            O => \N__55585\,
            I => \c0.data_in_frame_17_0\
        );

    \I__12622\ : CascadeMux
    port map (
            O => \N__55576\,
            I => \c0.n16_adj_4223_cascade_\
        );

    \I__12621\ : InMux
    port map (
            O => \N__55573\,
            I => \N__55570\
        );

    \I__12620\ : LocalMux
    port map (
            O => \N__55570\,
            I => \N__55567\
        );

    \I__12619\ : Odrv12
    port map (
            O => \N__55567\,
            I => \c0.n17\
        );

    \I__12618\ : InMux
    port map (
            O => \N__55564\,
            I => \N__55558\
        );

    \I__12617\ : InMux
    port map (
            O => \N__55563\,
            I => \N__55558\
        );

    \I__12616\ : LocalMux
    port map (
            O => \N__55558\,
            I => \N__55554\
        );

    \I__12615\ : InMux
    port map (
            O => \N__55557\,
            I => \N__55551\
        );

    \I__12614\ : Span4Mux_h
    port map (
            O => \N__55554\,
            I => \N__55548\
        );

    \I__12613\ : LocalMux
    port map (
            O => \N__55551\,
            I => \c0.n21187\
        );

    \I__12612\ : Odrv4
    port map (
            O => \N__55548\,
            I => \c0.n21187\
        );

    \I__12611\ : CascadeMux
    port map (
            O => \N__55543\,
            I => \c0.n22211_cascade_\
        );

    \I__12610\ : InMux
    port map (
            O => \N__55540\,
            I => \N__55536\
        );

    \I__12609\ : InMux
    port map (
            O => \N__55539\,
            I => \N__55531\
        );

    \I__12608\ : LocalMux
    port map (
            O => \N__55536\,
            I => \N__55528\
        );

    \I__12607\ : InMux
    port map (
            O => \N__55535\,
            I => \N__55525\
        );

    \I__12606\ : InMux
    port map (
            O => \N__55534\,
            I => \N__55522\
        );

    \I__12605\ : LocalMux
    port map (
            O => \N__55531\,
            I => \c0.n21140\
        );

    \I__12604\ : Odrv4
    port map (
            O => \N__55528\,
            I => \c0.n21140\
        );

    \I__12603\ : LocalMux
    port map (
            O => \N__55525\,
            I => \c0.n21140\
        );

    \I__12602\ : LocalMux
    port map (
            O => \N__55522\,
            I => \c0.n21140\
        );

    \I__12601\ : InMux
    port map (
            O => \N__55513\,
            I => \N__55510\
        );

    \I__12600\ : LocalMux
    port map (
            O => \N__55510\,
            I => \N__55506\
        );

    \I__12599\ : InMux
    port map (
            O => \N__55509\,
            I => \N__55503\
        );

    \I__12598\ : Odrv4
    port map (
            O => \N__55506\,
            I => \c0.n22311\
        );

    \I__12597\ : LocalMux
    port map (
            O => \N__55503\,
            I => \c0.n22311\
        );

    \I__12596\ : InMux
    port map (
            O => \N__55498\,
            I => \N__55494\
        );

    \I__12595\ : InMux
    port map (
            O => \N__55497\,
            I => \N__55491\
        );

    \I__12594\ : LocalMux
    port map (
            O => \N__55494\,
            I => \c0.n22211\
        );

    \I__12593\ : LocalMux
    port map (
            O => \N__55491\,
            I => \c0.n22211\
        );

    \I__12592\ : InMux
    port map (
            O => \N__55486\,
            I => \N__55482\
        );

    \I__12591\ : InMux
    port map (
            O => \N__55485\,
            I => \N__55479\
        );

    \I__12590\ : LocalMux
    port map (
            O => \N__55482\,
            I => \N__55476\
        );

    \I__12589\ : LocalMux
    port map (
            O => \N__55479\,
            I => \c0.n23298\
        );

    \I__12588\ : Odrv4
    port map (
            O => \N__55476\,
            I => \c0.n23298\
        );

    \I__12587\ : InMux
    port map (
            O => \N__55471\,
            I => \N__55468\
        );

    \I__12586\ : LocalMux
    port map (
            O => \N__55468\,
            I => \N__55465\
        );

    \I__12585\ : Odrv4
    port map (
            O => \N__55465\,
            I => \c0.n7\
        );

    \I__12584\ : CascadeMux
    port map (
            O => \N__55462\,
            I => \c0.n23298_cascade_\
        );

    \I__12583\ : InMux
    port map (
            O => \N__55459\,
            I => \N__55456\
        );

    \I__12582\ : LocalMux
    port map (
            O => \N__55456\,
            I => \N__55453\
        );

    \I__12581\ : Span4Mux_h
    port map (
            O => \N__55453\,
            I => \N__55450\
        );

    \I__12580\ : Odrv4
    port map (
            O => \N__55450\,
            I => \c0.n45_adj_4486\
        );

    \I__12579\ : InMux
    port map (
            O => \N__55447\,
            I => \N__55444\
        );

    \I__12578\ : LocalMux
    port map (
            O => \N__55444\,
            I => \c0.n22100\
        );

    \I__12577\ : CascadeMux
    port map (
            O => \N__55441\,
            I => \c0.n21054_cascade_\
        );

    \I__12576\ : InMux
    port map (
            O => \N__55438\,
            I => \N__55435\
        );

    \I__12575\ : LocalMux
    port map (
            O => \N__55435\,
            I => \c0.n21043\
        );

    \I__12574\ : InMux
    port map (
            O => \N__55432\,
            I => \N__55426\
        );

    \I__12573\ : InMux
    port map (
            O => \N__55431\,
            I => \N__55421\
        );

    \I__12572\ : InMux
    port map (
            O => \N__55430\,
            I => \N__55421\
        );

    \I__12571\ : CascadeMux
    port map (
            O => \N__55429\,
            I => \N__55418\
        );

    \I__12570\ : LocalMux
    port map (
            O => \N__55426\,
            I => \N__55412\
        );

    \I__12569\ : LocalMux
    port map (
            O => \N__55421\,
            I => \N__55412\
        );

    \I__12568\ : InMux
    port map (
            O => \N__55418\,
            I => \N__55409\
        );

    \I__12567\ : InMux
    port map (
            O => \N__55417\,
            I => \N__55406\
        );

    \I__12566\ : Span4Mux_h
    port map (
            O => \N__55412\,
            I => \N__55403\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__55409\,
            I => \c0.data_in_frame_17_3\
        );

    \I__12564\ : LocalMux
    port map (
            O => \N__55406\,
            I => \c0.data_in_frame_17_3\
        );

    \I__12563\ : Odrv4
    port map (
            O => \N__55403\,
            I => \c0.data_in_frame_17_3\
        );

    \I__12562\ : InMux
    port map (
            O => \N__55396\,
            I => \N__55389\
        );

    \I__12561\ : InMux
    port map (
            O => \N__55395\,
            I => \N__55389\
        );

    \I__12560\ : InMux
    port map (
            O => \N__55394\,
            I => \N__55386\
        );

    \I__12559\ : LocalMux
    port map (
            O => \N__55389\,
            I => \N__55382\
        );

    \I__12558\ : LocalMux
    port map (
            O => \N__55386\,
            I => \N__55379\
        );

    \I__12557\ : InMux
    port map (
            O => \N__55385\,
            I => \N__55376\
        );

    \I__12556\ : Span4Mux_v
    port map (
            O => \N__55382\,
            I => \N__55372\
        );

    \I__12555\ : Span4Mux_h
    port map (
            O => \N__55379\,
            I => \N__55367\
        );

    \I__12554\ : LocalMux
    port map (
            O => \N__55376\,
            I => \N__55367\
        );

    \I__12553\ : InMux
    port map (
            O => \N__55375\,
            I => \N__55364\
        );

    \I__12552\ : Span4Mux_h
    port map (
            O => \N__55372\,
            I => \N__55361\
        );

    \I__12551\ : Span4Mux_h
    port map (
            O => \N__55367\,
            I => \N__55358\
        );

    \I__12550\ : LocalMux
    port map (
            O => \N__55364\,
            I => \c0.data_in_frame_17_4\
        );

    \I__12549\ : Odrv4
    port map (
            O => \N__55361\,
            I => \c0.data_in_frame_17_4\
        );

    \I__12548\ : Odrv4
    port map (
            O => \N__55358\,
            I => \c0.data_in_frame_17_4\
        );

    \I__12547\ : InMux
    port map (
            O => \N__55351\,
            I => \N__55345\
        );

    \I__12546\ : InMux
    port map (
            O => \N__55350\,
            I => \N__55345\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__55345\,
            I => \N__55342\
        );

    \I__12544\ : Odrv4
    port map (
            O => \N__55342\,
            I => \c0.n22480\
        );

    \I__12543\ : InMux
    port map (
            O => \N__55339\,
            I => \N__55335\
        );

    \I__12542\ : CascadeMux
    port map (
            O => \N__55338\,
            I => \N__55332\
        );

    \I__12541\ : LocalMux
    port map (
            O => \N__55335\,
            I => \N__55329\
        );

    \I__12540\ : InMux
    port map (
            O => \N__55332\,
            I => \N__55323\
        );

    \I__12539\ : Span4Mux_h
    port map (
            O => \N__55329\,
            I => \N__55320\
        );

    \I__12538\ : InMux
    port map (
            O => \N__55328\,
            I => \N__55317\
        );

    \I__12537\ : InMux
    port map (
            O => \N__55327\,
            I => \N__55312\
        );

    \I__12536\ : InMux
    port map (
            O => \N__55326\,
            I => \N__55312\
        );

    \I__12535\ : LocalMux
    port map (
            O => \N__55323\,
            I => \c0.data_in_frame_17_5\
        );

    \I__12534\ : Odrv4
    port map (
            O => \N__55320\,
            I => \c0.data_in_frame_17_5\
        );

    \I__12533\ : LocalMux
    port map (
            O => \N__55317\,
            I => \c0.data_in_frame_17_5\
        );

    \I__12532\ : LocalMux
    port map (
            O => \N__55312\,
            I => \c0.data_in_frame_17_5\
        );

    \I__12531\ : InMux
    port map (
            O => \N__55303\,
            I => \N__55299\
        );

    \I__12530\ : InMux
    port map (
            O => \N__55302\,
            I => \N__55296\
        );

    \I__12529\ : LocalMux
    port map (
            O => \N__55299\,
            I => \N__55293\
        );

    \I__12528\ : LocalMux
    port map (
            O => \N__55296\,
            I => \N__55290\
        );

    \I__12527\ : Span4Mux_v
    port map (
            O => \N__55293\,
            I => \N__55287\
        );

    \I__12526\ : Odrv4
    port map (
            O => \N__55290\,
            I => \c0.n13719\
        );

    \I__12525\ : Odrv4
    port map (
            O => \N__55287\,
            I => \c0.n13719\
        );

    \I__12524\ : InMux
    port map (
            O => \N__55282\,
            I => \N__55279\
        );

    \I__12523\ : LocalMux
    port map (
            O => \N__55279\,
            I => \c0.n18\
        );

    \I__12522\ : CascadeMux
    port map (
            O => \N__55276\,
            I => \N__55273\
        );

    \I__12521\ : InMux
    port map (
            O => \N__55273\,
            I => \N__55270\
        );

    \I__12520\ : LocalMux
    port map (
            O => \N__55270\,
            I => \N__55267\
        );

    \I__12519\ : Span4Mux_h
    port map (
            O => \N__55267\,
            I => \N__55264\
        );

    \I__12518\ : Odrv4
    port map (
            O => \N__55264\,
            I => \c0.n22349\
        );

    \I__12517\ : InMux
    port map (
            O => \N__55261\,
            I => \N__55258\
        );

    \I__12516\ : LocalMux
    port map (
            O => \N__55258\,
            I => \c0.n30\
        );

    \I__12515\ : InMux
    port map (
            O => \N__55255\,
            I => \N__55252\
        );

    \I__12514\ : LocalMux
    port map (
            O => \N__55252\,
            I => \c0.n22\
        );

    \I__12513\ : InMux
    port map (
            O => \N__55249\,
            I => \N__55246\
        );

    \I__12512\ : LocalMux
    port map (
            O => \N__55246\,
            I => \N__55243\
        );

    \I__12511\ : Odrv4
    port map (
            O => \N__55243\,
            I => \c0.n7_adj_4235\
        );

    \I__12510\ : InMux
    port map (
            O => \N__55240\,
            I => \N__55237\
        );

    \I__12509\ : LocalMux
    port map (
            O => \N__55237\,
            I => \N__55234\
        );

    \I__12508\ : Odrv4
    port map (
            O => \N__55234\,
            I => \c0.n8_adj_4236\
        );

    \I__12507\ : CascadeMux
    port map (
            O => \N__55231\,
            I => \c0.n20203_cascade_\
        );

    \I__12506\ : InMux
    port map (
            O => \N__55228\,
            I => \N__55225\
        );

    \I__12505\ : LocalMux
    port map (
            O => \N__55225\,
            I => \N__55222\
        );

    \I__12504\ : Odrv4
    port map (
            O => \N__55222\,
            I => \c0.n21120\
        );

    \I__12503\ : InMux
    port map (
            O => \N__55219\,
            I => \N__55214\
        );

    \I__12502\ : CascadeMux
    port map (
            O => \N__55218\,
            I => \N__55211\
        );

    \I__12501\ : InMux
    port map (
            O => \N__55217\,
            I => \N__55207\
        );

    \I__12500\ : LocalMux
    port map (
            O => \N__55214\,
            I => \N__55204\
        );

    \I__12499\ : InMux
    port map (
            O => \N__55211\,
            I => \N__55201\
        );

    \I__12498\ : InMux
    port map (
            O => \N__55210\,
            I => \N__55198\
        );

    \I__12497\ : LocalMux
    port map (
            O => \N__55207\,
            I => \N__55195\
        );

    \I__12496\ : Sp12to4
    port map (
            O => \N__55204\,
            I => \N__55192\
        );

    \I__12495\ : LocalMux
    port map (
            O => \N__55201\,
            I => \c0.data_in_frame_15_2\
        );

    \I__12494\ : LocalMux
    port map (
            O => \N__55198\,
            I => \c0.data_in_frame_15_2\
        );

    \I__12493\ : Odrv4
    port map (
            O => \N__55195\,
            I => \c0.data_in_frame_15_2\
        );

    \I__12492\ : Odrv12
    port map (
            O => \N__55192\,
            I => \c0.data_in_frame_15_2\
        );

    \I__12491\ : InMux
    port map (
            O => \N__55183\,
            I => \N__55180\
        );

    \I__12490\ : LocalMux
    port map (
            O => \N__55180\,
            I => \N__55177\
        );

    \I__12489\ : Span4Mux_v
    port map (
            O => \N__55177\,
            I => \N__55174\
        );

    \I__12488\ : Odrv4
    port map (
            O => \N__55174\,
            I => \c0.n22242\
        );

    \I__12487\ : CascadeMux
    port map (
            O => \N__55171\,
            I => \N__55168\
        );

    \I__12486\ : InMux
    port map (
            O => \N__55168\,
            I => \N__55165\
        );

    \I__12485\ : LocalMux
    port map (
            O => \N__55165\,
            I => \N__55162\
        );

    \I__12484\ : Span4Mux_h
    port map (
            O => \N__55162\,
            I => \N__55159\
        );

    \I__12483\ : Odrv4
    port map (
            O => \N__55159\,
            I => \c0.n20402\
        );

    \I__12482\ : InMux
    port map (
            O => \N__55156\,
            I => \N__55152\
        );

    \I__12481\ : InMux
    port map (
            O => \N__55155\,
            I => \N__55149\
        );

    \I__12480\ : LocalMux
    port map (
            O => \N__55152\,
            I => \c0.n20196\
        );

    \I__12479\ : LocalMux
    port map (
            O => \N__55149\,
            I => \c0.n20196\
        );

    \I__12478\ : CascadeMux
    port map (
            O => \N__55144\,
            I => \c0.n13719_cascade_\
        );

    \I__12477\ : InMux
    port map (
            O => \N__55141\,
            I => \N__55138\
        );

    \I__12476\ : LocalMux
    port map (
            O => \N__55138\,
            I => \N__55134\
        );

    \I__12475\ : InMux
    port map (
            O => \N__55137\,
            I => \N__55131\
        );

    \I__12474\ : Odrv4
    port map (
            O => \N__55134\,
            I => \c0.n22221\
        );

    \I__12473\ : LocalMux
    port map (
            O => \N__55131\,
            I => \c0.n22221\
        );

    \I__12472\ : InMux
    port map (
            O => \N__55126\,
            I => \N__55123\
        );

    \I__12471\ : LocalMux
    port map (
            O => \N__55123\,
            I => \N__55120\
        );

    \I__12470\ : Span4Mux_h
    port map (
            O => \N__55120\,
            I => \N__55115\
        );

    \I__12469\ : InMux
    port map (
            O => \N__55119\,
            I => \N__55112\
        );

    \I__12468\ : InMux
    port map (
            O => \N__55118\,
            I => \N__55109\
        );

    \I__12467\ : Odrv4
    port map (
            O => \N__55115\,
            I => \c0.n13786\
        );

    \I__12466\ : LocalMux
    port map (
            O => \N__55112\,
            I => \c0.n13786\
        );

    \I__12465\ : LocalMux
    port map (
            O => \N__55109\,
            I => \c0.n13786\
        );

    \I__12464\ : InMux
    port map (
            O => \N__55102\,
            I => \N__55098\
        );

    \I__12463\ : InMux
    port map (
            O => \N__55101\,
            I => \N__55092\
        );

    \I__12462\ : LocalMux
    port map (
            O => \N__55098\,
            I => \N__55089\
        );

    \I__12461\ : InMux
    port map (
            O => \N__55097\,
            I => \N__55084\
        );

    \I__12460\ : InMux
    port map (
            O => \N__55096\,
            I => \N__55084\
        );

    \I__12459\ : InMux
    port map (
            O => \N__55095\,
            I => \N__55081\
        );

    \I__12458\ : LocalMux
    port map (
            O => \N__55092\,
            I => \N__55078\
        );

    \I__12457\ : Span4Mux_v
    port map (
            O => \N__55089\,
            I => \N__55073\
        );

    \I__12456\ : LocalMux
    port map (
            O => \N__55084\,
            I => \N__55073\
        );

    \I__12455\ : LocalMux
    port map (
            O => \N__55081\,
            I => data_in_frame_14_6
        );

    \I__12454\ : Odrv12
    port map (
            O => \N__55078\,
            I => data_in_frame_14_6
        );

    \I__12453\ : Odrv4
    port map (
            O => \N__55073\,
            I => data_in_frame_14_6
        );

    \I__12452\ : InMux
    port map (
            O => \N__55066\,
            I => \N__55061\
        );

    \I__12451\ : CascadeMux
    port map (
            O => \N__55065\,
            I => \N__55058\
        );

    \I__12450\ : InMux
    port map (
            O => \N__55064\,
            I => \N__55054\
        );

    \I__12449\ : LocalMux
    port map (
            O => \N__55061\,
            I => \N__55051\
        );

    \I__12448\ : InMux
    port map (
            O => \N__55058\,
            I => \N__55048\
        );

    \I__12447\ : InMux
    port map (
            O => \N__55057\,
            I => \N__55044\
        );

    \I__12446\ : LocalMux
    port map (
            O => \N__55054\,
            I => \N__55037\
        );

    \I__12445\ : Span4Mux_v
    port map (
            O => \N__55051\,
            I => \N__55037\
        );

    \I__12444\ : LocalMux
    port map (
            O => \N__55048\,
            I => \N__55037\
        );

    \I__12443\ : InMux
    port map (
            O => \N__55047\,
            I => \N__55034\
        );

    \I__12442\ : LocalMux
    port map (
            O => \N__55044\,
            I => data_in_frame_14_7
        );

    \I__12441\ : Odrv4
    port map (
            O => \N__55037\,
            I => data_in_frame_14_7
        );

    \I__12440\ : LocalMux
    port map (
            O => \N__55034\,
            I => data_in_frame_14_7
        );

    \I__12439\ : CascadeMux
    port map (
            O => \N__55027\,
            I => \N__55024\
        );

    \I__12438\ : InMux
    port map (
            O => \N__55024\,
            I => \N__55021\
        );

    \I__12437\ : LocalMux
    port map (
            O => \N__55021\,
            I => \c0.n5996\
        );

    \I__12436\ : CascadeMux
    port map (
            O => \N__55018\,
            I => \c0.n20222_cascade_\
        );

    \I__12435\ : InMux
    port map (
            O => \N__55015\,
            I => \N__55012\
        );

    \I__12434\ : LocalMux
    port map (
            O => \N__55012\,
            I => \N__55008\
        );

    \I__12433\ : InMux
    port map (
            O => \N__55011\,
            I => \N__55005\
        );

    \I__12432\ : Span4Mux_h
    port map (
            O => \N__55008\,
            I => \N__55000\
        );

    \I__12431\ : LocalMux
    port map (
            O => \N__55005\,
            I => \N__55000\
        );

    \I__12430\ : Span4Mux_v
    port map (
            O => \N__55000\,
            I => \N__54996\
        );

    \I__12429\ : InMux
    port map (
            O => \N__54999\,
            I => \N__54993\
        );

    \I__12428\ : Sp12to4
    port map (
            O => \N__54996\,
            I => \N__54988\
        );

    \I__12427\ : LocalMux
    port map (
            O => \N__54993\,
            I => \N__54988\
        );

    \I__12426\ : Odrv12
    port map (
            O => \N__54988\,
            I => \c0.n13677\
        );

    \I__12425\ : CascadeMux
    port map (
            O => \N__54985\,
            I => \c0.n28_adj_4232_cascade_\
        );

    \I__12424\ : CascadeMux
    port map (
            O => \N__54982\,
            I => \c0.n32_cascade_\
        );

    \I__12423\ : InMux
    port map (
            O => \N__54979\,
            I => \N__54976\
        );

    \I__12422\ : LocalMux
    port map (
            O => \N__54976\,
            I => \N__54973\
        );

    \I__12421\ : Odrv12
    port map (
            O => \N__54973\,
            I => \c0.n29_adj_4234\
        );

    \I__12420\ : InMux
    port map (
            O => \N__54970\,
            I => \N__54967\
        );

    \I__12419\ : LocalMux
    port map (
            O => \N__54967\,
            I => \N__54964\
        );

    \I__12418\ : Span4Mux_h
    port map (
            O => \N__54964\,
            I => \N__54961\
        );

    \I__12417\ : Odrv4
    port map (
            O => \N__54961\,
            I => \c0.n13681\
        );

    \I__12416\ : CascadeMux
    port map (
            O => \N__54958\,
            I => \c0.n21238_cascade_\
        );

    \I__12415\ : InMux
    port map (
            O => \N__54955\,
            I => \N__54952\
        );

    \I__12414\ : LocalMux
    port map (
            O => \N__54952\,
            I => \N__54948\
        );

    \I__12413\ : InMux
    port map (
            O => \N__54951\,
            I => \N__54945\
        );

    \I__12412\ : Span4Mux_h
    port map (
            O => \N__54948\,
            I => \N__54942\
        );

    \I__12411\ : LocalMux
    port map (
            O => \N__54945\,
            I => \c0.n21989\
        );

    \I__12410\ : Odrv4
    port map (
            O => \N__54942\,
            I => \c0.n21989\
        );

    \I__12409\ : InMux
    port map (
            O => \N__54937\,
            I => \N__54931\
        );

    \I__12408\ : InMux
    port map (
            O => \N__54936\,
            I => \N__54931\
        );

    \I__12407\ : LocalMux
    port map (
            O => \N__54931\,
            I => \c0.n21238\
        );

    \I__12406\ : InMux
    port map (
            O => \N__54928\,
            I => \N__54924\
        );

    \I__12405\ : InMux
    port map (
            O => \N__54927\,
            I => \N__54921\
        );

    \I__12404\ : LocalMux
    port map (
            O => \N__54924\,
            I => \N__54916\
        );

    \I__12403\ : LocalMux
    port map (
            O => \N__54921\,
            I => \N__54916\
        );

    \I__12402\ : Span4Mux_v
    port map (
            O => \N__54916\,
            I => \N__54913\
        );

    \I__12401\ : Odrv4
    port map (
            O => \N__54913\,
            I => \c0.n22430\
        );

    \I__12400\ : InMux
    port map (
            O => \N__54910\,
            I => \N__54907\
        );

    \I__12399\ : LocalMux
    port map (
            O => \N__54907\,
            I => \N__54903\
        );

    \I__12398\ : InMux
    port map (
            O => \N__54906\,
            I => \N__54900\
        );

    \I__12397\ : Odrv4
    port map (
            O => \N__54903\,
            I => \c0.n5810\
        );

    \I__12396\ : LocalMux
    port map (
            O => \N__54900\,
            I => \c0.n5810\
        );

    \I__12395\ : CascadeMux
    port map (
            O => \N__54895\,
            I => \N__54890\
        );

    \I__12394\ : InMux
    port map (
            O => \N__54894\,
            I => \N__54886\
        );

    \I__12393\ : CascadeMux
    port map (
            O => \N__54893\,
            I => \N__54883\
        );

    \I__12392\ : InMux
    port map (
            O => \N__54890\,
            I => \N__54880\
        );

    \I__12391\ : InMux
    port map (
            O => \N__54889\,
            I => \N__54877\
        );

    \I__12390\ : LocalMux
    port map (
            O => \N__54886\,
            I => \N__54874\
        );

    \I__12389\ : InMux
    port map (
            O => \N__54883\,
            I => \N__54871\
        );

    \I__12388\ : LocalMux
    port map (
            O => \N__54880\,
            I => \N__54866\
        );

    \I__12387\ : LocalMux
    port map (
            O => \N__54877\,
            I => \N__54866\
        );

    \I__12386\ : Odrv4
    port map (
            O => \N__54874\,
            I => \c0.data_in_frame_7_1\
        );

    \I__12385\ : LocalMux
    port map (
            O => \N__54871\,
            I => \c0.data_in_frame_7_1\
        );

    \I__12384\ : Odrv4
    port map (
            O => \N__54866\,
            I => \c0.data_in_frame_7_1\
        );

    \I__12383\ : InMux
    port map (
            O => \N__54859\,
            I => \N__54856\
        );

    \I__12382\ : LocalMux
    port map (
            O => \N__54856\,
            I => \c0.n6_adj_4273\
        );

    \I__12381\ : InMux
    port map (
            O => \N__54853\,
            I => \N__54850\
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__54850\,
            I => \c0.n22139\
        );

    \I__12379\ : CascadeMux
    port map (
            O => \N__54847\,
            I => \N__54844\
        );

    \I__12378\ : InMux
    port map (
            O => \N__54844\,
            I => \N__54841\
        );

    \I__12377\ : LocalMux
    port map (
            O => \N__54841\,
            I => \N__54838\
        );

    \I__12376\ : Span4Mux_h
    port map (
            O => \N__54838\,
            I => \N__54835\
        );

    \I__12375\ : Odrv4
    port map (
            O => \N__54835\,
            I => \c0.n6_adj_4243\
        );

    \I__12374\ : InMux
    port map (
            O => \N__54832\,
            I => \N__54829\
        );

    \I__12373\ : LocalMux
    port map (
            O => \N__54829\,
            I => \N__54825\
        );

    \I__12372\ : InMux
    port map (
            O => \N__54828\,
            I => \N__54822\
        );

    \I__12371\ : Span4Mux_v
    port map (
            O => \N__54825\,
            I => \N__54819\
        );

    \I__12370\ : LocalMux
    port map (
            O => \N__54822\,
            I => \N__54816\
        );

    \I__12369\ : Span4Mux_h
    port map (
            O => \N__54819\,
            I => \N__54812\
        );

    \I__12368\ : Span4Mux_v
    port map (
            O => \N__54816\,
            I => \N__54809\
        );

    \I__12367\ : InMux
    port map (
            O => \N__54815\,
            I => \N__54806\
        );

    \I__12366\ : Odrv4
    port map (
            O => \N__54812\,
            I => \c0.n13861\
        );

    \I__12365\ : Odrv4
    port map (
            O => \N__54809\,
            I => \c0.n13861\
        );

    \I__12364\ : LocalMux
    port map (
            O => \N__54806\,
            I => \c0.n13861\
        );

    \I__12363\ : CascadeMux
    port map (
            O => \N__54799\,
            I => \c0.n5813_cascade_\
        );

    \I__12362\ : InMux
    port map (
            O => \N__54796\,
            I => \N__54792\
        );

    \I__12361\ : InMux
    port map (
            O => \N__54795\,
            I => \N__54789\
        );

    \I__12360\ : LocalMux
    port map (
            O => \N__54792\,
            I => \N__54784\
        );

    \I__12359\ : LocalMux
    port map (
            O => \N__54789\,
            I => \N__54784\
        );

    \I__12358\ : Span4Mux_v
    port map (
            O => \N__54784\,
            I => \N__54781\
        );

    \I__12357\ : Odrv4
    port map (
            O => \N__54781\,
            I => \c0.n21967\
        );

    \I__12356\ : InMux
    port map (
            O => \N__54778\,
            I => \N__54773\
        );

    \I__12355\ : InMux
    port map (
            O => \N__54777\,
            I => \N__54768\
        );

    \I__12354\ : InMux
    port map (
            O => \N__54776\,
            I => \N__54768\
        );

    \I__12353\ : LocalMux
    port map (
            O => \N__54773\,
            I => \N__54761\
        );

    \I__12352\ : LocalMux
    port map (
            O => \N__54768\,
            I => \N__54761\
        );

    \I__12351\ : InMux
    port map (
            O => \N__54767\,
            I => \N__54756\
        );

    \I__12350\ : InMux
    port map (
            O => \N__54766\,
            I => \N__54756\
        );

    \I__12349\ : Odrv12
    port map (
            O => \N__54761\,
            I => \c0.n13237\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__54756\,
            I => \c0.n13237\
        );

    \I__12347\ : InMux
    port map (
            O => \N__54751\,
            I => \N__54748\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__54748\,
            I => \N__54743\
        );

    \I__12345\ : InMux
    port map (
            O => \N__54747\,
            I => \N__54740\
        );

    \I__12344\ : InMux
    port map (
            O => \N__54746\,
            I => \N__54737\
        );

    \I__12343\ : Span4Mux_h
    port map (
            O => \N__54743\,
            I => \N__54734\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__54740\,
            I => \N__54731\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__54737\,
            I => \N__54726\
        );

    \I__12340\ : Span4Mux_v
    port map (
            O => \N__54734\,
            I => \N__54726\
        );

    \I__12339\ : Span4Mux_v
    port map (
            O => \N__54731\,
            I => \N__54723\
        );

    \I__12338\ : Odrv4
    port map (
            O => \N__54726\,
            I => \c0.data_in_frame_7_6\
        );

    \I__12337\ : Odrv4
    port map (
            O => \N__54723\,
            I => \c0.data_in_frame_7_6\
        );

    \I__12336\ : InMux
    port map (
            O => \N__54718\,
            I => \N__54715\
        );

    \I__12335\ : LocalMux
    port map (
            O => \N__54715\,
            I => \N__54711\
        );

    \I__12334\ : InMux
    port map (
            O => \N__54714\,
            I => \N__54706\
        );

    \I__12333\ : Span4Mux_h
    port map (
            O => \N__54711\,
            I => \N__54703\
        );

    \I__12332\ : InMux
    port map (
            O => \N__54710\,
            I => \N__54700\
        );

    \I__12331\ : InMux
    port map (
            O => \N__54709\,
            I => \N__54697\
        );

    \I__12330\ : LocalMux
    port map (
            O => \N__54706\,
            I => \c0.data_in_frame_10_0\
        );

    \I__12329\ : Odrv4
    port map (
            O => \N__54703\,
            I => \c0.data_in_frame_10_0\
        );

    \I__12328\ : LocalMux
    port map (
            O => \N__54700\,
            I => \c0.data_in_frame_10_0\
        );

    \I__12327\ : LocalMux
    port map (
            O => \N__54697\,
            I => \c0.data_in_frame_10_0\
        );

    \I__12326\ : CascadeMux
    port map (
            O => \N__54688\,
            I => \c0.n10_adj_4245_cascade_\
        );

    \I__12325\ : InMux
    port map (
            O => \N__54685\,
            I => \N__54679\
        );

    \I__12324\ : InMux
    port map (
            O => \N__54684\,
            I => \N__54676\
        );

    \I__12323\ : InMux
    port map (
            O => \N__54683\,
            I => \N__54673\
        );

    \I__12322\ : InMux
    port map (
            O => \N__54682\,
            I => \N__54670\
        );

    \I__12321\ : LocalMux
    port map (
            O => \N__54679\,
            I => \N__54667\
        );

    \I__12320\ : LocalMux
    port map (
            O => \N__54676\,
            I => \N__54664\
        );

    \I__12319\ : LocalMux
    port map (
            O => \N__54673\,
            I => \N__54660\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__54670\,
            I => \N__54657\
        );

    \I__12317\ : Span4Mux_h
    port map (
            O => \N__54667\,
            I => \N__54654\
        );

    \I__12316\ : Span4Mux_v
    port map (
            O => \N__54664\,
            I => \N__54651\
        );

    \I__12315\ : InMux
    port map (
            O => \N__54663\,
            I => \N__54648\
        );

    \I__12314\ : Span4Mux_h
    port map (
            O => \N__54660\,
            I => \N__54643\
        );

    \I__12313\ : Span4Mux_v
    port map (
            O => \N__54657\,
            I => \N__54643\
        );

    \I__12312\ : Odrv4
    port map (
            O => \N__54654\,
            I => \c0.n13099\
        );

    \I__12311\ : Odrv4
    port map (
            O => \N__54651\,
            I => \c0.n13099\
        );

    \I__12310\ : LocalMux
    port map (
            O => \N__54648\,
            I => \c0.n13099\
        );

    \I__12309\ : Odrv4
    port map (
            O => \N__54643\,
            I => \c0.n13099\
        );

    \I__12308\ : InMux
    port map (
            O => \N__54634\,
            I => \N__54630\
        );

    \I__12307\ : CascadeMux
    port map (
            O => \N__54633\,
            I => \N__54627\
        );

    \I__12306\ : LocalMux
    port map (
            O => \N__54630\,
            I => \N__54623\
        );

    \I__12305\ : InMux
    port map (
            O => \N__54627\,
            I => \N__54618\
        );

    \I__12304\ : InMux
    port map (
            O => \N__54626\,
            I => \N__54618\
        );

    \I__12303\ : Odrv4
    port map (
            O => \N__54623\,
            I => \c0.data_in_frame_9_1\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__54618\,
            I => \c0.data_in_frame_9_1\
        );

    \I__12301\ : InMux
    port map (
            O => \N__54613\,
            I => \N__54610\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__54610\,
            I => \N__54607\
        );

    \I__12299\ : Span4Mux_v
    port map (
            O => \N__54607\,
            I => \N__54604\
        );

    \I__12298\ : Odrv4
    port map (
            O => \N__54604\,
            I => \c0.n14037\
        );

    \I__12297\ : InMux
    port map (
            O => \N__54601\,
            I => \N__54595\
        );

    \I__12296\ : InMux
    port map (
            O => \N__54600\,
            I => \N__54595\
        );

    \I__12295\ : LocalMux
    port map (
            O => \N__54595\,
            I => \c0.n22233\
        );

    \I__12294\ : CascadeMux
    port map (
            O => \N__54592\,
            I => \N__54589\
        );

    \I__12293\ : InMux
    port map (
            O => \N__54589\,
            I => \N__54584\
        );

    \I__12292\ : InMux
    port map (
            O => \N__54588\,
            I => \N__54581\
        );

    \I__12291\ : InMux
    port map (
            O => \N__54587\,
            I => \N__54578\
        );

    \I__12290\ : LocalMux
    port map (
            O => \N__54584\,
            I => \c0.data_in_frame_11_3\
        );

    \I__12289\ : LocalMux
    port map (
            O => \N__54581\,
            I => \c0.data_in_frame_11_3\
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__54578\,
            I => \c0.data_in_frame_11_3\
        );

    \I__12287\ : InMux
    port map (
            O => \N__54571\,
            I => \N__54568\
        );

    \I__12286\ : LocalMux
    port map (
            O => \N__54568\,
            I => \c0.n10_adj_4274\
        );

    \I__12285\ : InMux
    port map (
            O => \N__54565\,
            I => \N__54562\
        );

    \I__12284\ : LocalMux
    port map (
            O => \N__54562\,
            I => \N__54558\
        );

    \I__12283\ : InMux
    port map (
            O => \N__54561\,
            I => \N__54555\
        );

    \I__12282\ : Span4Mux_h
    port map (
            O => \N__54558\,
            I => \N__54552\
        );

    \I__12281\ : LocalMux
    port map (
            O => \N__54555\,
            I => \N__54549\
        );

    \I__12280\ : Odrv4
    port map (
            O => \N__54552\,
            I => \c0.n22108\
        );

    \I__12279\ : Odrv4
    port map (
            O => \N__54549\,
            I => \c0.n22108\
        );

    \I__12278\ : CascadeMux
    port map (
            O => \N__54544\,
            I => \c0.n4_adj_4240_cascade_\
        );

    \I__12277\ : InMux
    port map (
            O => \N__54541\,
            I => \N__54538\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__54538\,
            I => \N__54535\
        );

    \I__12275\ : Odrv4
    port map (
            O => \N__54535\,
            I => \c0.n22060\
        );

    \I__12274\ : CascadeMux
    port map (
            O => \N__54532\,
            I => \c0.n6_adj_4244_cascade_\
        );

    \I__12273\ : InMux
    port map (
            O => \N__54529\,
            I => \N__54525\
        );

    \I__12272\ : InMux
    port map (
            O => \N__54528\,
            I => \N__54522\
        );

    \I__12271\ : LocalMux
    port map (
            O => \N__54525\,
            I => \N__54519\
        );

    \I__12270\ : LocalMux
    port map (
            O => \N__54522\,
            I => \c0.n21097\
        );

    \I__12269\ : Odrv4
    port map (
            O => \N__54519\,
            I => \c0.n21097\
        );

    \I__12268\ : CascadeMux
    port map (
            O => \N__54514\,
            I => \c0.n20240_cascade_\
        );

    \I__12267\ : InMux
    port map (
            O => \N__54511\,
            I => \N__54508\
        );

    \I__12266\ : LocalMux
    port map (
            O => \N__54508\,
            I => \N__54504\
        );

    \I__12265\ : CascadeMux
    port map (
            O => \N__54507\,
            I => \N__54501\
        );

    \I__12264\ : Span4Mux_h
    port map (
            O => \N__54504\,
            I => \N__54497\
        );

    \I__12263\ : InMux
    port map (
            O => \N__54501\,
            I => \N__54494\
        );

    \I__12262\ : InMux
    port map (
            O => \N__54500\,
            I => \N__54491\
        );

    \I__12261\ : Span4Mux_v
    port map (
            O => \N__54497\,
            I => \N__54488\
        );

    \I__12260\ : LocalMux
    port map (
            O => \N__54494\,
            I => \c0.data_in_frame_15_0\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__54491\,
            I => \c0.data_in_frame_15_0\
        );

    \I__12258\ : Odrv4
    port map (
            O => \N__54488\,
            I => \c0.data_in_frame_15_0\
        );

    \I__12257\ : CascadeMux
    port map (
            O => \N__54481\,
            I => \c0.n22385_cascade_\
        );

    \I__12256\ : CascadeMux
    port map (
            O => \N__54478\,
            I => \N__54474\
        );

    \I__12255\ : InMux
    port map (
            O => \N__54477\,
            I => \N__54471\
        );

    \I__12254\ : InMux
    port map (
            O => \N__54474\,
            I => \N__54468\
        );

    \I__12253\ : LocalMux
    port map (
            O => \N__54471\,
            I => \N__54464\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__54468\,
            I => \N__54461\
        );

    \I__12251\ : InMux
    port map (
            O => \N__54467\,
            I => \N__54458\
        );

    \I__12250\ : Span4Mux_v
    port map (
            O => \N__54464\,
            I => \N__54453\
        );

    \I__12249\ : Span4Mux_h
    port map (
            O => \N__54461\,
            I => \N__54453\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__54458\,
            I => data_in_frame_14_5
        );

    \I__12247\ : Odrv4
    port map (
            O => \N__54453\,
            I => data_in_frame_14_5
        );

    \I__12246\ : InMux
    port map (
            O => \N__54448\,
            I => \N__54444\
        );

    \I__12245\ : InMux
    port map (
            O => \N__54447\,
            I => \N__54441\
        );

    \I__12244\ : LocalMux
    port map (
            O => \N__54444\,
            I => data_in_frame_14_3
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__54441\,
            I => data_in_frame_14_3
        );

    \I__12242\ : CascadeMux
    port map (
            O => \N__54436\,
            I => \N__54433\
        );

    \I__12241\ : InMux
    port map (
            O => \N__54433\,
            I => \N__54429\
        );

    \I__12240\ : InMux
    port map (
            O => \N__54432\,
            I => \N__54426\
        );

    \I__12239\ : LocalMux
    port map (
            O => \N__54429\,
            I => \c0.data_in_frame_4_0\
        );

    \I__12238\ : LocalMux
    port map (
            O => \N__54426\,
            I => \c0.data_in_frame_4_0\
        );

    \I__12237\ : InMux
    port map (
            O => \N__54421\,
            I => \N__54417\
        );

    \I__12236\ : InMux
    port map (
            O => \N__54420\,
            I => \N__54414\
        );

    \I__12235\ : LocalMux
    port map (
            O => \N__54417\,
            I => \N__54411\
        );

    \I__12234\ : LocalMux
    port map (
            O => \N__54414\,
            I => \N__54408\
        );

    \I__12233\ : Span4Mux_v
    port map (
            O => \N__54411\,
            I => \N__54404\
        );

    \I__12232\ : Span4Mux_v
    port map (
            O => \N__54408\,
            I => \N__54401\
        );

    \I__12231\ : CascadeMux
    port map (
            O => \N__54407\,
            I => \N__54396\
        );

    \I__12230\ : Span4Mux_v
    port map (
            O => \N__54404\,
            I => \N__54390\
        );

    \I__12229\ : Span4Mux_h
    port map (
            O => \N__54401\,
            I => \N__54390\
        );

    \I__12228\ : InMux
    port map (
            O => \N__54400\,
            I => \N__54387\
        );

    \I__12227\ : InMux
    port map (
            O => \N__54399\,
            I => \N__54384\
        );

    \I__12226\ : InMux
    port map (
            O => \N__54396\,
            I => \N__54379\
        );

    \I__12225\ : InMux
    port map (
            O => \N__54395\,
            I => \N__54379\
        );

    \I__12224\ : Sp12to4
    port map (
            O => \N__54390\,
            I => \N__54374\
        );

    \I__12223\ : LocalMux
    port map (
            O => \N__54387\,
            I => \N__54374\
        );

    \I__12222\ : LocalMux
    port map (
            O => \N__54384\,
            I => data_in_frame_1_4
        );

    \I__12221\ : LocalMux
    port map (
            O => \N__54379\,
            I => data_in_frame_1_4
        );

    \I__12220\ : Odrv12
    port map (
            O => \N__54374\,
            I => data_in_frame_1_4
        );

    \I__12219\ : InMux
    port map (
            O => \N__54367\,
            I => \N__54364\
        );

    \I__12218\ : LocalMux
    port map (
            O => \N__54364\,
            I => \N__54360\
        );

    \I__12217\ : InMux
    port map (
            O => \N__54363\,
            I => \N__54357\
        );

    \I__12216\ : Span4Mux_v
    port map (
            O => \N__54360\,
            I => \N__54352\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__54357\,
            I => \N__54352\
        );

    \I__12214\ : Span4Mux_h
    port map (
            O => \N__54352\,
            I => \N__54349\
        );

    \I__12213\ : Odrv4
    port map (
            O => \N__54349\,
            I => \c0.n21797\
        );

    \I__12212\ : CascadeMux
    port map (
            O => \N__54346\,
            I => \r_SM_Main_2_N_3681_2_cascade_\
        );

    \I__12211\ : CascadeMux
    port map (
            O => \N__54343\,
            I => \N__54340\
        );

    \I__12210\ : InMux
    port map (
            O => \N__54340\,
            I => \N__54337\
        );

    \I__12209\ : LocalMux
    port map (
            O => \N__54337\,
            I => \N__54334\
        );

    \I__12208\ : Span12Mux_h
    port map (
            O => \N__54334\,
            I => \N__54331\
        );

    \I__12207\ : Span12Mux_v
    port map (
            O => \N__54331\,
            I => \N__54328\
        );

    \I__12206\ : Span12Mux_h
    port map (
            O => \N__54328\,
            I => \N__54325\
        );

    \I__12205\ : Odrv12
    port map (
            O => \N__54325\,
            I => n14283
        );

    \I__12204\ : InMux
    port map (
            O => \N__54322\,
            I => \N__54316\
        );

    \I__12203\ : InMux
    port map (
            O => \N__54321\,
            I => \N__54313\
        );

    \I__12202\ : InMux
    port map (
            O => \N__54320\,
            I => \N__54308\
        );

    \I__12201\ : InMux
    port map (
            O => \N__54319\,
            I => \N__54308\
        );

    \I__12200\ : LocalMux
    port map (
            O => \N__54316\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__12199\ : LocalMux
    port map (
            O => \N__54313\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__12198\ : LocalMux
    port map (
            O => \N__54308\,
            I => \c0.rx.r_Clock_Count_4\
        );

    \I__12197\ : InMux
    port map (
            O => \N__54301\,
            I => \N__54297\
        );

    \I__12196\ : InMux
    port map (
            O => \N__54300\,
            I => \N__54294\
        );

    \I__12195\ : LocalMux
    port map (
            O => \N__54297\,
            I => \c0.rx.n18655\
        );

    \I__12194\ : LocalMux
    port map (
            O => \N__54294\,
            I => \c0.rx.n18655\
        );

    \I__12193\ : CascadeMux
    port map (
            O => \N__54289\,
            I => \N__54286\
        );

    \I__12192\ : InMux
    port map (
            O => \N__54286\,
            I => \N__54280\
        );

    \I__12191\ : InMux
    port map (
            O => \N__54285\,
            I => \N__54277\
        );

    \I__12190\ : InMux
    port map (
            O => \N__54284\,
            I => \N__54274\
        );

    \I__12189\ : InMux
    port map (
            O => \N__54283\,
            I => \N__54271\
        );

    \I__12188\ : LocalMux
    port map (
            O => \N__54280\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__12187\ : LocalMux
    port map (
            O => \N__54277\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__12186\ : LocalMux
    port map (
            O => \N__54274\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__12185\ : LocalMux
    port map (
            O => \N__54271\,
            I => \c0.rx.r_Clock_Count_0\
        );

    \I__12184\ : InMux
    port map (
            O => \N__54262\,
            I => \N__54258\
        );

    \I__12183\ : InMux
    port map (
            O => \N__54261\,
            I => \N__54255\
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__54258\,
            I => \c0.rx.n80\
        );

    \I__12181\ : LocalMux
    port map (
            O => \N__54255\,
            I => \c0.rx.n80\
        );

    \I__12180\ : SRMux
    port map (
            O => \N__54250\,
            I => \N__54247\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__54247\,
            I => \N__54244\
        );

    \I__12178\ : Span4Mux_h
    port map (
            O => \N__54244\,
            I => \N__54241\
        );

    \I__12177\ : Span4Mux_h
    port map (
            O => \N__54241\,
            I => \N__54238\
        );

    \I__12176\ : Span4Mux_v
    port map (
            O => \N__54238\,
            I => \N__54235\
        );

    \I__12175\ : Odrv4
    port map (
            O => \N__54235\,
            I => \c0.rx.n21783\
        );

    \I__12174\ : InMux
    port map (
            O => \N__54232\,
            I => \N__54229\
        );

    \I__12173\ : LocalMux
    port map (
            O => \N__54229\,
            I => \N__54226\
        );

    \I__12172\ : Span4Mux_v
    port map (
            O => \N__54226\,
            I => \N__54223\
        );

    \I__12171\ : Sp12to4
    port map (
            O => \N__54223\,
            I => \N__54220\
        );

    \I__12170\ : Span12Mux_h
    port map (
            O => \N__54220\,
            I => \N__54217\
        );

    \I__12169\ : Odrv12
    port map (
            O => \N__54217\,
            I => \c0.rx.r_Rx_Data_R\
        );

    \I__12168\ : InMux
    port map (
            O => \N__54214\,
            I => \N__54210\
        );

    \I__12167\ : CascadeMux
    port map (
            O => \N__54213\,
            I => \N__54207\
        );

    \I__12166\ : LocalMux
    port map (
            O => \N__54210\,
            I => \N__54204\
        );

    \I__12165\ : InMux
    port map (
            O => \N__54207\,
            I => \N__54201\
        );

    \I__12164\ : Span4Mux_v
    port map (
            O => \N__54204\,
            I => \N__54198\
        );

    \I__12163\ : LocalMux
    port map (
            O => \N__54201\,
            I => \c0.data_in_frame_12_6\
        );

    \I__12162\ : Odrv4
    port map (
            O => \N__54198\,
            I => \c0.data_in_frame_12_6\
        );

    \I__12161\ : InMux
    port map (
            O => \N__54193\,
            I => \N__54190\
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__54190\,
            I => \N__54185\
        );

    \I__12159\ : InMux
    port map (
            O => \N__54189\,
            I => \N__54180\
        );

    \I__12158\ : InMux
    port map (
            O => \N__54188\,
            I => \N__54180\
        );

    \I__12157\ : Odrv4
    port map (
            O => \N__54185\,
            I => \c0.data_in_frame_15_3\
        );

    \I__12156\ : LocalMux
    port map (
            O => \N__54180\,
            I => \c0.data_in_frame_15_3\
        );

    \I__12155\ : InMux
    port map (
            O => \N__54175\,
            I => \N__54171\
        );

    \I__12154\ : InMux
    port map (
            O => \N__54174\,
            I => \N__54168\
        );

    \I__12153\ : LocalMux
    port map (
            O => \N__54171\,
            I => \N__54165\
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__54168\,
            I => \N__54161\
        );

    \I__12151\ : Span4Mux_v
    port map (
            O => \N__54165\,
            I => \N__54158\
        );

    \I__12150\ : InMux
    port map (
            O => \N__54164\,
            I => \N__54155\
        );

    \I__12149\ : Odrv4
    port map (
            O => \N__54161\,
            I => \c0.n20927\
        );

    \I__12148\ : Odrv4
    port map (
            O => \N__54158\,
            I => \c0.n20927\
        );

    \I__12147\ : LocalMux
    port map (
            O => \N__54155\,
            I => \c0.n20927\
        );

    \I__12146\ : InMux
    port map (
            O => \N__54148\,
            I => \N__54145\
        );

    \I__12145\ : LocalMux
    port map (
            O => \N__54145\,
            I => \N__54142\
        );

    \I__12144\ : Odrv12
    port map (
            O => \N__54142\,
            I => \c0.n22119\
        );

    \I__12143\ : CascadeMux
    port map (
            O => \N__54139\,
            I => \c0.n21099_cascade_\
        );

    \I__12142\ : InMux
    port map (
            O => \N__54136\,
            I => \N__54132\
        );

    \I__12141\ : InMux
    port map (
            O => \N__54135\,
            I => \N__54127\
        );

    \I__12140\ : LocalMux
    port map (
            O => \N__54132\,
            I => \N__54124\
        );

    \I__12139\ : InMux
    port map (
            O => \N__54131\,
            I => \N__54119\
        );

    \I__12138\ : InMux
    port map (
            O => \N__54130\,
            I => \N__54119\
        );

    \I__12137\ : LocalMux
    port map (
            O => \N__54127\,
            I => \c0.n21160\
        );

    \I__12136\ : Odrv4
    port map (
            O => \N__54124\,
            I => \c0.n21160\
        );

    \I__12135\ : LocalMux
    port map (
            O => \N__54119\,
            I => \c0.n21160\
        );

    \I__12134\ : InMux
    port map (
            O => \N__54112\,
            I => \N__54108\
        );

    \I__12133\ : InMux
    port map (
            O => \N__54111\,
            I => \N__54105\
        );

    \I__12132\ : LocalMux
    port map (
            O => \N__54108\,
            I => \N__54100\
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__54105\,
            I => \N__54100\
        );

    \I__12130\ : Odrv4
    port map (
            O => \N__54100\,
            I => \c0.data_in_frame_29_6\
        );

    \I__12129\ : InMux
    port map (
            O => \N__54097\,
            I => \N__54094\
        );

    \I__12128\ : LocalMux
    port map (
            O => \N__54094\,
            I => \N__54090\
        );

    \I__12127\ : InMux
    port map (
            O => \N__54093\,
            I => \N__54087\
        );

    \I__12126\ : Span4Mux_h
    port map (
            O => \N__54090\,
            I => \N__54084\
        );

    \I__12125\ : LocalMux
    port map (
            O => \N__54087\,
            I => \c0.n63_adj_4293\
        );

    \I__12124\ : Odrv4
    port map (
            O => \N__54084\,
            I => \c0.n63_adj_4293\
        );

    \I__12123\ : CascadeMux
    port map (
            O => \N__54079\,
            I => \c0.n22148_cascade_\
        );

    \I__12122\ : InMux
    port map (
            O => \N__54076\,
            I => \N__54073\
        );

    \I__12121\ : LocalMux
    port map (
            O => \N__54073\,
            I => \c0.n21233\
        );

    \I__12120\ : InMux
    port map (
            O => \N__54070\,
            I => \N__54067\
        );

    \I__12119\ : LocalMux
    port map (
            O => \N__54067\,
            I => \N__54064\
        );

    \I__12118\ : Span4Mux_h
    port map (
            O => \N__54064\,
            I => \N__54061\
        );

    \I__12117\ : Odrv4
    port map (
            O => \N__54061\,
            I => \c0.n26_adj_4294\
        );

    \I__12116\ : CascadeMux
    port map (
            O => \N__54058\,
            I => \c0.rx.n12862_cascade_\
        );

    \I__12115\ : InMux
    port map (
            O => \N__54055\,
            I => \N__54051\
        );

    \I__12114\ : InMux
    port map (
            O => \N__54054\,
            I => \N__54048\
        );

    \I__12113\ : LocalMux
    port map (
            O => \N__54051\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__12112\ : LocalMux
    port map (
            O => \N__54048\,
            I => \c0.rx.r_Clock_Count_7\
        );

    \I__12111\ : InMux
    port map (
            O => \N__54043\,
            I => \N__54039\
        );

    \I__12110\ : InMux
    port map (
            O => \N__54042\,
            I => \N__54036\
        );

    \I__12109\ : LocalMux
    port map (
            O => \N__54039\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__12108\ : LocalMux
    port map (
            O => \N__54036\,
            I => \c0.rx.r_Clock_Count_5\
        );

    \I__12107\ : InMux
    port map (
            O => \N__54031\,
            I => \N__54027\
        );

    \I__12106\ : InMux
    port map (
            O => \N__54030\,
            I => \N__54024\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__54027\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__12104\ : LocalMux
    port map (
            O => \N__54024\,
            I => \c0.rx.r_Clock_Count_6\
        );

    \I__12103\ : CascadeMux
    port map (
            O => \N__54019\,
            I => \c0.rx.n80_cascade_\
        );

    \I__12102\ : InMux
    port map (
            O => \N__54016\,
            I => \N__54012\
        );

    \I__12101\ : InMux
    port map (
            O => \N__54015\,
            I => \N__54009\
        );

    \I__12100\ : LocalMux
    port map (
            O => \N__54012\,
            I => \N__54004\
        );

    \I__12099\ : LocalMux
    port map (
            O => \N__54009\,
            I => \N__54001\
        );

    \I__12098\ : InMux
    port map (
            O => \N__54008\,
            I => \N__53998\
        );

    \I__12097\ : InMux
    port map (
            O => \N__54007\,
            I => \N__53995\
        );

    \I__12096\ : Odrv4
    port map (
            O => \N__54004\,
            I => \c0.n13761\
        );

    \I__12095\ : Odrv4
    port map (
            O => \N__54001\,
            I => \c0.n13761\
        );

    \I__12094\ : LocalMux
    port map (
            O => \N__53998\,
            I => \c0.n13761\
        );

    \I__12093\ : LocalMux
    port map (
            O => \N__53995\,
            I => \c0.n13761\
        );

    \I__12092\ : InMux
    port map (
            O => \N__53986\,
            I => \N__53983\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__53983\,
            I => \c0.n22145\
        );

    \I__12090\ : InMux
    port map (
            O => \N__53980\,
            I => \N__53976\
        );

    \I__12089\ : InMux
    port map (
            O => \N__53979\,
            I => \N__53973\
        );

    \I__12088\ : LocalMux
    port map (
            O => \N__53976\,
            I => \c0.n21949\
        );

    \I__12087\ : LocalMux
    port map (
            O => \N__53973\,
            I => \c0.n21949\
        );

    \I__12086\ : CascadeMux
    port map (
            O => \N__53968\,
            I => \c0.n22145_cascade_\
        );

    \I__12085\ : InMux
    port map (
            O => \N__53965\,
            I => \N__53962\
        );

    \I__12084\ : LocalMux
    port map (
            O => \N__53962\,
            I => \c0.n10_adj_4297\
        );

    \I__12083\ : CascadeMux
    port map (
            O => \N__53959\,
            I => \c0.n23335_cascade_\
        );

    \I__12082\ : CascadeMux
    port map (
            O => \N__53956\,
            I => \N__53953\
        );

    \I__12081\ : InMux
    port map (
            O => \N__53953\,
            I => \N__53950\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__53950\,
            I => \N__53947\
        );

    \I__12079\ : Span4Mux_v
    port map (
            O => \N__53947\,
            I => \N__53944\
        );

    \I__12078\ : Odrv4
    port map (
            O => \N__53944\,
            I => \c0.n21_adj_4300\
        );

    \I__12077\ : CascadeMux
    port map (
            O => \N__53941\,
            I => \N__53937\
        );

    \I__12076\ : CascadeMux
    port map (
            O => \N__53940\,
            I => \N__53934\
        );

    \I__12075\ : InMux
    port map (
            O => \N__53937\,
            I => \N__53931\
        );

    \I__12074\ : InMux
    port map (
            O => \N__53934\,
            I => \N__53928\
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__53931\,
            I => \N__53925\
        );

    \I__12072\ : LocalMux
    port map (
            O => \N__53928\,
            I => \c0.data_in_frame_29_3\
        );

    \I__12071\ : Odrv4
    port map (
            O => \N__53925\,
            I => \c0.data_in_frame_29_3\
        );

    \I__12070\ : CascadeMux
    port map (
            O => \N__53920\,
            I => \N__53917\
        );

    \I__12069\ : InMux
    port map (
            O => \N__53917\,
            I => \N__53913\
        );

    \I__12068\ : InMux
    port map (
            O => \N__53916\,
            I => \N__53910\
        );

    \I__12067\ : LocalMux
    port map (
            O => \N__53913\,
            I => \c0.data_in_frame_28_0\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__53910\,
            I => \c0.data_in_frame_28_0\
        );

    \I__12065\ : InMux
    port map (
            O => \N__53905\,
            I => \N__53902\
        );

    \I__12064\ : LocalMux
    port map (
            O => \N__53902\,
            I => \N__53898\
        );

    \I__12063\ : InMux
    port map (
            O => \N__53901\,
            I => \N__53895\
        );

    \I__12062\ : Span4Mux_v
    port map (
            O => \N__53898\,
            I => \N__53892\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__53895\,
            I => \N__53889\
        );

    \I__12060\ : Span4Mux_h
    port map (
            O => \N__53892\,
            I => \N__53886\
        );

    \I__12059\ : Span4Mux_h
    port map (
            O => \N__53889\,
            I => \N__53883\
        );

    \I__12058\ : Span4Mux_v
    port map (
            O => \N__53886\,
            I => \N__53880\
        );

    \I__12057\ : Span4Mux_v
    port map (
            O => \N__53883\,
            I => \N__53877\
        );

    \I__12056\ : Span4Mux_v
    port map (
            O => \N__53880\,
            I => \N__53874\
        );

    \I__12055\ : Span4Mux_v
    port map (
            O => \N__53877\,
            I => \N__53871\
        );

    \I__12054\ : Odrv4
    port map (
            O => \N__53874\,
            I => \c0.n6404\
        );

    \I__12053\ : Odrv4
    port map (
            O => \N__53871\,
            I => \c0.n6404\
        );

    \I__12052\ : InMux
    port map (
            O => \N__53866\,
            I => \N__53863\
        );

    \I__12051\ : LocalMux
    port map (
            O => \N__53863\,
            I => \N__53859\
        );

    \I__12050\ : InMux
    port map (
            O => \N__53862\,
            I => \N__53856\
        );

    \I__12049\ : Span12Mux_v
    port map (
            O => \N__53859\,
            I => \N__53851\
        );

    \I__12048\ : LocalMux
    port map (
            O => \N__53856\,
            I => \N__53851\
        );

    \I__12047\ : Odrv12
    port map (
            O => \N__53851\,
            I => \c0.n21834\
        );

    \I__12046\ : InMux
    port map (
            O => \N__53848\,
            I => \N__53845\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__53845\,
            I => \N__53842\
        );

    \I__12044\ : Odrv4
    port map (
            O => \N__53842\,
            I => \c0.n22040\
        );

    \I__12043\ : CascadeMux
    port map (
            O => \N__53839\,
            I => \c0.n22040_cascade_\
        );

    \I__12042\ : InMux
    port map (
            O => \N__53836\,
            I => \N__53833\
        );

    \I__12041\ : LocalMux
    port map (
            O => \N__53833\,
            I => \N__53830\
        );

    \I__12040\ : Odrv4
    port map (
            O => \N__53830\,
            I => \c0.n21208\
        );

    \I__12039\ : InMux
    port map (
            O => \N__53827\,
            I => \N__53824\
        );

    \I__12038\ : LocalMux
    port map (
            O => \N__53824\,
            I => \c0.n21099\
        );

    \I__12037\ : CascadeMux
    port map (
            O => \N__53821\,
            I => \c0.n6_adj_4219_cascade_\
        );

    \I__12036\ : CascadeMux
    port map (
            O => \N__53818\,
            I => \N__53814\
        );

    \I__12035\ : InMux
    port map (
            O => \N__53817\,
            I => \N__53811\
        );

    \I__12034\ : InMux
    port map (
            O => \N__53814\,
            I => \N__53806\
        );

    \I__12033\ : LocalMux
    port map (
            O => \N__53811\,
            I => \N__53803\
        );

    \I__12032\ : InMux
    port map (
            O => \N__53810\,
            I => \N__53800\
        );

    \I__12031\ : InMux
    port map (
            O => \N__53809\,
            I => \N__53797\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__53806\,
            I => \c0.data_in_frame_21_2\
        );

    \I__12029\ : Odrv4
    port map (
            O => \N__53803\,
            I => \c0.data_in_frame_21_2\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__53800\,
            I => \c0.data_in_frame_21_2\
        );

    \I__12027\ : LocalMux
    port map (
            O => \N__53797\,
            I => \c0.data_in_frame_21_2\
        );

    \I__12026\ : InMux
    port map (
            O => \N__53788\,
            I => \N__53783\
        );

    \I__12025\ : InMux
    port map (
            O => \N__53787\,
            I => \N__53780\
        );

    \I__12024\ : InMux
    port map (
            O => \N__53786\,
            I => \N__53777\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__53783\,
            I => \c0.n22197\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__53780\,
            I => \c0.n22197\
        );

    \I__12021\ : LocalMux
    port map (
            O => \N__53777\,
            I => \c0.n22197\
        );

    \I__12020\ : CascadeMux
    port map (
            O => \N__53770\,
            I => \c0.n21949_cascade_\
        );

    \I__12019\ : InMux
    port map (
            O => \N__53767\,
            I => \N__53763\
        );

    \I__12018\ : CascadeMux
    port map (
            O => \N__53766\,
            I => \N__53759\
        );

    \I__12017\ : LocalMux
    port map (
            O => \N__53763\,
            I => \N__53756\
        );

    \I__12016\ : InMux
    port map (
            O => \N__53762\,
            I => \N__53751\
        );

    \I__12015\ : InMux
    port map (
            O => \N__53759\,
            I => \N__53751\
        );

    \I__12014\ : Odrv4
    port map (
            O => \N__53756\,
            I => \c0.n20137\
        );

    \I__12013\ : LocalMux
    port map (
            O => \N__53751\,
            I => \c0.n20137\
        );

    \I__12012\ : CascadeMux
    port map (
            O => \N__53746\,
            I => \c0.n22157_cascade_\
        );

    \I__12011\ : InMux
    port map (
            O => \N__53743\,
            I => \N__53740\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__53740\,
            I => \N__53737\
        );

    \I__12009\ : Span4Mux_h
    port map (
            O => \N__53737\,
            I => \N__53734\
        );

    \I__12008\ : Odrv4
    port map (
            O => \N__53734\,
            I => \c0.n20846\
        );

    \I__12007\ : CascadeMux
    port map (
            O => \N__53731\,
            I => \c0.n20846_cascade_\
        );

    \I__12006\ : InMux
    port map (
            O => \N__53728\,
            I => \N__53724\
        );

    \I__12005\ : CascadeMux
    port map (
            O => \N__53727\,
            I => \N__53721\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__53724\,
            I => \N__53716\
        );

    \I__12003\ : InMux
    port map (
            O => \N__53721\,
            I => \N__53713\
        );

    \I__12002\ : InMux
    port map (
            O => \N__53720\,
            I => \N__53710\
        );

    \I__12001\ : InMux
    port map (
            O => \N__53719\,
            I => \N__53707\
        );

    \I__12000\ : Sp12to4
    port map (
            O => \N__53716\,
            I => \N__53700\
        );

    \I__11999\ : LocalMux
    port map (
            O => \N__53713\,
            I => \N__53700\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__53710\,
            I => \N__53700\
        );

    \I__11997\ : LocalMux
    port map (
            O => \N__53707\,
            I => \c0.data_in_frame_25_4\
        );

    \I__11996\ : Odrv12
    port map (
            O => \N__53700\,
            I => \c0.data_in_frame_25_4\
        );

    \I__11995\ : InMux
    port map (
            O => \N__53695\,
            I => \N__53691\
        );

    \I__11994\ : CascadeMux
    port map (
            O => \N__53694\,
            I => \N__53686\
        );

    \I__11993\ : LocalMux
    port map (
            O => \N__53691\,
            I => \N__53683\
        );

    \I__11992\ : InMux
    port map (
            O => \N__53690\,
            I => \N__53678\
        );

    \I__11991\ : InMux
    port map (
            O => \N__53689\,
            I => \N__53678\
        );

    \I__11990\ : InMux
    port map (
            O => \N__53686\,
            I => \N__53675\
        );

    \I__11989\ : Span4Mux_h
    port map (
            O => \N__53683\,
            I => \N__53672\
        );

    \I__11988\ : LocalMux
    port map (
            O => \N__53678\,
            I => \N__53669\
        );

    \I__11987\ : LocalMux
    port map (
            O => \N__53675\,
            I => \N__53664\
        );

    \I__11986\ : Span4Mux_v
    port map (
            O => \N__53672\,
            I => \N__53664\
        );

    \I__11985\ : Span4Mux_h
    port map (
            O => \N__53669\,
            I => \N__53661\
        );

    \I__11984\ : Odrv4
    port map (
            O => \N__53664\,
            I => \c0.data_in_frame_25_2\
        );

    \I__11983\ : Odrv4
    port map (
            O => \N__53661\,
            I => \c0.data_in_frame_25_2\
        );

    \I__11982\ : InMux
    port map (
            O => \N__53656\,
            I => \N__53651\
        );

    \I__11981\ : CascadeMux
    port map (
            O => \N__53655\,
            I => \N__53647\
        );

    \I__11980\ : InMux
    port map (
            O => \N__53654\,
            I => \N__53644\
        );

    \I__11979\ : LocalMux
    port map (
            O => \N__53651\,
            I => \N__53641\
        );

    \I__11978\ : InMux
    port map (
            O => \N__53650\,
            I => \N__53636\
        );

    \I__11977\ : InMux
    port map (
            O => \N__53647\,
            I => \N__53636\
        );

    \I__11976\ : LocalMux
    port map (
            O => \N__53644\,
            I => \N__53633\
        );

    \I__11975\ : Span4Mux_v
    port map (
            O => \N__53641\,
            I => \N__53630\
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__53636\,
            I => \N__53627\
        );

    \I__11973\ : Span4Mux_h
    port map (
            O => \N__53633\,
            I => \N__53623\
        );

    \I__11972\ : Span4Mux_h
    port map (
            O => \N__53630\,
            I => \N__53618\
        );

    \I__11971\ : Span4Mux_h
    port map (
            O => \N__53627\,
            I => \N__53618\
        );

    \I__11970\ : InMux
    port map (
            O => \N__53626\,
            I => \N__53615\
        );

    \I__11969\ : Span4Mux_v
    port map (
            O => \N__53623\,
            I => \N__53612\
        );

    \I__11968\ : Span4Mux_v
    port map (
            O => \N__53618\,
            I => \N__53609\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__53615\,
            I => \c0.data_in_frame_25_3\
        );

    \I__11966\ : Odrv4
    port map (
            O => \N__53612\,
            I => \c0.data_in_frame_25_3\
        );

    \I__11965\ : Odrv4
    port map (
            O => \N__53609\,
            I => \c0.data_in_frame_25_3\
        );

    \I__11964\ : InMux
    port map (
            O => \N__53602\,
            I => \N__53595\
        );

    \I__11963\ : InMux
    port map (
            O => \N__53601\,
            I => \N__53590\
        );

    \I__11962\ : InMux
    port map (
            O => \N__53600\,
            I => \N__53590\
        );

    \I__11961\ : InMux
    port map (
            O => \N__53599\,
            I => \N__53587\
        );

    \I__11960\ : CascadeMux
    port map (
            O => \N__53598\,
            I => \N__53584\
        );

    \I__11959\ : LocalMux
    port map (
            O => \N__53595\,
            I => \N__53581\
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__53590\,
            I => \N__53576\
        );

    \I__11957\ : LocalMux
    port map (
            O => \N__53587\,
            I => \N__53576\
        );

    \I__11956\ : InMux
    port map (
            O => \N__53584\,
            I => \N__53573\
        );

    \I__11955\ : Span4Mux_h
    port map (
            O => \N__53581\,
            I => \N__53570\
        );

    \I__11954\ : Span4Mux_h
    port map (
            O => \N__53576\,
            I => \N__53567\
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__53573\,
            I => \c0.data_in_frame_25_5\
        );

    \I__11952\ : Odrv4
    port map (
            O => \N__53570\,
            I => \c0.data_in_frame_25_5\
        );

    \I__11951\ : Odrv4
    port map (
            O => \N__53567\,
            I => \c0.data_in_frame_25_5\
        );

    \I__11950\ : InMux
    port map (
            O => \N__53560\,
            I => \N__53557\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__53557\,
            I => \N__53554\
        );

    \I__11948\ : Span4Mux_h
    port map (
            O => \N__53554\,
            I => \N__53551\
        );

    \I__11947\ : Odrv4
    port map (
            O => \N__53551\,
            I => \c0.n22370\
        );

    \I__11946\ : InMux
    port map (
            O => \N__53548\,
            I => \N__53545\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__53545\,
            I => \c0.n12_adj_4491\
        );

    \I__11944\ : InMux
    port map (
            O => \N__53542\,
            I => \N__53539\
        );

    \I__11943\ : LocalMux
    port map (
            O => \N__53539\,
            I => \c0.n23009\
        );

    \I__11942\ : CascadeMux
    port map (
            O => \N__53536\,
            I => \c0.n22370_cascade_\
        );

    \I__11941\ : CascadeMux
    port map (
            O => \N__53533\,
            I => \N__53529\
        );

    \I__11940\ : InMux
    port map (
            O => \N__53532\,
            I => \N__53524\
        );

    \I__11939\ : InMux
    port map (
            O => \N__53529\,
            I => \N__53524\
        );

    \I__11938\ : LocalMux
    port map (
            O => \N__53524\,
            I => \N__53521\
        );

    \I__11937\ : Odrv4
    port map (
            O => \N__53521\,
            I => \c0.n23356\
        );

    \I__11936\ : SRMux
    port map (
            O => \N__53518\,
            I => \N__53515\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__53515\,
            I => \N__53512\
        );

    \I__11934\ : Span4Mux_h
    port map (
            O => \N__53512\,
            I => \N__53509\
        );

    \I__11933\ : Span4Mux_h
    port map (
            O => \N__53509\,
            I => \N__53506\
        );

    \I__11932\ : Odrv4
    port map (
            O => \N__53506\,
            I => \c0.n21366\
        );

    \I__11931\ : InMux
    port map (
            O => \N__53503\,
            I => \N__53499\
        );

    \I__11930\ : InMux
    port map (
            O => \N__53502\,
            I => \N__53496\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__53499\,
            I => \N__53493\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__53496\,
            I => \N__53490\
        );

    \I__11927\ : Span4Mux_h
    port map (
            O => \N__53493\,
            I => \N__53487\
        );

    \I__11926\ : Span4Mux_v
    port map (
            O => \N__53490\,
            I => \N__53482\
        );

    \I__11925\ : Span4Mux_v
    port map (
            O => \N__53487\,
            I => \N__53482\
        );

    \I__11924\ : Span4Mux_h
    port map (
            O => \N__53482\,
            I => \N__53479\
        );

    \I__11923\ : Odrv4
    port map (
            O => \N__53479\,
            I => \c0.n21855\
        );

    \I__11922\ : CascadeMux
    port map (
            O => \N__53476\,
            I => \N__53472\
        );

    \I__11921\ : InMux
    port map (
            O => \N__53475\,
            I => \N__53469\
        );

    \I__11920\ : InMux
    port map (
            O => \N__53472\,
            I => \N__53466\
        );

    \I__11919\ : LocalMux
    port map (
            O => \N__53469\,
            I => \N__53461\
        );

    \I__11918\ : LocalMux
    port map (
            O => \N__53466\,
            I => \N__53458\
        );

    \I__11917\ : InMux
    port map (
            O => \N__53465\,
            I => \N__53452\
        );

    \I__11916\ : InMux
    port map (
            O => \N__53464\,
            I => \N__53452\
        );

    \I__11915\ : Span4Mux_h
    port map (
            O => \N__53461\,
            I => \N__53449\
        );

    \I__11914\ : Span4Mux_h
    port map (
            O => \N__53458\,
            I => \N__53445\
        );

    \I__11913\ : InMux
    port map (
            O => \N__53457\,
            I => \N__53442\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__53452\,
            I => \N__53437\
        );

    \I__11911\ : Span4Mux_h
    port map (
            O => \N__53449\,
            I => \N__53437\
        );

    \I__11910\ : InMux
    port map (
            O => \N__53448\,
            I => \N__53433\
        );

    \I__11909\ : Span4Mux_v
    port map (
            O => \N__53445\,
            I => \N__53426\
        );

    \I__11908\ : LocalMux
    port map (
            O => \N__53442\,
            I => \N__53426\
        );

    \I__11907\ : Span4Mux_v
    port map (
            O => \N__53437\,
            I => \N__53426\
        );

    \I__11906\ : InMux
    port map (
            O => \N__53436\,
            I => \N__53423\
        );

    \I__11905\ : LocalMux
    port map (
            O => \N__53433\,
            I => encoder0_position_2
        );

    \I__11904\ : Odrv4
    port map (
            O => \N__53426\,
            I => encoder0_position_2
        );

    \I__11903\ : LocalMux
    port map (
            O => \N__53423\,
            I => encoder0_position_2
        );

    \I__11902\ : InMux
    port map (
            O => \N__53416\,
            I => \N__53413\
        );

    \I__11901\ : LocalMux
    port map (
            O => \N__53413\,
            I => \N__53410\
        );

    \I__11900\ : Span4Mux_h
    port map (
            O => \N__53410\,
            I => \N__53406\
        );

    \I__11899\ : InMux
    port map (
            O => \N__53409\,
            I => \N__53403\
        );

    \I__11898\ : Span4Mux_h
    port map (
            O => \N__53406\,
            I => \N__53400\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__53403\,
            I => \N__53397\
        );

    \I__11896\ : Odrv4
    port map (
            O => \N__53400\,
            I => \c0.n22248\
        );

    \I__11895\ : Odrv4
    port map (
            O => \N__53397\,
            I => \c0.n22248\
        );

    \I__11894\ : InMux
    port map (
            O => \N__53392\,
            I => \N__53389\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__53389\,
            I => \N__53383\
        );

    \I__11892\ : InMux
    port map (
            O => \N__53388\,
            I => \N__53380\
        );

    \I__11891\ : InMux
    port map (
            O => \N__53387\,
            I => \N__53375\
        );

    \I__11890\ : InMux
    port map (
            O => \N__53386\,
            I => \N__53375\
        );

    \I__11889\ : Span4Mux_h
    port map (
            O => \N__53383\,
            I => \N__53372\
        );

    \I__11888\ : LocalMux
    port map (
            O => \N__53380\,
            I => \N__53369\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__53375\,
            I => \N__53365\
        );

    \I__11886\ : Span4Mux_v
    port map (
            O => \N__53372\,
            I => \N__53360\
        );

    \I__11885\ : Span4Mux_h
    port map (
            O => \N__53369\,
            I => \N__53360\
        );

    \I__11884\ : InMux
    port map (
            O => \N__53368\,
            I => \N__53357\
        );

    \I__11883\ : Span4Mux_h
    port map (
            O => \N__53365\,
            I => \N__53354\
        );

    \I__11882\ : Span4Mux_h
    port map (
            O => \N__53360\,
            I => \N__53351\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__53357\,
            I => \N__53346\
        );

    \I__11880\ : Sp12to4
    port map (
            O => \N__53354\,
            I => \N__53346\
        );

    \I__11879\ : Span4Mux_v
    port map (
            O => \N__53351\,
            I => \N__53343\
        );

    \I__11878\ : Span12Mux_v
    port map (
            O => \N__53346\,
            I => \N__53340\
        );

    \I__11877\ : Odrv4
    port map (
            O => \N__53343\,
            I => \c0.n13379\
        );

    \I__11876\ : Odrv12
    port map (
            O => \N__53340\,
            I => \c0.n13379\
        );

    \I__11875\ : CascadeMux
    port map (
            O => \N__53335\,
            I => \N__53332\
        );

    \I__11874\ : InMux
    port map (
            O => \N__53332\,
            I => \N__53329\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__53329\,
            I => \N__53325\
        );

    \I__11872\ : InMux
    port map (
            O => \N__53328\,
            I => \N__53322\
        );

    \I__11871\ : Span4Mux_v
    port map (
            O => \N__53325\,
            I => \N__53318\
        );

    \I__11870\ : LocalMux
    port map (
            O => \N__53322\,
            I => \N__53315\
        );

    \I__11869\ : InMux
    port map (
            O => \N__53321\,
            I => \N__53312\
        );

    \I__11868\ : Span4Mux_h
    port map (
            O => \N__53318\,
            I => \N__53307\
        );

    \I__11867\ : Span4Mux_v
    port map (
            O => \N__53315\,
            I => \N__53307\
        );

    \I__11866\ : LocalMux
    port map (
            O => \N__53312\,
            I => \c0.data_in_frame_20_7\
        );

    \I__11865\ : Odrv4
    port map (
            O => \N__53307\,
            I => \c0.data_in_frame_20_7\
        );

    \I__11864\ : CascadeMux
    port map (
            O => \N__53302\,
            I => \c0.n28_cascade_\
        );

    \I__11863\ : CascadeMux
    port map (
            O => \N__53299\,
            I => \c0.n23640_cascade_\
        );

    \I__11862\ : CascadeMux
    port map (
            O => \N__53296\,
            I => \c0.n22305_cascade_\
        );

    \I__11861\ : InMux
    port map (
            O => \N__53293\,
            I => \N__53287\
        );

    \I__11860\ : InMux
    port map (
            O => \N__53292\,
            I => \N__53287\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__53287\,
            I => \N__53283\
        );

    \I__11858\ : InMux
    port map (
            O => \N__53286\,
            I => \N__53280\
        );

    \I__11857\ : Span4Mux_v
    port map (
            O => \N__53283\,
            I => \N__53274\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__53280\,
            I => \N__53274\
        );

    \I__11855\ : CascadeMux
    port map (
            O => \N__53279\,
            I => \N__53271\
        );

    \I__11854\ : Span4Mux_h
    port map (
            O => \N__53274\,
            I => \N__53268\
        );

    \I__11853\ : InMux
    port map (
            O => \N__53271\,
            I => \N__53265\
        );

    \I__11852\ : Span4Mux_h
    port map (
            O => \N__53268\,
            I => \N__53262\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__53265\,
            I => \c0.data_in_frame_21_1\
        );

    \I__11850\ : Odrv4
    port map (
            O => \N__53262\,
            I => \c0.data_in_frame_21_1\
        );

    \I__11849\ : InMux
    port map (
            O => \N__53257\,
            I => \N__53251\
        );

    \I__11848\ : InMux
    port map (
            O => \N__53256\,
            I => \N__53251\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__53251\,
            I => \c0.n23640\
        );

    \I__11846\ : InMux
    port map (
            O => \N__53248\,
            I => \N__53245\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__53245\,
            I => \c0.n22305\
        );

    \I__11844\ : InMux
    port map (
            O => \N__53242\,
            I => \N__53238\
        );

    \I__11843\ : InMux
    port map (
            O => \N__53241\,
            I => \N__53235\
        );

    \I__11842\ : LocalMux
    port map (
            O => \N__53238\,
            I => \N__53232\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__53235\,
            I => \c0.data_in_frame_20_1\
        );

    \I__11840\ : Odrv4
    port map (
            O => \N__53232\,
            I => \c0.data_in_frame_20_1\
        );

    \I__11839\ : CascadeMux
    port map (
            O => \N__53227\,
            I => \c0.n6_adj_4226_cascade_\
        );

    \I__11838\ : CascadeMux
    port map (
            O => \N__53224\,
            I => \c0.n23615_cascade_\
        );

    \I__11837\ : CascadeMux
    port map (
            O => \N__53221\,
            I => \c0.n22100_cascade_\
        );

    \I__11836\ : InMux
    port map (
            O => \N__53218\,
            I => \N__53214\
        );

    \I__11835\ : InMux
    port map (
            O => \N__53217\,
            I => \N__53211\
        );

    \I__11834\ : LocalMux
    port map (
            O => \N__53214\,
            I => \c0.n22081\
        );

    \I__11833\ : LocalMux
    port map (
            O => \N__53211\,
            I => \c0.n22081\
        );

    \I__11832\ : CascadeMux
    port map (
            O => \N__53206\,
            I => \N__53203\
        );

    \I__11831\ : InMux
    port map (
            O => \N__53203\,
            I => \N__53200\
        );

    \I__11830\ : LocalMux
    port map (
            O => \N__53200\,
            I => \c0.n6_adj_4224\
        );

    \I__11829\ : InMux
    port map (
            O => \N__53197\,
            I => \N__53190\
        );

    \I__11828\ : InMux
    port map (
            O => \N__53196\,
            I => \N__53185\
        );

    \I__11827\ : InMux
    port map (
            O => \N__53195\,
            I => \N__53182\
        );

    \I__11826\ : InMux
    port map (
            O => \N__53194\,
            I => \N__53178\
        );

    \I__11825\ : InMux
    port map (
            O => \N__53193\,
            I => \N__53171\
        );

    \I__11824\ : LocalMux
    port map (
            O => \N__53190\,
            I => \N__53165\
        );

    \I__11823\ : InMux
    port map (
            O => \N__53189\,
            I => \N__53162\
        );

    \I__11822\ : InMux
    port map (
            O => \N__53188\,
            I => \N__53159\
        );

    \I__11821\ : LocalMux
    port map (
            O => \N__53185\,
            I => \N__53156\
        );

    \I__11820\ : LocalMux
    port map (
            O => \N__53182\,
            I => \N__53153\
        );

    \I__11819\ : InMux
    port map (
            O => \N__53181\,
            I => \N__53150\
        );

    \I__11818\ : LocalMux
    port map (
            O => \N__53178\,
            I => \N__53147\
        );

    \I__11817\ : InMux
    port map (
            O => \N__53177\,
            I => \N__53144\
        );

    \I__11816\ : InMux
    port map (
            O => \N__53176\,
            I => \N__53141\
        );

    \I__11815\ : InMux
    port map (
            O => \N__53175\,
            I => \N__53138\
        );

    \I__11814\ : CascadeMux
    port map (
            O => \N__53174\,
            I => \N__53132\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__53171\,
            I => \N__53125\
        );

    \I__11812\ : InMux
    port map (
            O => \N__53170\,
            I => \N__53120\
        );

    \I__11811\ : InMux
    port map (
            O => \N__53169\,
            I => \N__53120\
        );

    \I__11810\ : CascadeMux
    port map (
            O => \N__53168\,
            I => \N__53117\
        );

    \I__11809\ : Span4Mux_v
    port map (
            O => \N__53165\,
            I => \N__53110\
        );

    \I__11808\ : LocalMux
    port map (
            O => \N__53162\,
            I => \N__53110\
        );

    \I__11807\ : LocalMux
    port map (
            O => \N__53159\,
            I => \N__53105\
        );

    \I__11806\ : Span4Mux_v
    port map (
            O => \N__53156\,
            I => \N__53105\
        );

    \I__11805\ : Span4Mux_v
    port map (
            O => \N__53153\,
            I => \N__53098\
        );

    \I__11804\ : LocalMux
    port map (
            O => \N__53150\,
            I => \N__53098\
        );

    \I__11803\ : Span4Mux_v
    port map (
            O => \N__53147\,
            I => \N__53098\
        );

    \I__11802\ : LocalMux
    port map (
            O => \N__53144\,
            I => \N__53093\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__53141\,
            I => \N__53093\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__53138\,
            I => \N__53090\
        );

    \I__11799\ : InMux
    port map (
            O => \N__53137\,
            I => \N__53087\
        );

    \I__11798\ : InMux
    port map (
            O => \N__53136\,
            I => \N__53084\
        );

    \I__11797\ : InMux
    port map (
            O => \N__53135\,
            I => \N__53077\
        );

    \I__11796\ : InMux
    port map (
            O => \N__53132\,
            I => \N__53077\
        );

    \I__11795\ : InMux
    port map (
            O => \N__53131\,
            I => \N__53077\
        );

    \I__11794\ : InMux
    port map (
            O => \N__53130\,
            I => \N__53070\
        );

    \I__11793\ : InMux
    port map (
            O => \N__53129\,
            I => \N__53070\
        );

    \I__11792\ : InMux
    port map (
            O => \N__53128\,
            I => \N__53070\
        );

    \I__11791\ : Span4Mux_v
    port map (
            O => \N__53125\,
            I => \N__53065\
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__53120\,
            I => \N__53065\
        );

    \I__11789\ : InMux
    port map (
            O => \N__53117\,
            I => \N__53058\
        );

    \I__11788\ : InMux
    port map (
            O => \N__53116\,
            I => \N__53058\
        );

    \I__11787\ : InMux
    port map (
            O => \N__53115\,
            I => \N__53058\
        );

    \I__11786\ : Span4Mux_h
    port map (
            O => \N__53110\,
            I => \N__53053\
        );

    \I__11785\ : Span4Mux_h
    port map (
            O => \N__53105\,
            I => \N__53053\
        );

    \I__11784\ : Span4Mux_h
    port map (
            O => \N__53098\,
            I => \N__53046\
        );

    \I__11783\ : Span4Mux_v
    port map (
            O => \N__53093\,
            I => \N__53046\
        );

    \I__11782\ : Span4Mux_h
    port map (
            O => \N__53090\,
            I => \N__53046\
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__53087\,
            I => \c0.n21737\
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__53084\,
            I => \c0.n21737\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__53077\,
            I => \c0.n21737\
        );

    \I__11778\ : LocalMux
    port map (
            O => \N__53070\,
            I => \c0.n21737\
        );

    \I__11777\ : Odrv4
    port map (
            O => \N__53065\,
            I => \c0.n21737\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__53058\,
            I => \c0.n21737\
        );

    \I__11775\ : Odrv4
    port map (
            O => \N__53053\,
            I => \c0.n21737\
        );

    \I__11774\ : Odrv4
    port map (
            O => \N__53046\,
            I => \c0.n21737\
        );

    \I__11773\ : InMux
    port map (
            O => \N__53029\,
            I => \N__53023\
        );

    \I__11772\ : InMux
    port map (
            O => \N__53028\,
            I => \N__53016\
        );

    \I__11771\ : InMux
    port map (
            O => \N__53027\,
            I => \N__53013\
        );

    \I__11770\ : InMux
    port map (
            O => \N__53026\,
            I => \N__53006\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__53023\,
            I => \N__53003\
        );

    \I__11768\ : InMux
    port map (
            O => \N__53022\,
            I => \N__53000\
        );

    \I__11767\ : InMux
    port map (
            O => \N__53021\,
            I => \N__52993\
        );

    \I__11766\ : InMux
    port map (
            O => \N__53020\,
            I => \N__52993\
        );

    \I__11765\ : InMux
    port map (
            O => \N__53019\,
            I => \N__52993\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__53016\,
            I => \N__52988\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__53013\,
            I => \N__52988\
        );

    \I__11762\ : InMux
    port map (
            O => \N__53012\,
            I => \N__52985\
        );

    \I__11761\ : InMux
    port map (
            O => \N__53011\,
            I => \N__52982\
        );

    \I__11760\ : InMux
    port map (
            O => \N__53010\,
            I => \N__52978\
        );

    \I__11759\ : InMux
    port map (
            O => \N__53009\,
            I => \N__52975\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__53006\,
            I => \N__52967\
        );

    \I__11757\ : Span4Mux_h
    port map (
            O => \N__53003\,
            I => \N__52964\
        );

    \I__11756\ : LocalMux
    port map (
            O => \N__53000\,
            I => \N__52961\
        );

    \I__11755\ : LocalMux
    port map (
            O => \N__52993\,
            I => \N__52958\
        );

    \I__11754\ : Span4Mux_v
    port map (
            O => \N__52988\,
            I => \N__52951\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__52985\,
            I => \N__52951\
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__52982\,
            I => \N__52951\
        );

    \I__11751\ : InMux
    port map (
            O => \N__52981\,
            I => \N__52948\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__52978\,
            I => \N__52942\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__52975\,
            I => \N__52942\
        );

    \I__11748\ : InMux
    port map (
            O => \N__52974\,
            I => \N__52939\
        );

    \I__11747\ : InMux
    port map (
            O => \N__52973\,
            I => \N__52934\
        );

    \I__11746\ : InMux
    port map (
            O => \N__52972\,
            I => \N__52934\
        );

    \I__11745\ : InMux
    port map (
            O => \N__52971\,
            I => \N__52929\
        );

    \I__11744\ : InMux
    port map (
            O => \N__52970\,
            I => \N__52929\
        );

    \I__11743\ : Span4Mux_h
    port map (
            O => \N__52967\,
            I => \N__52924\
        );

    \I__11742\ : Span4Mux_h
    port map (
            O => \N__52964\,
            I => \N__52924\
        );

    \I__11741\ : Span4Mux_v
    port map (
            O => \N__52961\,
            I => \N__52919\
        );

    \I__11740\ : Span4Mux_h
    port map (
            O => \N__52958\,
            I => \N__52919\
        );

    \I__11739\ : Span4Mux_v
    port map (
            O => \N__52951\,
            I => \N__52914\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__52948\,
            I => \N__52914\
        );

    \I__11737\ : InMux
    port map (
            O => \N__52947\,
            I => \N__52911\
        );

    \I__11736\ : Span4Mux_v
    port map (
            O => \N__52942\,
            I => \N__52902\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__52939\,
            I => \N__52902\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__52934\,
            I => \N__52902\
        );

    \I__11733\ : LocalMux
    port map (
            O => \N__52929\,
            I => \N__52902\
        );

    \I__11732\ : Odrv4
    port map (
            O => \N__52924\,
            I => \c0.n6_adj_4353\
        );

    \I__11731\ : Odrv4
    port map (
            O => \N__52919\,
            I => \c0.n6_adj_4353\
        );

    \I__11730\ : Odrv4
    port map (
            O => \N__52914\,
            I => \c0.n6_adj_4353\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__52911\,
            I => \c0.n6_adj_4353\
        );

    \I__11728\ : Odrv4
    port map (
            O => \N__52902\,
            I => \c0.n6_adj_4353\
        );

    \I__11727\ : InMux
    port map (
            O => \N__52891\,
            I => \N__52881\
        );

    \I__11726\ : InMux
    port map (
            O => \N__52890\,
            I => \N__52878\
        );

    \I__11725\ : InMux
    port map (
            O => \N__52889\,
            I => \N__52875\
        );

    \I__11724\ : InMux
    port map (
            O => \N__52888\,
            I => \N__52864\
        );

    \I__11723\ : InMux
    port map (
            O => \N__52887\,
            I => \N__52861\
        );

    \I__11722\ : InMux
    port map (
            O => \N__52886\,
            I => \N__52855\
        );

    \I__11721\ : InMux
    port map (
            O => \N__52885\,
            I => \N__52852\
        );

    \I__11720\ : InMux
    port map (
            O => \N__52884\,
            I => \N__52849\
        );

    \I__11719\ : LocalMux
    port map (
            O => \N__52881\,
            I => \N__52840\
        );

    \I__11718\ : LocalMux
    port map (
            O => \N__52878\,
            I => \N__52837\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__52875\,
            I => \N__52834\
        );

    \I__11716\ : InMux
    port map (
            O => \N__52874\,
            I => \N__52831\
        );

    \I__11715\ : InMux
    port map (
            O => \N__52873\,
            I => \N__52828\
        );

    \I__11714\ : InMux
    port map (
            O => \N__52872\,
            I => \N__52825\
        );

    \I__11713\ : InMux
    port map (
            O => \N__52871\,
            I => \N__52822\
        );

    \I__11712\ : InMux
    port map (
            O => \N__52870\,
            I => \N__52819\
        );

    \I__11711\ : InMux
    port map (
            O => \N__52869\,
            I => \N__52816\
        );

    \I__11710\ : InMux
    port map (
            O => \N__52868\,
            I => \N__52812\
        );

    \I__11709\ : InMux
    port map (
            O => \N__52867\,
            I => \N__52809\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__52864\,
            I => \N__52804\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__52861\,
            I => \N__52804\
        );

    \I__11706\ : InMux
    port map (
            O => \N__52860\,
            I => \N__52801\
        );

    \I__11705\ : InMux
    port map (
            O => \N__52859\,
            I => \N__52798\
        );

    \I__11704\ : InMux
    port map (
            O => \N__52858\,
            I => \N__52795\
        );

    \I__11703\ : LocalMux
    port map (
            O => \N__52855\,
            I => \N__52792\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__52852\,
            I => \N__52787\
        );

    \I__11701\ : LocalMux
    port map (
            O => \N__52849\,
            I => \N__52787\
        );

    \I__11700\ : InMux
    port map (
            O => \N__52848\,
            I => \N__52784\
        );

    \I__11699\ : InMux
    port map (
            O => \N__52847\,
            I => \N__52781\
        );

    \I__11698\ : InMux
    port map (
            O => \N__52846\,
            I => \N__52778\
        );

    \I__11697\ : InMux
    port map (
            O => \N__52845\,
            I => \N__52775\
        );

    \I__11696\ : InMux
    port map (
            O => \N__52844\,
            I => \N__52772\
        );

    \I__11695\ : InMux
    port map (
            O => \N__52843\,
            I => \N__52769\
        );

    \I__11694\ : Span4Mux_h
    port map (
            O => \N__52840\,
            I => \N__52764\
        );

    \I__11693\ : Span4Mux_v
    port map (
            O => \N__52837\,
            I => \N__52764\
        );

    \I__11692\ : Span4Mux_v
    port map (
            O => \N__52834\,
            I => \N__52749\
        );

    \I__11691\ : LocalMux
    port map (
            O => \N__52831\,
            I => \N__52749\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__52828\,
            I => \N__52749\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__52825\,
            I => \N__52749\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__52822\,
            I => \N__52749\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__52819\,
            I => \N__52749\
        );

    \I__11686\ : LocalMux
    port map (
            O => \N__52816\,
            I => \N__52749\
        );

    \I__11685\ : InMux
    port map (
            O => \N__52815\,
            I => \N__52746\
        );

    \I__11684\ : LocalMux
    port map (
            O => \N__52812\,
            I => \N__52741\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__52809\,
            I => \N__52738\
        );

    \I__11682\ : Span4Mux_v
    port map (
            O => \N__52804\,
            I => \N__52731\
        );

    \I__11681\ : LocalMux
    port map (
            O => \N__52801\,
            I => \N__52731\
        );

    \I__11680\ : LocalMux
    port map (
            O => \N__52798\,
            I => \N__52731\
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__52795\,
            I => \N__52728\
        );

    \I__11678\ : Span4Mux_v
    port map (
            O => \N__52792\,
            I => \N__52725\
        );

    \I__11677\ : Span4Mux_h
    port map (
            O => \N__52787\,
            I => \N__52710\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__52784\,
            I => \N__52710\
        );

    \I__11675\ : LocalMux
    port map (
            O => \N__52781\,
            I => \N__52710\
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__52778\,
            I => \N__52710\
        );

    \I__11673\ : LocalMux
    port map (
            O => \N__52775\,
            I => \N__52710\
        );

    \I__11672\ : LocalMux
    port map (
            O => \N__52772\,
            I => \N__52710\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__52769\,
            I => \N__52710\
        );

    \I__11670\ : Span4Mux_h
    port map (
            O => \N__52764\,
            I => \N__52703\
        );

    \I__11669\ : Span4Mux_v
    port map (
            O => \N__52749\,
            I => \N__52703\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__52746\,
            I => \N__52703\
        );

    \I__11667\ : InMux
    port map (
            O => \N__52745\,
            I => \N__52700\
        );

    \I__11666\ : InMux
    port map (
            O => \N__52744\,
            I => \N__52697\
        );

    \I__11665\ : Span12Mux_h
    port map (
            O => \N__52741\,
            I => \N__52694\
        );

    \I__11664\ : Span4Mux_h
    port map (
            O => \N__52738\,
            I => \N__52691\
        );

    \I__11663\ : Span4Mux_v
    port map (
            O => \N__52731\,
            I => \N__52686\
        );

    \I__11662\ : Span4Mux_h
    port map (
            O => \N__52728\,
            I => \N__52686\
        );

    \I__11661\ : Span4Mux_v
    port map (
            O => \N__52725\,
            I => \N__52679\
        );

    \I__11660\ : Span4Mux_v
    port map (
            O => \N__52710\,
            I => \N__52679\
        );

    \I__11659\ : Span4Mux_h
    port map (
            O => \N__52703\,
            I => \N__52679\
        );

    \I__11658\ : LocalMux
    port map (
            O => \N__52700\,
            I => \N__52674\
        );

    \I__11657\ : LocalMux
    port map (
            O => \N__52697\,
            I => \N__52674\
        );

    \I__11656\ : Odrv12
    port map (
            O => \N__52694\,
            I => \c0.n5_adj_4342\
        );

    \I__11655\ : Odrv4
    port map (
            O => \N__52691\,
            I => \c0.n5_adj_4342\
        );

    \I__11654\ : Odrv4
    port map (
            O => \N__52686\,
            I => \c0.n5_adj_4342\
        );

    \I__11653\ : Odrv4
    port map (
            O => \N__52679\,
            I => \c0.n5_adj_4342\
        );

    \I__11652\ : Odrv12
    port map (
            O => \N__52674\,
            I => \c0.n5_adj_4342\
        );

    \I__11651\ : CascadeMux
    port map (
            O => \N__52663\,
            I => \N__52660\
        );

    \I__11650\ : InMux
    port map (
            O => \N__52660\,
            I => \N__52654\
        );

    \I__11649\ : InMux
    port map (
            O => \N__52659\,
            I => \N__52654\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__52654\,
            I => \N__52651\
        );

    \I__11647\ : Span4Mux_h
    port map (
            O => \N__52651\,
            I => \N__52646\
        );

    \I__11646\ : InMux
    port map (
            O => \N__52650\,
            I => \N__52641\
        );

    \I__11645\ : InMux
    port map (
            O => \N__52649\,
            I => \N__52641\
        );

    \I__11644\ : Span4Mux_v
    port map (
            O => \N__52646\,
            I => \N__52638\
        );

    \I__11643\ : LocalMux
    port map (
            O => \N__52641\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__11642\ : Odrv4
    port map (
            O => \N__52638\,
            I => \c0.FRAME_MATCHER_state_20\
        );

    \I__11641\ : InMux
    port map (
            O => \N__52633\,
            I => \N__52630\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__52630\,
            I => \N__52626\
        );

    \I__11639\ : InMux
    port map (
            O => \N__52629\,
            I => \N__52623\
        );

    \I__11638\ : Span4Mux_v
    port map (
            O => \N__52626\,
            I => \N__52618\
        );

    \I__11637\ : LocalMux
    port map (
            O => \N__52623\,
            I => \N__52618\
        );

    \I__11636\ : Span4Mux_h
    port map (
            O => \N__52618\,
            I => \N__52615\
        );

    \I__11635\ : Odrv4
    port map (
            O => \N__52615\,
            I => \c0.n13190\
        );

    \I__11634\ : CascadeMux
    port map (
            O => \N__52612\,
            I => \c0.n18_adj_4222_cascade_\
        );

    \I__11633\ : InMux
    port map (
            O => \N__52609\,
            I => \N__52605\
        );

    \I__11632\ : InMux
    port map (
            O => \N__52608\,
            I => \N__52602\
        );

    \I__11631\ : LocalMux
    port map (
            O => \N__52605\,
            I => \N__52597\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__52602\,
            I => \N__52597\
        );

    \I__11629\ : Span4Mux_v
    port map (
            O => \N__52597\,
            I => \N__52593\
        );

    \I__11628\ : InMux
    port map (
            O => \N__52596\,
            I => \N__52590\
        );

    \I__11627\ : Odrv4
    port map (
            O => \N__52593\,
            I => \c0.n22270\
        );

    \I__11626\ : LocalMux
    port map (
            O => \N__52590\,
            I => \c0.n22270\
        );

    \I__11625\ : InMux
    port map (
            O => \N__52585\,
            I => \N__52582\
        );

    \I__11624\ : LocalMux
    port map (
            O => \N__52582\,
            I => \N__52579\
        );

    \I__11623\ : Odrv12
    port map (
            O => \N__52579\,
            I => \c0.n6_adj_4221\
        );

    \I__11622\ : InMux
    port map (
            O => \N__52576\,
            I => \N__52573\
        );

    \I__11621\ : LocalMux
    port map (
            O => \N__52573\,
            I => \N__52570\
        );

    \I__11620\ : Span4Mux_h
    port map (
            O => \N__52570\,
            I => \N__52567\
        );

    \I__11619\ : Odrv4
    port map (
            O => \N__52567\,
            I => \c0.n22308\
        );

    \I__11618\ : CascadeMux
    port map (
            O => \N__52564\,
            I => \c0.n22003_cascade_\
        );

    \I__11617\ : InMux
    port map (
            O => \N__52561\,
            I => \N__52558\
        );

    \I__11616\ : LocalMux
    port map (
            O => \N__52558\,
            I => \c0.n5943\
        );

    \I__11615\ : CascadeMux
    port map (
            O => \N__52555\,
            I => \c0.n6221_cascade_\
        );

    \I__11614\ : InMux
    port map (
            O => \N__52552\,
            I => \N__52549\
        );

    \I__11613\ : LocalMux
    port map (
            O => \N__52549\,
            I => \c0.n22003\
        );

    \I__11612\ : InMux
    port map (
            O => \N__52546\,
            I => \N__52543\
        );

    \I__11611\ : LocalMux
    port map (
            O => \N__52543\,
            I => \N__52540\
        );

    \I__11610\ : Span4Mux_h
    port map (
            O => \N__52540\,
            I => \N__52536\
        );

    \I__11609\ : InMux
    port map (
            O => \N__52539\,
            I => \N__52531\
        );

    \I__11608\ : Span4Mux_v
    port map (
            O => \N__52536\,
            I => \N__52528\
        );

    \I__11607\ : InMux
    port map (
            O => \N__52535\,
            I => \N__52525\
        );

    \I__11606\ : InMux
    port map (
            O => \N__52534\,
            I => \N__52522\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__52531\,
            I => \c0.data_in_frame_10_2\
        );

    \I__11604\ : Odrv4
    port map (
            O => \N__52528\,
            I => \c0.data_in_frame_10_2\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__52525\,
            I => \c0.data_in_frame_10_2\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__52522\,
            I => \c0.data_in_frame_10_2\
        );

    \I__11601\ : CascadeMux
    port map (
            O => \N__52513\,
            I => \c0.n20402_cascade_\
        );

    \I__11600\ : InMux
    port map (
            O => \N__52510\,
            I => \N__52506\
        );

    \I__11599\ : CascadeMux
    port map (
            O => \N__52509\,
            I => \N__52502\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__52506\,
            I => \N__52499\
        );

    \I__11597\ : InMux
    port map (
            O => \N__52505\,
            I => \N__52496\
        );

    \I__11596\ : InMux
    port map (
            O => \N__52502\,
            I => \N__52493\
        );

    \I__11595\ : Span4Mux_v
    port map (
            O => \N__52499\,
            I => \N__52490\
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__52496\,
            I => \N__52487\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__52493\,
            I => \c0.data_in_frame_9_6\
        );

    \I__11592\ : Odrv4
    port map (
            O => \N__52490\,
            I => \c0.data_in_frame_9_6\
        );

    \I__11591\ : Odrv4
    port map (
            O => \N__52487\,
            I => \c0.data_in_frame_9_6\
        );

    \I__11590\ : CascadeMux
    port map (
            O => \N__52480\,
            I => \N__52477\
        );

    \I__11589\ : InMux
    port map (
            O => \N__52477\,
            I => \N__52470\
        );

    \I__11588\ : InMux
    port map (
            O => \N__52476\,
            I => \N__52470\
        );

    \I__11587\ : InMux
    port map (
            O => \N__52475\,
            I => \N__52467\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__52470\,
            I => \c0.data_in_frame_9_4\
        );

    \I__11585\ : LocalMux
    port map (
            O => \N__52467\,
            I => \c0.data_in_frame_9_4\
        );

    \I__11584\ : InMux
    port map (
            O => \N__52462\,
            I => \N__52456\
        );

    \I__11583\ : InMux
    port map (
            O => \N__52461\,
            I => \N__52456\
        );

    \I__11582\ : LocalMux
    port map (
            O => \N__52456\,
            I => \N__52453\
        );

    \I__11581\ : Odrv4
    port map (
            O => \N__52453\,
            I => \c0.n21873\
        );

    \I__11580\ : InMux
    port map (
            O => \N__52450\,
            I => \N__52447\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__52447\,
            I => \N__52444\
        );

    \I__11578\ : Span4Mux_v
    port map (
            O => \N__52444\,
            I => \N__52440\
        );

    \I__11577\ : InMux
    port map (
            O => \N__52443\,
            I => \N__52437\
        );

    \I__11576\ : Span4Mux_h
    port map (
            O => \N__52440\,
            I => \N__52432\
        );

    \I__11575\ : LocalMux
    port map (
            O => \N__52437\,
            I => \N__52432\
        );

    \I__11574\ : Span4Mux_h
    port map (
            O => \N__52432\,
            I => \N__52429\
        );

    \I__11573\ : Odrv4
    port map (
            O => \N__52429\,
            I => \c0.n13287\
        );

    \I__11572\ : InMux
    port map (
            O => \N__52426\,
            I => \N__52423\
        );

    \I__11571\ : LocalMux
    port map (
            O => \N__52423\,
            I => \N__52420\
        );

    \I__11570\ : Span4Mux_h
    port map (
            O => \N__52420\,
            I => \N__52417\
        );

    \I__11569\ : Span4Mux_v
    port map (
            O => \N__52417\,
            I => \N__52414\
        );

    \I__11568\ : Odrv4
    port map (
            O => \N__52414\,
            I => \c0.n22443\
        );

    \I__11567\ : CascadeMux
    port map (
            O => \N__52411\,
            I => \c0.n10_adj_4242_cascade_\
        );

    \I__11566\ : InMux
    port map (
            O => \N__52408\,
            I => \N__52404\
        );

    \I__11565\ : CascadeMux
    port map (
            O => \N__52407\,
            I => \N__52401\
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__52404\,
            I => \N__52398\
        );

    \I__11563\ : InMux
    port map (
            O => \N__52401\,
            I => \N__52395\
        );

    \I__11562\ : Span4Mux_h
    port map (
            O => \N__52398\,
            I => \N__52392\
        );

    \I__11561\ : LocalMux
    port map (
            O => \N__52395\,
            I => \N__52386\
        );

    \I__11560\ : Span4Mux_h
    port map (
            O => \N__52392\,
            I => \N__52386\
        );

    \I__11559\ : InMux
    port map (
            O => \N__52391\,
            I => \N__52383\
        );

    \I__11558\ : Odrv4
    port map (
            O => \N__52386\,
            I => \c0.data_in_frame_8_1\
        );

    \I__11557\ : LocalMux
    port map (
            O => \N__52383\,
            I => \c0.data_in_frame_8_1\
        );

    \I__11556\ : InMux
    port map (
            O => \N__52378\,
            I => \N__52372\
        );

    \I__11555\ : InMux
    port map (
            O => \N__52377\,
            I => \N__52367\
        );

    \I__11554\ : InMux
    port map (
            O => \N__52376\,
            I => \N__52367\
        );

    \I__11553\ : InMux
    port map (
            O => \N__52375\,
            I => \N__52364\
        );

    \I__11552\ : LocalMux
    port map (
            O => \N__52372\,
            I => \N__52361\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__52367\,
            I => \N__52358\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__52364\,
            I => \c0.data_in_frame_16_6\
        );

    \I__11549\ : Odrv4
    port map (
            O => \N__52361\,
            I => \c0.data_in_frame_16_6\
        );

    \I__11548\ : Odrv4
    port map (
            O => \N__52358\,
            I => \c0.data_in_frame_16_6\
        );

    \I__11547\ : CascadeMux
    port map (
            O => \N__52351\,
            I => \c0.n13786_cascade_\
        );

    \I__11546\ : InMux
    port map (
            O => \N__52348\,
            I => \N__52345\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__52345\,
            I => \N__52340\
        );

    \I__11544\ : InMux
    port map (
            O => \N__52344\,
            I => \N__52335\
        );

    \I__11543\ : InMux
    port map (
            O => \N__52343\,
            I => \N__52335\
        );

    \I__11542\ : Odrv12
    port map (
            O => \N__52340\,
            I => \c0.n21170\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__52335\,
            I => \c0.n21170\
        );

    \I__11540\ : InMux
    port map (
            O => \N__52330\,
            I => \N__52326\
        );

    \I__11539\ : CascadeMux
    port map (
            O => \N__52329\,
            I => \N__52323\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__52326\,
            I => \N__52320\
        );

    \I__11537\ : InMux
    port map (
            O => \N__52323\,
            I => \N__52317\
        );

    \I__11536\ : Span4Mux_h
    port map (
            O => \N__52320\,
            I => \N__52314\
        );

    \I__11535\ : LocalMux
    port map (
            O => \N__52317\,
            I => \c0.n13974\
        );

    \I__11534\ : Odrv4
    port map (
            O => \N__52314\,
            I => \c0.n13974\
        );

    \I__11533\ : InMux
    port map (
            O => \N__52309\,
            I => \N__52306\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__52306\,
            I => \c0.n22245\
        );

    \I__11531\ : CascadeMux
    port map (
            O => \N__52303\,
            I => \N__52300\
        );

    \I__11530\ : InMux
    port map (
            O => \N__52300\,
            I => \N__52297\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__52297\,
            I => \N__52294\
        );

    \I__11528\ : Odrv4
    port map (
            O => \N__52294\,
            I => \c0.n22379\
        );

    \I__11527\ : CascadeMux
    port map (
            O => \N__52291\,
            I => \N__52288\
        );

    \I__11526\ : InMux
    port map (
            O => \N__52288\,
            I => \N__52285\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__52285\,
            I => \c0.n38_adj_4260\
        );

    \I__11524\ : InMux
    port map (
            O => \N__52282\,
            I => \N__52279\
        );

    \I__11523\ : LocalMux
    port map (
            O => \N__52279\,
            I => \c0.n6_adj_4256\
        );

    \I__11522\ : InMux
    port map (
            O => \N__52276\,
            I => \N__52271\
        );

    \I__11521\ : CascadeMux
    port map (
            O => \N__52275\,
            I => \N__52268\
        );

    \I__11520\ : InMux
    port map (
            O => \N__52274\,
            I => \N__52265\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__52271\,
            I => \N__52262\
        );

    \I__11518\ : InMux
    port map (
            O => \N__52268\,
            I => \N__52259\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__52265\,
            I => \N__52256\
        );

    \I__11516\ : Span4Mux_v
    port map (
            O => \N__52262\,
            I => \N__52253\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__52259\,
            I => \c0.data_in_frame_7_3\
        );

    \I__11514\ : Odrv4
    port map (
            O => \N__52256\,
            I => \c0.data_in_frame_7_3\
        );

    \I__11513\ : Odrv4
    port map (
            O => \N__52253\,
            I => \c0.data_in_frame_7_3\
        );

    \I__11512\ : CascadeMux
    port map (
            O => \N__52246\,
            I => \N__52243\
        );

    \I__11511\ : InMux
    port map (
            O => \N__52243\,
            I => \N__52240\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__52240\,
            I => \N__52237\
        );

    \I__11509\ : Span4Mux_v
    port map (
            O => \N__52237\,
            I => \N__52234\
        );

    \I__11508\ : Span4Mux_v
    port map (
            O => \N__52234\,
            I => \N__52230\
        );

    \I__11507\ : InMux
    port map (
            O => \N__52233\,
            I => \N__52226\
        );

    \I__11506\ : Span4Mux_h
    port map (
            O => \N__52230\,
            I => \N__52223\
        );

    \I__11505\ : InMux
    port map (
            O => \N__52229\,
            I => \N__52220\
        );

    \I__11504\ : LocalMux
    port map (
            O => \N__52226\,
            I => \N__52217\
        );

    \I__11503\ : Odrv4
    port map (
            O => \N__52223\,
            I => \c0.n13488\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__52220\,
            I => \c0.n13488\
        );

    \I__11501\ : Odrv4
    port map (
            O => \N__52217\,
            I => \c0.n13488\
        );

    \I__11500\ : CascadeMux
    port map (
            O => \N__52210\,
            I => \c0.n22139_cascade_\
        );

    \I__11499\ : CascadeMux
    port map (
            O => \N__52207\,
            I => \N__52203\
        );

    \I__11498\ : InMux
    port map (
            O => \N__52206\,
            I => \N__52199\
        );

    \I__11497\ : InMux
    port map (
            O => \N__52203\,
            I => \N__52196\
        );

    \I__11496\ : InMux
    port map (
            O => \N__52202\,
            I => \N__52193\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__52199\,
            I => \N__52190\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__52196\,
            I => \c0.data_in_frame_9_0\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__52193\,
            I => \c0.data_in_frame_9_0\
        );

    \I__11492\ : Odrv12
    port map (
            O => \N__52190\,
            I => \c0.data_in_frame_9_0\
        );

    \I__11491\ : InMux
    port map (
            O => \N__52183\,
            I => \N__52180\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__52180\,
            I => \N__52175\
        );

    \I__11489\ : InMux
    port map (
            O => \N__52179\,
            I => \N__52172\
        );

    \I__11488\ : InMux
    port map (
            O => \N__52178\,
            I => \N__52168\
        );

    \I__11487\ : Span4Mux_v
    port map (
            O => \N__52175\,
            I => \N__52165\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__52172\,
            I => \N__52162\
        );

    \I__11485\ : InMux
    port map (
            O => \N__52171\,
            I => \N__52159\
        );

    \I__11484\ : LocalMux
    port map (
            O => \N__52168\,
            I => \N__52156\
        );

    \I__11483\ : Span4Mux_h
    port map (
            O => \N__52165\,
            I => \N__52149\
        );

    \I__11482\ : Span4Mux_v
    port map (
            O => \N__52162\,
            I => \N__52149\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__52159\,
            I => \N__52149\
        );

    \I__11480\ : Odrv4
    port map (
            O => \N__52156\,
            I => \c0.n13605\
        );

    \I__11479\ : Odrv4
    port map (
            O => \N__52149\,
            I => \c0.n13605\
        );

    \I__11478\ : InMux
    port map (
            O => \N__52144\,
            I => \N__52138\
        );

    \I__11477\ : InMux
    port map (
            O => \N__52143\,
            I => \N__52138\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__52138\,
            I => \N__52135\
        );

    \I__11475\ : Span4Mux_h
    port map (
            O => \N__52135\,
            I => \N__52129\
        );

    \I__11474\ : InMux
    port map (
            O => \N__52134\,
            I => \N__52122\
        );

    \I__11473\ : InMux
    port map (
            O => \N__52133\,
            I => \N__52122\
        );

    \I__11472\ : InMux
    port map (
            O => \N__52132\,
            I => \N__52122\
        );

    \I__11471\ : Span4Mux_v
    port map (
            O => \N__52129\,
            I => \N__52119\
        );

    \I__11470\ : LocalMux
    port map (
            O => \N__52122\,
            I => \N__52116\
        );

    \I__11469\ : Odrv4
    port map (
            O => \N__52119\,
            I => \c0.n13043\
        );

    \I__11468\ : Odrv12
    port map (
            O => \N__52116\,
            I => \c0.n13043\
        );

    \I__11467\ : InMux
    port map (
            O => \N__52111\,
            I => \N__52108\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__52108\,
            I => \N__52102\
        );

    \I__11465\ : InMux
    port map (
            O => \N__52107\,
            I => \N__52099\
        );

    \I__11464\ : InMux
    port map (
            O => \N__52106\,
            I => \N__52095\
        );

    \I__11463\ : InMux
    port map (
            O => \N__52105\,
            I => \N__52092\
        );

    \I__11462\ : Span4Mux_v
    port map (
            O => \N__52102\,
            I => \N__52089\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__52099\,
            I => \N__52086\
        );

    \I__11460\ : InMux
    port map (
            O => \N__52098\,
            I => \N__52083\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__52095\,
            I => \c0.data_in_frame_8_6\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__52092\,
            I => \c0.data_in_frame_8_6\
        );

    \I__11457\ : Odrv4
    port map (
            O => \N__52089\,
            I => \c0.data_in_frame_8_6\
        );

    \I__11456\ : Odrv12
    port map (
            O => \N__52086\,
            I => \c0.data_in_frame_8_6\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__52083\,
            I => \c0.data_in_frame_8_6\
        );

    \I__11454\ : CascadeMux
    port map (
            O => \N__52072\,
            I => \c0.n21822_cascade_\
        );

    \I__11453\ : InMux
    port map (
            O => \N__52069\,
            I => \N__52065\
        );

    \I__11452\ : CascadeMux
    port map (
            O => \N__52068\,
            I => \N__52062\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__52065\,
            I => \N__52059\
        );

    \I__11450\ : InMux
    port map (
            O => \N__52062\,
            I => \N__52055\
        );

    \I__11449\ : Span4Mux_h
    port map (
            O => \N__52059\,
            I => \N__52051\
        );

    \I__11448\ : CascadeMux
    port map (
            O => \N__52058\,
            I => \N__52047\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__52055\,
            I => \N__52044\
        );

    \I__11446\ : InMux
    port map (
            O => \N__52054\,
            I => \N__52041\
        );

    \I__11445\ : Sp12to4
    port map (
            O => \N__52051\,
            I => \N__52038\
        );

    \I__11444\ : InMux
    port map (
            O => \N__52050\,
            I => \N__52035\
        );

    \I__11443\ : InMux
    port map (
            O => \N__52047\,
            I => \N__52031\
        );

    \I__11442\ : Span4Mux_v
    port map (
            O => \N__52044\,
            I => \N__52028\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__52041\,
            I => \N__52025\
        );

    \I__11440\ : Span12Mux_v
    port map (
            O => \N__52038\,
            I => \N__52020\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__52035\,
            I => \N__52020\
        );

    \I__11438\ : InMux
    port map (
            O => \N__52034\,
            I => \N__52017\
        );

    \I__11437\ : LocalMux
    port map (
            O => \N__52031\,
            I => data_in_frame_1_2
        );

    \I__11436\ : Odrv4
    port map (
            O => \N__52028\,
            I => data_in_frame_1_2
        );

    \I__11435\ : Odrv4
    port map (
            O => \N__52025\,
            I => data_in_frame_1_2
        );

    \I__11434\ : Odrv12
    port map (
            O => \N__52020\,
            I => data_in_frame_1_2
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__52017\,
            I => data_in_frame_1_2
        );

    \I__11432\ : InMux
    port map (
            O => \N__52006\,
            I => \N__52003\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__52003\,
            I => \c0.n22334\
        );

    \I__11430\ : CascadeMux
    port map (
            O => \N__52000\,
            I => \c0.n22334_cascade_\
        );

    \I__11429\ : InMux
    port map (
            O => \N__51997\,
            I => \N__51991\
        );

    \I__11428\ : InMux
    port map (
            O => \N__51996\,
            I => \N__51991\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__51991\,
            I => \N__51987\
        );

    \I__11426\ : InMux
    port map (
            O => \N__51990\,
            I => \N__51984\
        );

    \I__11425\ : Odrv4
    port map (
            O => \N__51987\,
            I => \c0.n22051\
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__51984\,
            I => \c0.n22051\
        );

    \I__11423\ : InMux
    port map (
            O => \N__51979\,
            I => \N__51975\
        );

    \I__11422\ : InMux
    port map (
            O => \N__51978\,
            I => \N__51971\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__51975\,
            I => \N__51967\
        );

    \I__11420\ : InMux
    port map (
            O => \N__51974\,
            I => \N__51964\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__51971\,
            I => \N__51961\
        );

    \I__11418\ : InMux
    port map (
            O => \N__51970\,
            I => \N__51958\
        );

    \I__11417\ : Span4Mux_h
    port map (
            O => \N__51967\,
            I => \N__51953\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__51964\,
            I => \N__51953\
        );

    \I__11415\ : Span4Mux_h
    port map (
            O => \N__51961\,
            I => \N__51950\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__51958\,
            I => \c0.n15_adj_4404\
        );

    \I__11413\ : Odrv4
    port map (
            O => \N__51953\,
            I => \c0.n15_adj_4404\
        );

    \I__11412\ : Odrv4
    port map (
            O => \N__51950\,
            I => \c0.n15_adj_4404\
        );

    \I__11411\ : InMux
    port map (
            O => \N__51943\,
            I => \N__51939\
        );

    \I__11410\ : CascadeMux
    port map (
            O => \N__51942\,
            I => \N__51935\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__51939\,
            I => \N__51932\
        );

    \I__11408\ : InMux
    port map (
            O => \N__51938\,
            I => \N__51927\
        );

    \I__11407\ : InMux
    port map (
            O => \N__51935\,
            I => \N__51927\
        );

    \I__11406\ : Span4Mux_v
    port map (
            O => \N__51932\,
            I => \N__51924\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__51927\,
            I => \c0.data_in_frame_8_0\
        );

    \I__11404\ : Odrv4
    port map (
            O => \N__51924\,
            I => \c0.data_in_frame_8_0\
        );

    \I__11403\ : CascadeMux
    port map (
            O => \N__51919\,
            I => \N__51915\
        );

    \I__11402\ : CascadeMux
    port map (
            O => \N__51918\,
            I => \N__51911\
        );

    \I__11401\ : InMux
    port map (
            O => \N__51915\,
            I => \N__51907\
        );

    \I__11400\ : InMux
    port map (
            O => \N__51914\,
            I => \N__51904\
        );

    \I__11399\ : InMux
    port map (
            O => \N__51911\,
            I => \N__51899\
        );

    \I__11398\ : InMux
    port map (
            O => \N__51910\,
            I => \N__51899\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__51907\,
            I => \c0.data_in_frame_7_7\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__51904\,
            I => \c0.data_in_frame_7_7\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__51899\,
            I => \c0.data_in_frame_7_7\
        );

    \I__11394\ : InMux
    port map (
            O => \N__51892\,
            I => \N__51889\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__51889\,
            I => \c0.n6_adj_4259\
        );

    \I__11392\ : InMux
    port map (
            O => \N__51886\,
            I => \N__51883\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__51883\,
            I => \N__51880\
        );

    \I__11390\ : Odrv4
    port map (
            O => \N__51880\,
            I => \c0.n39_adj_4263\
        );

    \I__11389\ : InMux
    port map (
            O => \N__51877\,
            I => \N__51874\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__51874\,
            I => \N__51871\
        );

    \I__11387\ : Odrv4
    port map (
            O => \N__51871\,
            I => \c0.n40_adj_4261\
        );

    \I__11386\ : CascadeMux
    port map (
            O => \N__51868\,
            I => \c0.n22060_cascade_\
        );

    \I__11385\ : InMux
    port map (
            O => \N__51865\,
            I => \N__51862\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__51862\,
            I => \c0.n44_adj_4262\
        );

    \I__11383\ : CascadeMux
    port map (
            O => \N__51859\,
            I => \c0.n11_adj_4266_cascade_\
        );

    \I__11382\ : InMux
    port map (
            O => \N__51856\,
            I => \N__51851\
        );

    \I__11381\ : InMux
    port map (
            O => \N__51855\,
            I => \N__51846\
        );

    \I__11380\ : InMux
    port map (
            O => \N__51854\,
            I => \N__51846\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__51851\,
            I => \c0.n13425\
        );

    \I__11378\ : LocalMux
    port map (
            O => \N__51846\,
            I => \c0.n13425\
        );

    \I__11377\ : CascadeMux
    port map (
            O => \N__51841\,
            I => \c0.n22842_cascade_\
        );

    \I__11376\ : InMux
    port map (
            O => \N__51838\,
            I => \N__51833\
        );

    \I__11375\ : InMux
    port map (
            O => \N__51837\,
            I => \N__51830\
        );

    \I__11374\ : InMux
    port map (
            O => \N__51836\,
            I => \N__51827\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__51833\,
            I => \c0.data_in_frame_5_6\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__51830\,
            I => \c0.data_in_frame_5_6\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__51827\,
            I => \c0.data_in_frame_5_6\
        );

    \I__11370\ : InMux
    port map (
            O => \N__51820\,
            I => \N__51816\
        );

    \I__11369\ : InMux
    port map (
            O => \N__51819\,
            I => \N__51813\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__51816\,
            I => \N__51810\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__51813\,
            I => \c0.n22283\
        );

    \I__11366\ : Odrv12
    port map (
            O => \N__51810\,
            I => \c0.n22283\
        );

    \I__11365\ : CascadeMux
    port map (
            O => \N__51805\,
            I => \c0.n13488_cascade_\
        );

    \I__11364\ : InMux
    port map (
            O => \N__51802\,
            I => \N__51797\
        );

    \I__11363\ : InMux
    port map (
            O => \N__51801\,
            I => \N__51794\
        );

    \I__11362\ : InMux
    port map (
            O => \N__51800\,
            I => \N__51791\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__51797\,
            I => \N__51788\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__51794\,
            I => \N__51785\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__51791\,
            I => \c0.n13180\
        );

    \I__11358\ : Odrv12
    port map (
            O => \N__51788\,
            I => \c0.n13180\
        );

    \I__11357\ : Odrv12
    port map (
            O => \N__51785\,
            I => \c0.n13180\
        );

    \I__11356\ : InMux
    port map (
            O => \N__51778\,
            I => \N__51768\
        );

    \I__11355\ : InMux
    port map (
            O => \N__51777\,
            I => \N__51768\
        );

    \I__11354\ : InMux
    port map (
            O => \N__51776\,
            I => \N__51765\
        );

    \I__11353\ : InMux
    port map (
            O => \N__51775\,
            I => \N__51762\
        );

    \I__11352\ : InMux
    port map (
            O => \N__51774\,
            I => \N__51759\
        );

    \I__11351\ : CascadeMux
    port map (
            O => \N__51773\,
            I => \N__51756\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__51768\,
            I => \N__51750\
        );

    \I__11349\ : LocalMux
    port map (
            O => \N__51765\,
            I => \N__51747\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__51762\,
            I => \N__51744\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__51759\,
            I => \N__51741\
        );

    \I__11346\ : InMux
    port map (
            O => \N__51756\,
            I => \N__51738\
        );

    \I__11345\ : InMux
    port map (
            O => \N__51755\,
            I => \N__51733\
        );

    \I__11344\ : InMux
    port map (
            O => \N__51754\,
            I => \N__51733\
        );

    \I__11343\ : InMux
    port map (
            O => \N__51753\,
            I => \N__51730\
        );

    \I__11342\ : Span4Mux_h
    port map (
            O => \N__51750\,
            I => \N__51721\
        );

    \I__11341\ : Span4Mux_v
    port map (
            O => \N__51747\,
            I => \N__51721\
        );

    \I__11340\ : Span4Mux_h
    port map (
            O => \N__51744\,
            I => \N__51721\
        );

    \I__11339\ : Span4Mux_v
    port map (
            O => \N__51741\,
            I => \N__51721\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__51738\,
            I => \c0.data_in_frame_0_5\
        );

    \I__11337\ : LocalMux
    port map (
            O => \N__51733\,
            I => \c0.data_in_frame_0_5\
        );

    \I__11336\ : LocalMux
    port map (
            O => \N__51730\,
            I => \c0.data_in_frame_0_5\
        );

    \I__11335\ : Odrv4
    port map (
            O => \N__51721\,
            I => \c0.data_in_frame_0_5\
        );

    \I__11334\ : InMux
    port map (
            O => \N__51712\,
            I => \N__51707\
        );

    \I__11333\ : InMux
    port map (
            O => \N__51711\,
            I => \N__51704\
        );

    \I__11332\ : InMux
    port map (
            O => \N__51710\,
            I => \N__51701\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__51707\,
            I => \N__51697\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__51704\,
            I => \N__51694\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__51701\,
            I => \N__51691\
        );

    \I__11328\ : InMux
    port map (
            O => \N__51700\,
            I => \N__51688\
        );

    \I__11327\ : Span4Mux_h
    port map (
            O => \N__51697\,
            I => \N__51680\
        );

    \I__11326\ : Span4Mux_v
    port map (
            O => \N__51694\,
            I => \N__51673\
        );

    \I__11325\ : Span4Mux_h
    port map (
            O => \N__51691\,
            I => \N__51673\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__51688\,
            I => \N__51673\
        );

    \I__11323\ : InMux
    port map (
            O => \N__51687\,
            I => \N__51670\
        );

    \I__11322\ : InMux
    port map (
            O => \N__51686\,
            I => \N__51665\
        );

    \I__11321\ : InMux
    port map (
            O => \N__51685\,
            I => \N__51665\
        );

    \I__11320\ : InMux
    port map (
            O => \N__51684\,
            I => \N__51660\
        );

    \I__11319\ : InMux
    port map (
            O => \N__51683\,
            I => \N__51660\
        );

    \I__11318\ : Odrv4
    port map (
            O => \N__51680\,
            I => \c0.data_in_frame_0_6\
        );

    \I__11317\ : Odrv4
    port map (
            O => \N__51673\,
            I => \c0.data_in_frame_0_6\
        );

    \I__11316\ : LocalMux
    port map (
            O => \N__51670\,
            I => \c0.data_in_frame_0_6\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__51665\,
            I => \c0.data_in_frame_0_6\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__51660\,
            I => \c0.data_in_frame_0_6\
        );

    \I__11313\ : CascadeMux
    port map (
            O => \N__51649\,
            I => \N__51646\
        );

    \I__11312\ : InMux
    port map (
            O => \N__51646\,
            I => \N__51643\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__51643\,
            I => \N__51640\
        );

    \I__11310\ : Span4Mux_h
    port map (
            O => \N__51640\,
            I => \N__51637\
        );

    \I__11309\ : Span4Mux_v
    port map (
            O => \N__51637\,
            I => \N__51634\
        );

    \I__11308\ : Odrv4
    port map (
            O => \N__51634\,
            I => \c0.n23827\
        );

    \I__11307\ : InMux
    port map (
            O => \N__51631\,
            I => \N__51627\
        );

    \I__11306\ : CascadeMux
    port map (
            O => \N__51630\,
            I => \N__51624\
        );

    \I__11305\ : LocalMux
    port map (
            O => \N__51627\,
            I => \N__51619\
        );

    \I__11304\ : InMux
    port map (
            O => \N__51624\,
            I => \N__51616\
        );

    \I__11303\ : InMux
    port map (
            O => \N__51623\,
            I => \N__51613\
        );

    \I__11302\ : InMux
    port map (
            O => \N__51622\,
            I => \N__51610\
        );

    \I__11301\ : Sp12to4
    port map (
            O => \N__51619\,
            I => \N__51607\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__51616\,
            I => \c0.data_in_frame_5_3\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__51613\,
            I => \c0.data_in_frame_5_3\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__51610\,
            I => \c0.data_in_frame_5_3\
        );

    \I__11297\ : Odrv12
    port map (
            O => \N__51607\,
            I => \c0.data_in_frame_5_3\
        );

    \I__11296\ : CascadeMux
    port map (
            O => \N__51598\,
            I => \N__51593\
        );

    \I__11295\ : CascadeMux
    port map (
            O => \N__51597\,
            I => \N__51589\
        );

    \I__11294\ : InMux
    port map (
            O => \N__51596\,
            I => \N__51586\
        );

    \I__11293\ : InMux
    port map (
            O => \N__51593\,
            I => \N__51581\
        );

    \I__11292\ : InMux
    port map (
            O => \N__51592\,
            I => \N__51581\
        );

    \I__11291\ : InMux
    port map (
            O => \N__51589\,
            I => \N__51578\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__51586\,
            I => \c0.data_in_frame_7_5\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__51581\,
            I => \c0.data_in_frame_7_5\
        );

    \I__11288\ : LocalMux
    port map (
            O => \N__51578\,
            I => \c0.data_in_frame_7_5\
        );

    \I__11287\ : InMux
    port map (
            O => \N__51571\,
            I => \N__51568\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__51568\,
            I => \N__51563\
        );

    \I__11285\ : InMux
    port map (
            O => \N__51567\,
            I => \N__51560\
        );

    \I__11284\ : InMux
    port map (
            O => \N__51566\,
            I => \N__51557\
        );

    \I__11283\ : Odrv4
    port map (
            O => \N__51563\,
            I => \c0.n12484\
        );

    \I__11282\ : LocalMux
    port map (
            O => \N__51560\,
            I => \c0.n12484\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__51557\,
            I => \c0.n12484\
        );

    \I__11280\ : CascadeMux
    port map (
            O => \N__51550\,
            I => \c0.n20368_cascade_\
        );

    \I__11279\ : CascadeMux
    port map (
            O => \N__51547\,
            I => \N__51544\
        );

    \I__11278\ : InMux
    port map (
            O => \N__51544\,
            I => \N__51540\
        );

    \I__11277\ : InMux
    port map (
            O => \N__51543\,
            I => \N__51537\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__51540\,
            I => \N__51534\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__51537\,
            I => \N__51531\
        );

    \I__11274\ : Odrv4
    port map (
            O => \N__51534\,
            I => \c0.data_in_frame_10_1\
        );

    \I__11273\ : Odrv4
    port map (
            O => \N__51531\,
            I => \c0.data_in_frame_10_1\
        );

    \I__11272\ : CascadeMux
    port map (
            O => \N__51526\,
            I => \c0.n22133_cascade_\
        );

    \I__11271\ : InMux
    port map (
            O => \N__51523\,
            I => \N__51520\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__51520\,
            I => \c0.n21925\
        );

    \I__11269\ : CascadeMux
    port map (
            O => \N__51517\,
            I => \c0.n20927_cascade_\
        );

    \I__11268\ : InMux
    port map (
            O => \N__51514\,
            I => \N__51511\
        );

    \I__11267\ : LocalMux
    port map (
            O => \N__51511\,
            I => \c0.n22133\
        );

    \I__11266\ : InMux
    port map (
            O => \N__51508\,
            I => \N__51505\
        );

    \I__11265\ : LocalMux
    port map (
            O => \N__51505\,
            I => \c0.n36\
        );

    \I__11264\ : InMux
    port map (
            O => \N__51502\,
            I => \c0.rx.n19539\
        );

    \I__11263\ : CEMux
    port map (
            O => \N__51499\,
            I => \N__51496\
        );

    \I__11262\ : LocalMux
    port map (
            O => \N__51496\,
            I => \N__51493\
        );

    \I__11261\ : Span4Mux_h
    port map (
            O => \N__51493\,
            I => \N__51490\
        );

    \I__11260\ : Span4Mux_h
    port map (
            O => \N__51490\,
            I => \N__51487\
        );

    \I__11259\ : Odrv4
    port map (
            O => \N__51487\,
            I => \c0.rx.n14391\
        );

    \I__11258\ : SRMux
    port map (
            O => \N__51484\,
            I => \N__51481\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__51481\,
            I => \N__51478\
        );

    \I__11256\ : Odrv12
    port map (
            O => \N__51478\,
            I => \c0.rx.n17411\
        );

    \I__11255\ : InMux
    port map (
            O => \N__51475\,
            I => \N__51467\
        );

    \I__11254\ : InMux
    port map (
            O => \N__51474\,
            I => \N__51458\
        );

    \I__11253\ : InMux
    port map (
            O => \N__51473\,
            I => \N__51458\
        );

    \I__11252\ : InMux
    port map (
            O => \N__51472\,
            I => \N__51455\
        );

    \I__11251\ : InMux
    port map (
            O => \N__51471\,
            I => \N__51452\
        );

    \I__11250\ : InMux
    port map (
            O => \N__51470\,
            I => \N__51445\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__51467\,
            I => \N__51440\
        );

    \I__11248\ : InMux
    port map (
            O => \N__51466\,
            I => \N__51437\
        );

    \I__11247\ : InMux
    port map (
            O => \N__51465\,
            I => \N__51426\
        );

    \I__11246\ : InMux
    port map (
            O => \N__51464\,
            I => \N__51426\
        );

    \I__11245\ : InMux
    port map (
            O => \N__51463\,
            I => \N__51426\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__51458\,
            I => \N__51423\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__51455\,
            I => \N__51420\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__51452\,
            I => \N__51417\
        );

    \I__11241\ : InMux
    port map (
            O => \N__51451\,
            I => \N__51414\
        );

    \I__11240\ : InMux
    port map (
            O => \N__51450\,
            I => \N__51404\
        );

    \I__11239\ : InMux
    port map (
            O => \N__51449\,
            I => \N__51404\
        );

    \I__11238\ : InMux
    port map (
            O => \N__51448\,
            I => \N__51399\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__51445\,
            I => \N__51395\
        );

    \I__11236\ : InMux
    port map (
            O => \N__51444\,
            I => \N__51390\
        );

    \I__11235\ : InMux
    port map (
            O => \N__51443\,
            I => \N__51390\
        );

    \I__11234\ : Span4Mux_h
    port map (
            O => \N__51440\,
            I => \N__51383\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__51437\,
            I => \N__51383\
        );

    \I__11232\ : InMux
    port map (
            O => \N__51436\,
            I => \N__51380\
        );

    \I__11231\ : InMux
    port map (
            O => \N__51435\,
            I => \N__51373\
        );

    \I__11230\ : InMux
    port map (
            O => \N__51434\,
            I => \N__51373\
        );

    \I__11229\ : InMux
    port map (
            O => \N__51433\,
            I => \N__51373\
        );

    \I__11228\ : LocalMux
    port map (
            O => \N__51426\,
            I => \N__51368\
        );

    \I__11227\ : Span4Mux_v
    port map (
            O => \N__51423\,
            I => \N__51363\
        );

    \I__11226\ : Span4Mux_h
    port map (
            O => \N__51420\,
            I => \N__51356\
        );

    \I__11225\ : Span4Mux_v
    port map (
            O => \N__51417\,
            I => \N__51356\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__51414\,
            I => \N__51356\
        );

    \I__11223\ : InMux
    port map (
            O => \N__51413\,
            I => \N__51351\
        );

    \I__11222\ : InMux
    port map (
            O => \N__51412\,
            I => \N__51351\
        );

    \I__11221\ : InMux
    port map (
            O => \N__51411\,
            I => \N__51348\
        );

    \I__11220\ : InMux
    port map (
            O => \N__51410\,
            I => \N__51343\
        );

    \I__11219\ : InMux
    port map (
            O => \N__51409\,
            I => \N__51343\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__51404\,
            I => \N__51340\
        );

    \I__11217\ : InMux
    port map (
            O => \N__51403\,
            I => \N__51335\
        );

    \I__11216\ : InMux
    port map (
            O => \N__51402\,
            I => \N__51335\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__51399\,
            I => \N__51332\
        );

    \I__11214\ : InMux
    port map (
            O => \N__51398\,
            I => \N__51329\
        );

    \I__11213\ : Span4Mux_h
    port map (
            O => \N__51395\,
            I => \N__51326\
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__51390\,
            I => \N__51323\
        );

    \I__11211\ : InMux
    port map (
            O => \N__51389\,
            I => \N__51317\
        );

    \I__11210\ : InMux
    port map (
            O => \N__51388\,
            I => \N__51317\
        );

    \I__11209\ : Span4Mux_v
    port map (
            O => \N__51383\,
            I => \N__51312\
        );

    \I__11208\ : LocalMux
    port map (
            O => \N__51380\,
            I => \N__51312\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__51373\,
            I => \N__51309\
        );

    \I__11206\ : InMux
    port map (
            O => \N__51372\,
            I => \N__51304\
        );

    \I__11205\ : InMux
    port map (
            O => \N__51371\,
            I => \N__51304\
        );

    \I__11204\ : Span4Mux_h
    port map (
            O => \N__51368\,
            I => \N__51301\
        );

    \I__11203\ : InMux
    port map (
            O => \N__51367\,
            I => \N__51296\
        );

    \I__11202\ : InMux
    port map (
            O => \N__51366\,
            I => \N__51296\
        );

    \I__11201\ : Sp12to4
    port map (
            O => \N__51363\,
            I => \N__51293\
        );

    \I__11200\ : Span4Mux_h
    port map (
            O => \N__51356\,
            I => \N__51290\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__51351\,
            I => \N__51287\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__51348\,
            I => \N__51282\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__51343\,
            I => \N__51282\
        );

    \I__11196\ : Span4Mux_v
    port map (
            O => \N__51340\,
            I => \N__51277\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__51335\,
            I => \N__51277\
        );

    \I__11194\ : Span4Mux_v
    port map (
            O => \N__51332\,
            I => \N__51272\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__51329\,
            I => \N__51272\
        );

    \I__11192\ : Span4Mux_h
    port map (
            O => \N__51326\,
            I => \N__51267\
        );

    \I__11191\ : Span4Mux_h
    port map (
            O => \N__51323\,
            I => \N__51267\
        );

    \I__11190\ : InMux
    port map (
            O => \N__51322\,
            I => \N__51264\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__51317\,
            I => \N__51257\
        );

    \I__11188\ : Span4Mux_v
    port map (
            O => \N__51312\,
            I => \N__51257\
        );

    \I__11187\ : Span4Mux_v
    port map (
            O => \N__51309\,
            I => \N__51257\
        );

    \I__11186\ : LocalMux
    port map (
            O => \N__51304\,
            I => \N__51250\
        );

    \I__11185\ : Span4Mux_h
    port map (
            O => \N__51301\,
            I => \N__51250\
        );

    \I__11184\ : LocalMux
    port map (
            O => \N__51296\,
            I => \N__51250\
        );

    \I__11183\ : Span12Mux_h
    port map (
            O => \N__51293\,
            I => \N__51247\
        );

    \I__11182\ : Sp12to4
    port map (
            O => \N__51290\,
            I => \N__51244\
        );

    \I__11181\ : Span4Mux_v
    port map (
            O => \N__51287\,
            I => \N__51239\
        );

    \I__11180\ : Span4Mux_v
    port map (
            O => \N__51282\,
            I => \N__51239\
        );

    \I__11179\ : Span4Mux_h
    port map (
            O => \N__51277\,
            I => \N__51236\
        );

    \I__11178\ : Span4Mux_h
    port map (
            O => \N__51272\,
            I => \N__51231\
        );

    \I__11177\ : Span4Mux_v
    port map (
            O => \N__51267\,
            I => \N__51231\
        );

    \I__11176\ : LocalMux
    port map (
            O => \N__51264\,
            I => \N__51224\
        );

    \I__11175\ : Span4Mux_h
    port map (
            O => \N__51257\,
            I => \N__51224\
        );

    \I__11174\ : Span4Mux_v
    port map (
            O => \N__51250\,
            I => \N__51224\
        );

    \I__11173\ : Span12Mux_v
    port map (
            O => \N__51247\,
            I => \N__51221\
        );

    \I__11172\ : Span12Mux_s10_v
    port map (
            O => \N__51244\,
            I => \N__51218\
        );

    \I__11171\ : Odrv4
    port map (
            O => \N__51239\,
            I => \c0.data_out_frame_29_7_N_1483_0\
        );

    \I__11170\ : Odrv4
    port map (
            O => \N__51236\,
            I => \c0.data_out_frame_29_7_N_1483_0\
        );

    \I__11169\ : Odrv4
    port map (
            O => \N__51231\,
            I => \c0.data_out_frame_29_7_N_1483_0\
        );

    \I__11168\ : Odrv4
    port map (
            O => \N__51224\,
            I => \c0.data_out_frame_29_7_N_1483_0\
        );

    \I__11167\ : Odrv12
    port map (
            O => \N__51221\,
            I => \c0.data_out_frame_29_7_N_1483_0\
        );

    \I__11166\ : Odrv12
    port map (
            O => \N__51218\,
            I => \c0.data_out_frame_29_7_N_1483_0\
        );

    \I__11165\ : InMux
    port map (
            O => \N__51205\,
            I => \N__51200\
        );

    \I__11164\ : InMux
    port map (
            O => \N__51204\,
            I => \N__51197\
        );

    \I__11163\ : InMux
    port map (
            O => \N__51203\,
            I => \N__51194\
        );

    \I__11162\ : LocalMux
    port map (
            O => \N__51200\,
            I => \N__51182\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__51197\,
            I => \N__51182\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__51194\,
            I => \N__51182\
        );

    \I__11159\ : InMux
    port map (
            O => \N__51193\,
            I => \N__51179\
        );

    \I__11158\ : InMux
    port map (
            O => \N__51192\,
            I => \N__51176\
        );

    \I__11157\ : InMux
    port map (
            O => \N__51191\,
            I => \N__51169\
        );

    \I__11156\ : InMux
    port map (
            O => \N__51190\,
            I => \N__51166\
        );

    \I__11155\ : InMux
    port map (
            O => \N__51189\,
            I => \N__51163\
        );

    \I__11154\ : Span4Mux_v
    port map (
            O => \N__51182\,
            I => \N__51151\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__51179\,
            I => \N__51151\
        );

    \I__11152\ : LocalMux
    port map (
            O => \N__51176\,
            I => \N__51151\
        );

    \I__11151\ : InMux
    port map (
            O => \N__51175\,
            I => \N__51148\
        );

    \I__11150\ : InMux
    port map (
            O => \N__51174\,
            I => \N__51145\
        );

    \I__11149\ : InMux
    port map (
            O => \N__51173\,
            I => \N__51142\
        );

    \I__11148\ : InMux
    port map (
            O => \N__51172\,
            I => \N__51139\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__51169\,
            I => \N__51132\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__51166\,
            I => \N__51132\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__51163\,
            I => \N__51132\
        );

    \I__11144\ : InMux
    port map (
            O => \N__51162\,
            I => \N__51127\
        );

    \I__11143\ : InMux
    port map (
            O => \N__51161\,
            I => \N__51124\
        );

    \I__11142\ : InMux
    port map (
            O => \N__51160\,
            I => \N__51119\
        );

    \I__11141\ : InMux
    port map (
            O => \N__51159\,
            I => \N__51114\
        );

    \I__11140\ : InMux
    port map (
            O => \N__51158\,
            I => \N__51114\
        );

    \I__11139\ : Span4Mux_v
    port map (
            O => \N__51151\,
            I => \N__51104\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__51148\,
            I => \N__51104\
        );

    \I__11137\ : LocalMux
    port map (
            O => \N__51145\,
            I => \N__51104\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__51142\,
            I => \N__51101\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__51139\,
            I => \N__51093\
        );

    \I__11134\ : Span4Mux_h
    port map (
            O => \N__51132\,
            I => \N__51090\
        );

    \I__11133\ : InMux
    port map (
            O => \N__51131\,
            I => \N__51082\
        );

    \I__11132\ : InMux
    port map (
            O => \N__51130\,
            I => \N__51079\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__51127\,
            I => \N__51074\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__51124\,
            I => \N__51074\
        );

    \I__11129\ : InMux
    port map (
            O => \N__51123\,
            I => \N__51071\
        );

    \I__11128\ : InMux
    port map (
            O => \N__51122\,
            I => \N__51061\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__51119\,
            I => \N__51056\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__51114\,
            I => \N__51056\
        );

    \I__11125\ : InMux
    port map (
            O => \N__51113\,
            I => \N__51049\
        );

    \I__11124\ : InMux
    port map (
            O => \N__51112\,
            I => \N__51046\
        );

    \I__11123\ : CascadeMux
    port map (
            O => \N__51111\,
            I => \N__51043\
        );

    \I__11122\ : Span4Mux_v
    port map (
            O => \N__51104\,
            I => \N__51036\
        );

    \I__11121\ : Span4Mux_s1_v
    port map (
            O => \N__51101\,
            I => \N__51036\
        );

    \I__11120\ : InMux
    port map (
            O => \N__51100\,
            I => \N__51033\
        );

    \I__11119\ : InMux
    port map (
            O => \N__51099\,
            I => \N__51030\
        );

    \I__11118\ : InMux
    port map (
            O => \N__51098\,
            I => \N__51027\
        );

    \I__11117\ : InMux
    port map (
            O => \N__51097\,
            I => \N__51024\
        );

    \I__11116\ : InMux
    port map (
            O => \N__51096\,
            I => \N__51021\
        );

    \I__11115\ : Span4Mux_h
    port map (
            O => \N__51093\,
            I => \N__51016\
        );

    \I__11114\ : Span4Mux_v
    port map (
            O => \N__51090\,
            I => \N__51016\
        );

    \I__11113\ : CascadeMux
    port map (
            O => \N__51089\,
            I => \N__51013\
        );

    \I__11112\ : InMux
    port map (
            O => \N__51088\,
            I => \N__51007\
        );

    \I__11111\ : InMux
    port map (
            O => \N__51087\,
            I => \N__51004\
        );

    \I__11110\ : InMux
    port map (
            O => \N__51086\,
            I => \N__51001\
        );

    \I__11109\ : InMux
    port map (
            O => \N__51085\,
            I => \N__50998\
        );

    \I__11108\ : LocalMux
    port map (
            O => \N__51082\,
            I => \N__50995\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__51079\,
            I => \N__50988\
        );

    \I__11106\ : Span4Mux_s2_v
    port map (
            O => \N__51074\,
            I => \N__50988\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__51071\,
            I => \N__50988\
        );

    \I__11104\ : CascadeMux
    port map (
            O => \N__51070\,
            I => \N__50984\
        );

    \I__11103\ : InMux
    port map (
            O => \N__51069\,
            I => \N__50981\
        );

    \I__11102\ : InMux
    port map (
            O => \N__51068\,
            I => \N__50975\
        );

    \I__11101\ : InMux
    port map (
            O => \N__51067\,
            I => \N__50975\
        );

    \I__11100\ : CascadeMux
    port map (
            O => \N__51066\,
            I => \N__50970\
        );

    \I__11099\ : CascadeMux
    port map (
            O => \N__51065\,
            I => \N__50966\
        );

    \I__11098\ : InMux
    port map (
            O => \N__51064\,
            I => \N__50963\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__51061\,
            I => \N__50956\
        );

    \I__11096\ : Span4Mux_h
    port map (
            O => \N__51056\,
            I => \N__50956\
        );

    \I__11095\ : InMux
    port map (
            O => \N__51055\,
            I => \N__50951\
        );

    \I__11094\ : InMux
    port map (
            O => \N__51054\,
            I => \N__50948\
        );

    \I__11093\ : InMux
    port map (
            O => \N__51053\,
            I => \N__50945\
        );

    \I__11092\ : InMux
    port map (
            O => \N__51052\,
            I => \N__50942\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__51049\,
            I => \N__50937\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__51046\,
            I => \N__50937\
        );

    \I__11089\ : InMux
    port map (
            O => \N__51043\,
            I => \N__50930\
        );

    \I__11088\ : InMux
    port map (
            O => \N__51042\,
            I => \N__50930\
        );

    \I__11087\ : InMux
    port map (
            O => \N__51041\,
            I => \N__50930\
        );

    \I__11086\ : Sp12to4
    port map (
            O => \N__51036\,
            I => \N__50924\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__51033\,
            I => \N__50924\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__51030\,
            I => \N__50919\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__51027\,
            I => \N__50919\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__51024\,
            I => \N__50914\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__51021\,
            I => \N__50914\
        );

    \I__11080\ : Span4Mux_v
    port map (
            O => \N__51016\,
            I => \N__50911\
        );

    \I__11079\ : InMux
    port map (
            O => \N__51013\,
            I => \N__50904\
        );

    \I__11078\ : InMux
    port map (
            O => \N__51012\,
            I => \N__50904\
        );

    \I__11077\ : InMux
    port map (
            O => \N__51011\,
            I => \N__50904\
        );

    \I__11076\ : InMux
    port map (
            O => \N__51010\,
            I => \N__50901\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__51007\,
            I => \N__50888\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__51004\,
            I => \N__50888\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__51001\,
            I => \N__50888\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__50998\,
            I => \N__50888\
        );

    \I__11071\ : Span4Mux_v
    port map (
            O => \N__50995\,
            I => \N__50888\
        );

    \I__11070\ : Span4Mux_v
    port map (
            O => \N__50988\,
            I => \N__50888\
        );

    \I__11069\ : InMux
    port map (
            O => \N__50987\,
            I => \N__50883\
        );

    \I__11068\ : InMux
    port map (
            O => \N__50984\,
            I => \N__50883\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__50981\,
            I => \N__50880\
        );

    \I__11066\ : InMux
    port map (
            O => \N__50980\,
            I => \N__50877\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__50975\,
            I => \N__50874\
        );

    \I__11064\ : InMux
    port map (
            O => \N__50974\,
            I => \N__50871\
        );

    \I__11063\ : InMux
    port map (
            O => \N__50973\,
            I => \N__50866\
        );

    \I__11062\ : InMux
    port map (
            O => \N__50970\,
            I => \N__50866\
        );

    \I__11061\ : InMux
    port map (
            O => \N__50969\,
            I => \N__50861\
        );

    \I__11060\ : InMux
    port map (
            O => \N__50966\,
            I => \N__50861\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__50963\,
            I => \N__50858\
        );

    \I__11058\ : InMux
    port map (
            O => \N__50962\,
            I => \N__50853\
        );

    \I__11057\ : InMux
    port map (
            O => \N__50961\,
            I => \N__50853\
        );

    \I__11056\ : Sp12to4
    port map (
            O => \N__50956\,
            I => \N__50850\
        );

    \I__11055\ : InMux
    port map (
            O => \N__50955\,
            I => \N__50846\
        );

    \I__11054\ : InMux
    port map (
            O => \N__50954\,
            I => \N__50843\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__50951\,
            I => \N__50830\
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__50948\,
            I => \N__50830\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__50945\,
            I => \N__50830\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__50942\,
            I => \N__50830\
        );

    \I__11049\ : Span4Mux_v
    port map (
            O => \N__50937\,
            I => \N__50830\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__50930\,
            I => \N__50830\
        );

    \I__11047\ : InMux
    port map (
            O => \N__50929\,
            I => \N__50827\
        );

    \I__11046\ : Span12Mux_h
    port map (
            O => \N__50924\,
            I => \N__50823\
        );

    \I__11045\ : Span4Mux_h
    port map (
            O => \N__50919\,
            I => \N__50820\
        );

    \I__11044\ : Span4Mux_h
    port map (
            O => \N__50914\,
            I => \N__50813\
        );

    \I__11043\ : Span4Mux_v
    port map (
            O => \N__50911\,
            I => \N__50813\
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__50904\,
            I => \N__50813\
        );

    \I__11041\ : LocalMux
    port map (
            O => \N__50901\,
            I => \N__50810\
        );

    \I__11040\ : Span4Mux_v
    port map (
            O => \N__50888\,
            I => \N__50803\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__50883\,
            I => \N__50803\
        );

    \I__11038\ : Span4Mux_h
    port map (
            O => \N__50880\,
            I => \N__50803\
        );

    \I__11037\ : LocalMux
    port map (
            O => \N__50877\,
            I => \N__50791\
        );

    \I__11036\ : Sp12to4
    port map (
            O => \N__50874\,
            I => \N__50791\
        );

    \I__11035\ : LocalMux
    port map (
            O => \N__50871\,
            I => \N__50791\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__50866\,
            I => \N__50791\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__50861\,
            I => \N__50791\
        );

    \I__11032\ : Span12Mux_h
    port map (
            O => \N__50858\,
            I => \N__50784\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__50853\,
            I => \N__50784\
        );

    \I__11030\ : Span12Mux_s7_v
    port map (
            O => \N__50850\,
            I => \N__50784\
        );

    \I__11029\ : CascadeMux
    port map (
            O => \N__50849\,
            I => \N__50781\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__50846\,
            I => \N__50768\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__50843\,
            I => \N__50768\
        );

    \I__11026\ : Span4Mux_v
    port map (
            O => \N__50830\,
            I => \N__50768\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__50827\,
            I => \N__50768\
        );

    \I__11024\ : InMux
    port map (
            O => \N__50826\,
            I => \N__50765\
        );

    \I__11023\ : Span12Mux_v
    port map (
            O => \N__50823\,
            I => \N__50762\
        );

    \I__11022\ : Span4Mux_v
    port map (
            O => \N__50820\,
            I => \N__50757\
        );

    \I__11021\ : Span4Mux_v
    port map (
            O => \N__50813\,
            I => \N__50757\
        );

    \I__11020\ : Span4Mux_h
    port map (
            O => \N__50810\,
            I => \N__50752\
        );

    \I__11019\ : Span4Mux_h
    port map (
            O => \N__50803\,
            I => \N__50752\
        );

    \I__11018\ : InMux
    port map (
            O => \N__50802\,
            I => \N__50749\
        );

    \I__11017\ : Span12Mux_v
    port map (
            O => \N__50791\,
            I => \N__50744\
        );

    \I__11016\ : Span12Mux_v
    port map (
            O => \N__50784\,
            I => \N__50744\
        );

    \I__11015\ : InMux
    port map (
            O => \N__50781\,
            I => \N__50739\
        );

    \I__11014\ : InMux
    port map (
            O => \N__50780\,
            I => \N__50739\
        );

    \I__11013\ : InMux
    port map (
            O => \N__50779\,
            I => \N__50732\
        );

    \I__11012\ : InMux
    port map (
            O => \N__50778\,
            I => \N__50732\
        );

    \I__11011\ : InMux
    port map (
            O => \N__50777\,
            I => \N__50732\
        );

    \I__11010\ : Span4Mux_h
    port map (
            O => \N__50768\,
            I => \N__50729\
        );

    \I__11009\ : LocalMux
    port map (
            O => \N__50765\,
            I => \c0.n1220\
        );

    \I__11008\ : Odrv12
    port map (
            O => \N__50762\,
            I => \c0.n1220\
        );

    \I__11007\ : Odrv4
    port map (
            O => \N__50757\,
            I => \c0.n1220\
        );

    \I__11006\ : Odrv4
    port map (
            O => \N__50752\,
            I => \c0.n1220\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__50749\,
            I => \c0.n1220\
        );

    \I__11004\ : Odrv12
    port map (
            O => \N__50744\,
            I => \c0.n1220\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__50739\,
            I => \c0.n1220\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__50732\,
            I => \c0.n1220\
        );

    \I__11001\ : Odrv4
    port map (
            O => \N__50729\,
            I => \c0.n1220\
        );

    \I__11000\ : InMux
    port map (
            O => \N__50710\,
            I => \N__50706\
        );

    \I__10999\ : CascadeMux
    port map (
            O => \N__50709\,
            I => \N__50703\
        );

    \I__10998\ : LocalMux
    port map (
            O => \N__50706\,
            I => \N__50700\
        );

    \I__10997\ : InMux
    port map (
            O => \N__50703\,
            I => \N__50696\
        );

    \I__10996\ : Span4Mux_v
    port map (
            O => \N__50700\,
            I => \N__50693\
        );

    \I__10995\ : InMux
    port map (
            O => \N__50699\,
            I => \N__50690\
        );

    \I__10994\ : LocalMux
    port map (
            O => \N__50696\,
            I => \N__50685\
        );

    \I__10993\ : Span4Mux_v
    port map (
            O => \N__50693\,
            I => \N__50685\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__50690\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__10991\ : Odrv4
    port map (
            O => \N__50685\,
            I => \c0.FRAME_MATCHER_i_28\
        );

    \I__10990\ : InMux
    port map (
            O => \N__50680\,
            I => \N__50675\
        );

    \I__10989\ : CascadeMux
    port map (
            O => \N__50679\,
            I => \N__50670\
        );

    \I__10988\ : InMux
    port map (
            O => \N__50678\,
            I => \N__50655\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__50675\,
            I => \N__50652\
        );

    \I__10986\ : InMux
    port map (
            O => \N__50674\,
            I => \N__50643\
        );

    \I__10985\ : InMux
    port map (
            O => \N__50673\,
            I => \N__50640\
        );

    \I__10984\ : InMux
    port map (
            O => \N__50670\,
            I => \N__50637\
        );

    \I__10983\ : InMux
    port map (
            O => \N__50669\,
            I => \N__50632\
        );

    \I__10982\ : InMux
    port map (
            O => \N__50668\,
            I => \N__50632\
        );

    \I__10981\ : InMux
    port map (
            O => \N__50667\,
            I => \N__50629\
        );

    \I__10980\ : InMux
    port map (
            O => \N__50666\,
            I => \N__50622\
        );

    \I__10979\ : InMux
    port map (
            O => \N__50665\,
            I => \N__50622\
        );

    \I__10978\ : InMux
    port map (
            O => \N__50664\,
            I => \N__50622\
        );

    \I__10977\ : InMux
    port map (
            O => \N__50663\,
            I => \N__50617\
        );

    \I__10976\ : InMux
    port map (
            O => \N__50662\,
            I => \N__50612\
        );

    \I__10975\ : InMux
    port map (
            O => \N__50661\,
            I => \N__50612\
        );

    \I__10974\ : InMux
    port map (
            O => \N__50660\,
            I => \N__50606\
        );

    \I__10973\ : InMux
    port map (
            O => \N__50659\,
            I => \N__50601\
        );

    \I__10972\ : InMux
    port map (
            O => \N__50658\,
            I => \N__50601\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__50655\,
            I => \N__50596\
        );

    \I__10970\ : Span4Mux_v
    port map (
            O => \N__50652\,
            I => \N__50596\
        );

    \I__10969\ : InMux
    port map (
            O => \N__50651\,
            I => \N__50591\
        );

    \I__10968\ : InMux
    port map (
            O => \N__50650\,
            I => \N__50588\
        );

    \I__10967\ : InMux
    port map (
            O => \N__50649\,
            I => \N__50583\
        );

    \I__10966\ : InMux
    port map (
            O => \N__50648\,
            I => \N__50583\
        );

    \I__10965\ : InMux
    port map (
            O => \N__50647\,
            I => \N__50578\
        );

    \I__10964\ : InMux
    port map (
            O => \N__50646\,
            I => \N__50578\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__50643\,
            I => \N__50567\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__50640\,
            I => \N__50567\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__50637\,
            I => \N__50567\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__50632\,
            I => \N__50567\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__50629\,
            I => \N__50567\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__50622\,
            I => \N__50564\
        );

    \I__10957\ : InMux
    port map (
            O => \N__50621\,
            I => \N__50561\
        );

    \I__10956\ : InMux
    port map (
            O => \N__50620\,
            I => \N__50558\
        );

    \I__10955\ : LocalMux
    port map (
            O => \N__50617\,
            I => \N__50553\
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__50612\,
            I => \N__50553\
        );

    \I__10953\ : InMux
    port map (
            O => \N__50611\,
            I => \N__50546\
        );

    \I__10952\ : InMux
    port map (
            O => \N__50610\,
            I => \N__50546\
        );

    \I__10951\ : InMux
    port map (
            O => \N__50609\,
            I => \N__50546\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__50606\,
            I => \N__50541\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__50601\,
            I => \N__50541\
        );

    \I__10948\ : Span4Mux_h
    port map (
            O => \N__50596\,
            I => \N__50538\
        );

    \I__10947\ : InMux
    port map (
            O => \N__50595\,
            I => \N__50532\
        );

    \I__10946\ : InMux
    port map (
            O => \N__50594\,
            I => \N__50532\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__50591\,
            I => \N__50527\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__50588\,
            I => \N__50527\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__50583\,
            I => \N__50520\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__50578\,
            I => \N__50520\
        );

    \I__10941\ : Span4Mux_v
    port map (
            O => \N__50567\,
            I => \N__50520\
        );

    \I__10940\ : Span4Mux_h
    port map (
            O => \N__50564\,
            I => \N__50517\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__50561\,
            I => \N__50512\
        );

    \I__10938\ : LocalMux
    port map (
            O => \N__50558\,
            I => \N__50512\
        );

    \I__10937\ : Span12Mux_s7_v
    port map (
            O => \N__50553\,
            I => \N__50507\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__50546\,
            I => \N__50507\
        );

    \I__10935\ : Span4Mux_h
    port map (
            O => \N__50541\,
            I => \N__50504\
        );

    \I__10934\ : Span4Mux_v
    port map (
            O => \N__50538\,
            I => \N__50501\
        );

    \I__10933\ : InMux
    port map (
            O => \N__50537\,
            I => \N__50495\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__50532\,
            I => \N__50486\
        );

    \I__10931\ : Span4Mux_v
    port map (
            O => \N__50527\,
            I => \N__50486\
        );

    \I__10930\ : Span4Mux_v
    port map (
            O => \N__50520\,
            I => \N__50486\
        );

    \I__10929\ : Span4Mux_v
    port map (
            O => \N__50517\,
            I => \N__50486\
        );

    \I__10928\ : Span12Mux_v
    port map (
            O => \N__50512\,
            I => \N__50481\
        );

    \I__10927\ : Span12Mux_v
    port map (
            O => \N__50507\,
            I => \N__50481\
        );

    \I__10926\ : Span4Mux_v
    port map (
            O => \N__50504\,
            I => \N__50478\
        );

    \I__10925\ : Sp12to4
    port map (
            O => \N__50501\,
            I => \N__50475\
        );

    \I__10924\ : InMux
    port map (
            O => \N__50500\,
            I => \N__50468\
        );

    \I__10923\ : InMux
    port map (
            O => \N__50499\,
            I => \N__50468\
        );

    \I__10922\ : InMux
    port map (
            O => \N__50498\,
            I => \N__50468\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__50495\,
            I => \c0.n31_adj_4271\
        );

    \I__10920\ : Odrv4
    port map (
            O => \N__50486\,
            I => \c0.n31_adj_4271\
        );

    \I__10919\ : Odrv12
    port map (
            O => \N__50481\,
            I => \c0.n31_adj_4271\
        );

    \I__10918\ : Odrv4
    port map (
            O => \N__50478\,
            I => \c0.n31_adj_4271\
        );

    \I__10917\ : Odrv12
    port map (
            O => \N__50475\,
            I => \c0.n31_adj_4271\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__50468\,
            I => \c0.n31_adj_4271\
        );

    \I__10915\ : SRMux
    port map (
            O => \N__50455\,
            I => \N__50452\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__50452\,
            I => \N__50449\
        );

    \I__10913\ : Span4Mux_h
    port map (
            O => \N__50449\,
            I => \N__50446\
        );

    \I__10912\ : Odrv4
    port map (
            O => \N__50446\,
            I => \c0.n3_adj_4430\
        );

    \I__10911\ : InMux
    port map (
            O => \N__50443\,
            I => \N__50440\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__50440\,
            I => \N__50435\
        );

    \I__10909\ : InMux
    port map (
            O => \N__50439\,
            I => \N__50432\
        );

    \I__10908\ : InMux
    port map (
            O => \N__50438\,
            I => \N__50429\
        );

    \I__10907\ : Span4Mux_v
    port map (
            O => \N__50435\,
            I => \N__50426\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__50432\,
            I => \N__50423\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__50429\,
            I => \c0.data_in_frame_7_4\
        );

    \I__10904\ : Odrv4
    port map (
            O => \N__50426\,
            I => \c0.data_in_frame_7_4\
        );

    \I__10903\ : Odrv12
    port map (
            O => \N__50423\,
            I => \c0.data_in_frame_7_4\
        );

    \I__10902\ : CascadeMux
    port map (
            O => \N__50416\,
            I => \c0.n13555_cascade_\
        );

    \I__10901\ : InMux
    port map (
            O => \N__50413\,
            I => \N__50410\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__50410\,
            I => \N__50407\
        );

    \I__10899\ : Span4Mux_h
    port map (
            O => \N__50407\,
            I => \N__50404\
        );

    \I__10898\ : Span4Mux_v
    port map (
            O => \N__50404\,
            I => \N__50400\
        );

    \I__10897\ : InMux
    port map (
            O => \N__50403\,
            I => \N__50397\
        );

    \I__10896\ : Odrv4
    port map (
            O => \N__50400\,
            I => \c0.n13555\
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__50397\,
            I => \c0.n13555\
        );

    \I__10894\ : CascadeMux
    port map (
            O => \N__50392\,
            I => \c0.n22043_cascade_\
        );

    \I__10893\ : InMux
    port map (
            O => \N__50389\,
            I => \N__50385\
        );

    \I__10892\ : InMux
    port map (
            O => \N__50388\,
            I => \N__50382\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__50385\,
            I => \N__50378\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__50382\,
            I => \N__50375\
        );

    \I__10889\ : InMux
    port map (
            O => \N__50381\,
            I => \N__50372\
        );

    \I__10888\ : Span4Mux_h
    port map (
            O => \N__50378\,
            I => \N__50369\
        );

    \I__10887\ : Span4Mux_v
    port map (
            O => \N__50375\,
            I => \N__50365\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__50372\,
            I => \N__50360\
        );

    \I__10885\ : Span4Mux_v
    port map (
            O => \N__50369\,
            I => \N__50360\
        );

    \I__10884\ : InMux
    port map (
            O => \N__50368\,
            I => \N__50357\
        );

    \I__10883\ : Odrv4
    port map (
            O => \N__50365\,
            I => \c0.data_in_frame_2_6\
        );

    \I__10882\ : Odrv4
    port map (
            O => \N__50360\,
            I => \c0.data_in_frame_2_6\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__50357\,
            I => \c0.data_in_frame_2_6\
        );

    \I__10880\ : InMux
    port map (
            O => \N__50350\,
            I => \N__50346\
        );

    \I__10879\ : InMux
    port map (
            O => \N__50349\,
            I => \N__50342\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__50346\,
            I => \N__50336\
        );

    \I__10877\ : InMux
    port map (
            O => \N__50345\,
            I => \N__50333\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__50342\,
            I => \N__50330\
        );

    \I__10875\ : InMux
    port map (
            O => \N__50341\,
            I => \N__50325\
        );

    \I__10874\ : InMux
    port map (
            O => \N__50340\,
            I => \N__50325\
        );

    \I__10873\ : InMux
    port map (
            O => \N__50339\,
            I => \N__50322\
        );

    \I__10872\ : Span4Mux_h
    port map (
            O => \N__50336\,
            I => \N__50318\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__50333\,
            I => \N__50315\
        );

    \I__10870\ : Span4Mux_v
    port map (
            O => \N__50330\,
            I => \N__50308\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__50325\,
            I => \N__50308\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__50322\,
            I => \N__50308\
        );

    \I__10867\ : InMux
    port map (
            O => \N__50321\,
            I => \N__50303\
        );

    \I__10866\ : Span4Mux_v
    port map (
            O => \N__50318\,
            I => \N__50300\
        );

    \I__10865\ : Span4Mux_v
    port map (
            O => \N__50315\,
            I => \N__50295\
        );

    \I__10864\ : Span4Mux_h
    port map (
            O => \N__50308\,
            I => \N__50295\
        );

    \I__10863\ : InMux
    port map (
            O => \N__50307\,
            I => \N__50290\
        );

    \I__10862\ : InMux
    port map (
            O => \N__50306\,
            I => \N__50290\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__50303\,
            I => \c0.data_in_frame_0_4\
        );

    \I__10860\ : Odrv4
    port map (
            O => \N__50300\,
            I => \c0.data_in_frame_0_4\
        );

    \I__10859\ : Odrv4
    port map (
            O => \N__50295\,
            I => \c0.data_in_frame_0_4\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__50290\,
            I => \c0.data_in_frame_0_4\
        );

    \I__10857\ : CascadeMux
    port map (
            O => \N__50281\,
            I => \N__50278\
        );

    \I__10856\ : InMux
    port map (
            O => \N__50278\,
            I => \N__50275\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__50275\,
            I => \N__50272\
        );

    \I__10854\ : Odrv12
    port map (
            O => \N__50272\,
            I => \c0.n10_adj_4363\
        );

    \I__10853\ : CascadeMux
    port map (
            O => \N__50269\,
            I => \c0.rx.n22573_cascade_\
        );

    \I__10852\ : CascadeMux
    port map (
            O => \N__50266\,
            I => \c0.rx.n12_cascade_\
        );

    \I__10851\ : InMux
    port map (
            O => \N__50263\,
            I => \bfn_20_24_0_\
        );

    \I__10850\ : InMux
    port map (
            O => \N__50260\,
            I => \N__50256\
        );

    \I__10849\ : InMux
    port map (
            O => \N__50259\,
            I => \N__50253\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__50256\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__50253\,
            I => \c0.rx.r_Clock_Count_1\
        );

    \I__10846\ : InMux
    port map (
            O => \N__50248\,
            I => \c0.rx.n19533\
        );

    \I__10845\ : InMux
    port map (
            O => \N__50245\,
            I => \N__50241\
        );

    \I__10844\ : InMux
    port map (
            O => \N__50244\,
            I => \N__50238\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__50241\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__50238\,
            I => \c0.rx.r_Clock_Count_2\
        );

    \I__10841\ : InMux
    port map (
            O => \N__50233\,
            I => \c0.rx.n19534\
        );

    \I__10840\ : InMux
    port map (
            O => \N__50230\,
            I => \N__50226\
        );

    \I__10839\ : InMux
    port map (
            O => \N__50229\,
            I => \N__50223\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__50226\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__50223\,
            I => \c0.rx.r_Clock_Count_3\
        );

    \I__10836\ : InMux
    port map (
            O => \N__50218\,
            I => \c0.rx.n19535\
        );

    \I__10835\ : InMux
    port map (
            O => \N__50215\,
            I => \c0.rx.n19536\
        );

    \I__10834\ : InMux
    port map (
            O => \N__50212\,
            I => \c0.rx.n19537\
        );

    \I__10833\ : InMux
    port map (
            O => \N__50209\,
            I => \c0.rx.n19538\
        );

    \I__10832\ : InMux
    port map (
            O => \N__50206\,
            I => \N__50201\
        );

    \I__10831\ : InMux
    port map (
            O => \N__50205\,
            I => \N__50198\
        );

    \I__10830\ : InMux
    port map (
            O => \N__50204\,
            I => \N__50195\
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__50201\,
            I => \N__50192\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__50198\,
            I => \N__50186\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__50195\,
            I => \N__50186\
        );

    \I__10826\ : Span4Mux_h
    port map (
            O => \N__50192\,
            I => \N__50183\
        );

    \I__10825\ : InMux
    port map (
            O => \N__50191\,
            I => \N__50180\
        );

    \I__10824\ : Span4Mux_h
    port map (
            O => \N__50186\,
            I => \N__50177\
        );

    \I__10823\ : Span4Mux_v
    port map (
            O => \N__50183\,
            I => \N__50174\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__50180\,
            I => \c0.data_in_frame_27_1\
        );

    \I__10821\ : Odrv4
    port map (
            O => \N__50177\,
            I => \c0.data_in_frame_27_1\
        );

    \I__10820\ : Odrv4
    port map (
            O => \N__50174\,
            I => \c0.data_in_frame_27_1\
        );

    \I__10819\ : CascadeMux
    port map (
            O => \N__50167\,
            I => \N__50164\
        );

    \I__10818\ : InMux
    port map (
            O => \N__50164\,
            I => \N__50161\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__50161\,
            I => \N__50158\
        );

    \I__10816\ : Span4Mux_v
    port map (
            O => \N__50158\,
            I => \N__50154\
        );

    \I__10815\ : InMux
    port map (
            O => \N__50157\,
            I => \N__50151\
        );

    \I__10814\ : Span4Mux_v
    port map (
            O => \N__50154\,
            I => \N__50148\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__50151\,
            I => \N__50145\
        );

    \I__10812\ : Span4Mux_v
    port map (
            O => \N__50148\,
            I => \N__50142\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__50145\,
            I => \N__50139\
        );

    \I__10810\ : Span4Mux_v
    port map (
            O => \N__50142\,
            I => \N__50135\
        );

    \I__10809\ : Span4Mux_v
    port map (
            O => \N__50139\,
            I => \N__50132\
        );

    \I__10808\ : InMux
    port map (
            O => \N__50138\,
            I => \N__50129\
        );

    \I__10807\ : Odrv4
    port map (
            O => \N__50135\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__10806\ : Odrv4
    port map (
            O => \N__50132\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__50129\,
            I => \c0.FRAME_MATCHER_i_10\
        );

    \I__10804\ : SRMux
    port map (
            O => \N__50122\,
            I => \N__50119\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__50119\,
            I => \N__50116\
        );

    \I__10802\ : Span4Mux_v
    port map (
            O => \N__50116\,
            I => \N__50113\
        );

    \I__10801\ : Sp12to4
    port map (
            O => \N__50113\,
            I => \N__50110\
        );

    \I__10800\ : Odrv12
    port map (
            O => \N__50110\,
            I => \c0.n3_adj_4460\
        );

    \I__10799\ : InMux
    port map (
            O => \N__50107\,
            I => \N__50103\
        );

    \I__10798\ : InMux
    port map (
            O => \N__50106\,
            I => \N__50100\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__50103\,
            I => \N__50097\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__50100\,
            I => \N__50094\
        );

    \I__10795\ : Span4Mux_v
    port map (
            O => \N__50097\,
            I => \N__50091\
        );

    \I__10794\ : Span12Mux_h
    port map (
            O => \N__50094\,
            I => \N__50088\
        );

    \I__10793\ : Span4Mux_v
    port map (
            O => \N__50091\,
            I => \N__50085\
        );

    \I__10792\ : Odrv12
    port map (
            O => \N__50088\,
            I => n18678
        );

    \I__10791\ : Odrv4
    port map (
            O => \N__50085\,
            I => n18678
        );

    \I__10790\ : CascadeMux
    port map (
            O => \N__50080\,
            I => \c0.rx.n18655_cascade_\
        );

    \I__10789\ : CascadeMux
    port map (
            O => \N__50077\,
            I => \c0.rx.n21704_cascade_\
        );

    \I__10788\ : InMux
    port map (
            O => \N__50074\,
            I => \N__50065\
        );

    \I__10787\ : InMux
    port map (
            O => \N__50073\,
            I => \N__50065\
        );

    \I__10786\ : InMux
    port map (
            O => \N__50072\,
            I => \N__50065\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__50065\,
            I => \c0.data_in_frame_23_4\
        );

    \I__10784\ : CascadeMux
    port map (
            O => \N__50062\,
            I => \c0.n10_adj_4287_cascade_\
        );

    \I__10783\ : InMux
    port map (
            O => \N__50059\,
            I => \N__50056\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__50056\,
            I => \N__50053\
        );

    \I__10781\ : Span4Mux_h
    port map (
            O => \N__50053\,
            I => \N__50050\
        );

    \I__10780\ : Odrv4
    port map (
            O => \N__50050\,
            I => \c0.n22_adj_4298\
        );

    \I__10779\ : InMux
    port map (
            O => \N__50047\,
            I => \N__50044\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__50044\,
            I => \N__50041\
        );

    \I__10777\ : Odrv4
    port map (
            O => \N__50041\,
            I => \c0.n13266\
        );

    \I__10776\ : InMux
    port map (
            O => \N__50038\,
            I => \N__50035\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__50035\,
            I => \N__50031\
        );

    \I__10774\ : InMux
    port map (
            O => \N__50034\,
            I => \N__50028\
        );

    \I__10773\ : Span4Mux_h
    port map (
            O => \N__50031\,
            I => \N__50025\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__50028\,
            I => \c0.data_in_frame_29_7\
        );

    \I__10771\ : Odrv4
    port map (
            O => \N__50025\,
            I => \c0.data_in_frame_29_7\
        );

    \I__10770\ : CascadeMux
    port map (
            O => \N__50020\,
            I => \c0.n21233_cascade_\
        );

    \I__10769\ : InMux
    port map (
            O => \N__50017\,
            I => \N__50014\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__50014\,
            I => \c0.n23506\
        );

    \I__10767\ : CascadeMux
    port map (
            O => \N__50011\,
            I => \N__50007\
        );

    \I__10766\ : CascadeMux
    port map (
            O => \N__50010\,
            I => \N__50004\
        );

    \I__10765\ : InMux
    port map (
            O => \N__50007\,
            I => \N__50001\
        );

    \I__10764\ : InMux
    port map (
            O => \N__50004\,
            I => \N__49998\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__50001\,
            I => \N__49993\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__49998\,
            I => \N__49993\
        );

    \I__10761\ : Span4Mux_h
    port map (
            O => \N__49993\,
            I => \N__49989\
        );

    \I__10760\ : InMux
    port map (
            O => \N__49992\,
            I => \N__49986\
        );

    \I__10759\ : Odrv4
    port map (
            O => \N__49989\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__49986\,
            I => \c0.FRAME_MATCHER_i_20\
        );

    \I__10757\ : SRMux
    port map (
            O => \N__49981\,
            I => \N__49978\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__49978\,
            I => \N__49975\
        );

    \I__10755\ : Span4Mux_v
    port map (
            O => \N__49975\,
            I => \N__49972\
        );

    \I__10754\ : Odrv4
    port map (
            O => \N__49972\,
            I => \c0.n3_adj_4442\
        );

    \I__10753\ : CascadeMux
    port map (
            O => \N__49969\,
            I => \N__49966\
        );

    \I__10752\ : InMux
    port map (
            O => \N__49966\,
            I => \N__49963\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__49963\,
            I => \N__49959\
        );

    \I__10750\ : CascadeMux
    port map (
            O => \N__49962\,
            I => \N__49956\
        );

    \I__10749\ : Span4Mux_h
    port map (
            O => \N__49959\,
            I => \N__49953\
        );

    \I__10748\ : InMux
    port map (
            O => \N__49956\,
            I => \N__49950\
        );

    \I__10747\ : Span4Mux_h
    port map (
            O => \N__49953\,
            I => \N__49947\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__49950\,
            I => \c0.data_in_frame_28_1\
        );

    \I__10745\ : Odrv4
    port map (
            O => \N__49947\,
            I => \c0.data_in_frame_28_1\
        );

    \I__10744\ : CascadeMux
    port map (
            O => \N__49942\,
            I => \c0.n21870_cascade_\
        );

    \I__10743\ : CascadeMux
    port map (
            O => \N__49939\,
            I => \N__49936\
        );

    \I__10742\ : InMux
    port map (
            O => \N__49936\,
            I => \N__49931\
        );

    \I__10741\ : InMux
    port map (
            O => \N__49935\,
            I => \N__49926\
        );

    \I__10740\ : InMux
    port map (
            O => \N__49934\,
            I => \N__49926\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__49931\,
            I => \c0.data_in_frame_21_3\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__49926\,
            I => \c0.data_in_frame_21_3\
        );

    \I__10737\ : InMux
    port map (
            O => \N__49921\,
            I => \N__49916\
        );

    \I__10736\ : InMux
    port map (
            O => \N__49920\,
            I => \N__49913\
        );

    \I__10735\ : InMux
    port map (
            O => \N__49919\,
            I => \N__49910\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__49916\,
            I => \N__49905\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__49913\,
            I => \N__49905\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__49910\,
            I => \c0.data_in_frame_23_5\
        );

    \I__10731\ : Odrv4
    port map (
            O => \N__49905\,
            I => \c0.data_in_frame_23_5\
        );

    \I__10730\ : CascadeMux
    port map (
            O => \N__49900\,
            I => \c0.n21858_cascade_\
        );

    \I__10729\ : CascadeMux
    port map (
            O => \N__49897\,
            I => \N__49894\
        );

    \I__10728\ : InMux
    port map (
            O => \N__49894\,
            I => \N__49891\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__49891\,
            I => \N__49886\
        );

    \I__10726\ : InMux
    port map (
            O => \N__49890\,
            I => \N__49883\
        );

    \I__10725\ : InMux
    port map (
            O => \N__49889\,
            I => \N__49880\
        );

    \I__10724\ : Odrv4
    port map (
            O => \N__49886\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__49883\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__49880\,
            I => \c0.FRAME_MATCHER_i_16\
        );

    \I__10721\ : InMux
    port map (
            O => \N__49873\,
            I => \N__49870\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__49870\,
            I => \N__49867\
        );

    \I__10719\ : Span4Mux_v
    port map (
            O => \N__49867\,
            I => \N__49864\
        );

    \I__10718\ : Odrv4
    port map (
            O => \N__49864\,
            I => \c0.n16_adj_4375\
        );

    \I__10717\ : CascadeMux
    port map (
            O => \N__49861\,
            I => \N__49858\
        );

    \I__10716\ : InMux
    port map (
            O => \N__49858\,
            I => \N__49852\
        );

    \I__10715\ : InMux
    port map (
            O => \N__49857\,
            I => \N__49852\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__49852\,
            I => \N__49848\
        );

    \I__10713\ : InMux
    port map (
            O => \N__49851\,
            I => \N__49845\
        );

    \I__10712\ : Span4Mux_v
    port map (
            O => \N__49848\,
            I => \N__49842\
        );

    \I__10711\ : LocalMux
    port map (
            O => \N__49845\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__10710\ : Odrv4
    port map (
            O => \N__49842\,
            I => \c0.FRAME_MATCHER_i_13\
        );

    \I__10709\ : SRMux
    port map (
            O => \N__49837\,
            I => \N__49834\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__49834\,
            I => \N__49831\
        );

    \I__10707\ : Span4Mux_h
    port map (
            O => \N__49831\,
            I => \N__49828\
        );

    \I__10706\ : Span4Mux_h
    port map (
            O => \N__49828\,
            I => \N__49825\
        );

    \I__10705\ : Odrv4
    port map (
            O => \N__49825\,
            I => \c0.n3_adj_4454\
        );

    \I__10704\ : InMux
    port map (
            O => \N__49822\,
            I => \N__49818\
        );

    \I__10703\ : InMux
    port map (
            O => \N__49821\,
            I => \N__49815\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__49818\,
            I => \N__49811\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__49815\,
            I => \N__49808\
        );

    \I__10700\ : InMux
    port map (
            O => \N__49814\,
            I => \N__49805\
        );

    \I__10699\ : Span4Mux_v
    port map (
            O => \N__49811\,
            I => \N__49802\
        );

    \I__10698\ : Odrv4
    port map (
            O => \N__49808\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__49805\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__10696\ : Odrv4
    port map (
            O => \N__49802\,
            I => \c0.FRAME_MATCHER_i_15\
        );

    \I__10695\ : SRMux
    port map (
            O => \N__49795\,
            I => \N__49792\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__49792\,
            I => \N__49789\
        );

    \I__10693\ : Span4Mux_h
    port map (
            O => \N__49789\,
            I => \N__49786\
        );

    \I__10692\ : Odrv4
    port map (
            O => \N__49786\,
            I => \c0.n3_adj_4452\
        );

    \I__10691\ : InMux
    port map (
            O => \N__49783\,
            I => \N__49780\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__49780\,
            I => \N__49776\
        );

    \I__10689\ : InMux
    port map (
            O => \N__49779\,
            I => \N__49773\
        );

    \I__10688\ : Span4Mux_v
    port map (
            O => \N__49776\,
            I => \N__49768\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__49773\,
            I => \N__49768\
        );

    \I__10686\ : Span4Mux_v
    port map (
            O => \N__49768\,
            I => \N__49765\
        );

    \I__10685\ : Odrv4
    port map (
            O => \N__49765\,
            I => \c0.n13697\
        );

    \I__10684\ : CascadeMux
    port map (
            O => \N__49762\,
            I => \c0.n22440_cascade_\
        );

    \I__10683\ : InMux
    port map (
            O => \N__49759\,
            I => \N__49756\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__49756\,
            I => \N__49750\
        );

    \I__10681\ : InMux
    port map (
            O => \N__49755\,
            I => \N__49745\
        );

    \I__10680\ : InMux
    port map (
            O => \N__49754\,
            I => \N__49745\
        );

    \I__10679\ : CascadeMux
    port map (
            O => \N__49753\,
            I => \N__49742\
        );

    \I__10678\ : Span4Mux_v
    port map (
            O => \N__49750\,
            I => \N__49737\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__49745\,
            I => \N__49737\
        );

    \I__10676\ : InMux
    port map (
            O => \N__49742\,
            I => \N__49733\
        );

    \I__10675\ : Span4Mux_v
    port map (
            O => \N__49737\,
            I => \N__49730\
        );

    \I__10674\ : InMux
    port map (
            O => \N__49736\,
            I => \N__49727\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__49733\,
            I => \c0.data_in_frame_10_7\
        );

    \I__10672\ : Odrv4
    port map (
            O => \N__49730\,
            I => \c0.data_in_frame_10_7\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__49727\,
            I => \c0.data_in_frame_10_7\
        );

    \I__10670\ : CascadeMux
    port map (
            O => \N__49720\,
            I => \c0.n10_adj_4229_cascade_\
        );

    \I__10669\ : CascadeMux
    port map (
            O => \N__49717\,
            I => \c0.n5943_cascade_\
        );

    \I__10668\ : CascadeMux
    port map (
            O => \N__49714\,
            I => \c0.n22081_cascade_\
        );

    \I__10667\ : CascadeMux
    port map (
            O => \N__49711\,
            I => \c0.n22349_cascade_\
        );

    \I__10666\ : InMux
    port map (
            O => \N__49708\,
            I => \N__49704\
        );

    \I__10665\ : InMux
    port map (
            O => \N__49707\,
            I => \N__49700\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__49704\,
            I => \N__49697\
        );

    \I__10663\ : InMux
    port map (
            O => \N__49703\,
            I => \N__49694\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__49700\,
            I => \N__49688\
        );

    \I__10661\ : Span4Mux_v
    port map (
            O => \N__49697\,
            I => \N__49683\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__49694\,
            I => \N__49683\
        );

    \I__10659\ : InMux
    port map (
            O => \N__49693\,
            I => \N__49680\
        );

    \I__10658\ : InMux
    port map (
            O => \N__49692\,
            I => \N__49675\
        );

    \I__10657\ : InMux
    port map (
            O => \N__49691\,
            I => \N__49675\
        );

    \I__10656\ : Span4Mux_v
    port map (
            O => \N__49688\,
            I => \N__49669\
        );

    \I__10655\ : Span4Mux_h
    port map (
            O => \N__49683\,
            I => \N__49669\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__49680\,
            I => \N__49664\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__49675\,
            I => \N__49664\
        );

    \I__10652\ : InMux
    port map (
            O => \N__49674\,
            I => \N__49661\
        );

    \I__10651\ : Odrv4
    port map (
            O => \N__49669\,
            I => n21744
        );

    \I__10650\ : Odrv12
    port map (
            O => \N__49664\,
            I => n21744
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__49661\,
            I => n21744
        );

    \I__10648\ : InMux
    port map (
            O => \N__49654\,
            I => \N__49651\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__49651\,
            I => \N__49648\
        );

    \I__10646\ : Span4Mux_h
    port map (
            O => \N__49648\,
            I => \N__49645\
        );

    \I__10645\ : Odrv4
    port map (
            O => \N__49645\,
            I => \c0.n6_adj_4386\
        );

    \I__10644\ : CascadeMux
    port map (
            O => \N__49642\,
            I => \N__49638\
        );

    \I__10643\ : InMux
    port map (
            O => \N__49641\,
            I => \N__49635\
        );

    \I__10642\ : InMux
    port map (
            O => \N__49638\,
            I => \N__49631\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__49635\,
            I => \N__49628\
        );

    \I__10640\ : InMux
    port map (
            O => \N__49634\,
            I => \N__49625\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__49631\,
            I => \N__49622\
        );

    \I__10638\ : Span4Mux_h
    port map (
            O => \N__49628\,
            I => \N__49619\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__49625\,
            I => \N__49616\
        );

    \I__10636\ : Odrv12
    port map (
            O => \N__49622\,
            I => \c0.data_in_frame_4_3\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__49619\,
            I => \c0.data_in_frame_4_3\
        );

    \I__10634\ : Odrv12
    port map (
            O => \N__49616\,
            I => \c0.data_in_frame_4_3\
        );

    \I__10633\ : CascadeMux
    port map (
            O => \N__49609\,
            I => \N__49605\
        );

    \I__10632\ : InMux
    port map (
            O => \N__49608\,
            I => \N__49600\
        );

    \I__10631\ : InMux
    port map (
            O => \N__49605\,
            I => \N__49600\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__49600\,
            I => data_in_frame_6_4
        );

    \I__10629\ : InMux
    port map (
            O => \N__49597\,
            I => \N__49593\
        );

    \I__10628\ : CascadeMux
    port map (
            O => \N__49596\,
            I => \N__49590\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__49593\,
            I => \N__49586\
        );

    \I__10626\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49581\
        );

    \I__10625\ : InMux
    port map (
            O => \N__49589\,
            I => \N__49581\
        );

    \I__10624\ : Span4Mux_h
    port map (
            O => \N__49586\,
            I => \N__49578\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__49581\,
            I => \N__49573\
        );

    \I__10622\ : Span4Mux_v
    port map (
            O => \N__49578\,
            I => \N__49573\
        );

    \I__10621\ : Odrv4
    port map (
            O => \N__49573\,
            I => \c0.data_in_frame_4_2\
        );

    \I__10620\ : InMux
    port map (
            O => \N__49570\,
            I => \N__49566\
        );

    \I__10619\ : InMux
    port map (
            O => \N__49569\,
            I => \N__49562\
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__49566\,
            I => \N__49558\
        );

    \I__10617\ : InMux
    port map (
            O => \N__49565\,
            I => \N__49555\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__49562\,
            I => \N__49545\
        );

    \I__10615\ : InMux
    port map (
            O => \N__49561\,
            I => \N__49542\
        );

    \I__10614\ : Span4Mux_h
    port map (
            O => \N__49558\,
            I => \N__49539\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__49555\,
            I => \N__49536\
        );

    \I__10612\ : InMux
    port map (
            O => \N__49554\,
            I => \N__49531\
        );

    \I__10611\ : InMux
    port map (
            O => \N__49553\,
            I => \N__49531\
        );

    \I__10610\ : CascadeMux
    port map (
            O => \N__49552\,
            I => \N__49528\
        );

    \I__10609\ : CascadeMux
    port map (
            O => \N__49551\,
            I => \N__49525\
        );

    \I__10608\ : InMux
    port map (
            O => \N__49550\,
            I => \N__49520\
        );

    \I__10607\ : InMux
    port map (
            O => \N__49549\,
            I => \N__49520\
        );

    \I__10606\ : InMux
    port map (
            O => \N__49548\,
            I => \N__49514\
        );

    \I__10605\ : Span4Mux_v
    port map (
            O => \N__49545\,
            I => \N__49501\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__49542\,
            I => \N__49501\
        );

    \I__10603\ : Span4Mux_h
    port map (
            O => \N__49539\,
            I => \N__49501\
        );

    \I__10602\ : Span4Mux_h
    port map (
            O => \N__49536\,
            I => \N__49501\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__49531\,
            I => \N__49501\
        );

    \I__10600\ : InMux
    port map (
            O => \N__49528\,
            I => \N__49496\
        );

    \I__10599\ : InMux
    port map (
            O => \N__49525\,
            I => \N__49496\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__49520\,
            I => \N__49493\
        );

    \I__10597\ : InMux
    port map (
            O => \N__49519\,
            I => \N__49488\
        );

    \I__10596\ : InMux
    port map (
            O => \N__49518\,
            I => \N__49488\
        );

    \I__10595\ : InMux
    port map (
            O => \N__49517\,
            I => \N__49485\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__49514\,
            I => \N__49482\
        );

    \I__10593\ : InMux
    port map (
            O => \N__49513\,
            I => \N__49477\
        );

    \I__10592\ : InMux
    port map (
            O => \N__49512\,
            I => \N__49477\
        );

    \I__10591\ : Span4Mux_v
    port map (
            O => \N__49501\,
            I => \N__49457\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__49496\,
            I => \N__49457\
        );

    \I__10589\ : Span4Mux_h
    port map (
            O => \N__49493\,
            I => \N__49457\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__49488\,
            I => \N__49457\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__49485\,
            I => \N__49457\
        );

    \I__10586\ : Span4Mux_h
    port map (
            O => \N__49482\,
            I => \N__49457\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__49477\,
            I => \N__49457\
        );

    \I__10584\ : InMux
    port map (
            O => \N__49476\,
            I => \N__49438\
        );

    \I__10583\ : InMux
    port map (
            O => \N__49475\,
            I => \N__49438\
        );

    \I__10582\ : InMux
    port map (
            O => \N__49474\,
            I => \N__49431\
        );

    \I__10581\ : InMux
    port map (
            O => \N__49473\,
            I => \N__49431\
        );

    \I__10580\ : InMux
    port map (
            O => \N__49472\,
            I => \N__49431\
        );

    \I__10579\ : Span4Mux_v
    port map (
            O => \N__49457\,
            I => \N__49428\
        );

    \I__10578\ : InMux
    port map (
            O => \N__49456\,
            I => \N__49416\
        );

    \I__10577\ : InMux
    port map (
            O => \N__49455\,
            I => \N__49416\
        );

    \I__10576\ : InMux
    port map (
            O => \N__49454\,
            I => \N__49416\
        );

    \I__10575\ : InMux
    port map (
            O => \N__49453\,
            I => \N__49416\
        );

    \I__10574\ : CascadeMux
    port map (
            O => \N__49452\,
            I => \N__49407\
        );

    \I__10573\ : CascadeMux
    port map (
            O => \N__49451\,
            I => \N__49404\
        );

    \I__10572\ : InMux
    port map (
            O => \N__49450\,
            I => \N__49397\
        );

    \I__10571\ : InMux
    port map (
            O => \N__49449\,
            I => \N__49397\
        );

    \I__10570\ : InMux
    port map (
            O => \N__49448\,
            I => \N__49394\
        );

    \I__10569\ : InMux
    port map (
            O => \N__49447\,
            I => \N__49386\
        );

    \I__10568\ : InMux
    port map (
            O => \N__49446\,
            I => \N__49386\
        );

    \I__10567\ : InMux
    port map (
            O => \N__49445\,
            I => \N__49383\
        );

    \I__10566\ : InMux
    port map (
            O => \N__49444\,
            I => \N__49374\
        );

    \I__10565\ : InMux
    port map (
            O => \N__49443\,
            I => \N__49374\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__49438\,
            I => \N__49371\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__49431\,
            I => \N__49366\
        );

    \I__10562\ : Span4Mux_h
    port map (
            O => \N__49428\,
            I => \N__49366\
        );

    \I__10561\ : InMux
    port map (
            O => \N__49427\,
            I => \N__49359\
        );

    \I__10560\ : InMux
    port map (
            O => \N__49426\,
            I => \N__49359\
        );

    \I__10559\ : InMux
    port map (
            O => \N__49425\,
            I => \N__49359\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__49416\,
            I => \N__49353\
        );

    \I__10557\ : InMux
    port map (
            O => \N__49415\,
            I => \N__49348\
        );

    \I__10556\ : InMux
    port map (
            O => \N__49414\,
            I => \N__49348\
        );

    \I__10555\ : InMux
    port map (
            O => \N__49413\,
            I => \N__49345\
        );

    \I__10554\ : InMux
    port map (
            O => \N__49412\,
            I => \N__49340\
        );

    \I__10553\ : InMux
    port map (
            O => \N__49411\,
            I => \N__49340\
        );

    \I__10552\ : InMux
    port map (
            O => \N__49410\,
            I => \N__49337\
        );

    \I__10551\ : InMux
    port map (
            O => \N__49407\,
            I => \N__49326\
        );

    \I__10550\ : InMux
    port map (
            O => \N__49404\,
            I => \N__49326\
        );

    \I__10549\ : InMux
    port map (
            O => \N__49403\,
            I => \N__49323\
        );

    \I__10548\ : InMux
    port map (
            O => \N__49402\,
            I => \N__49317\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__49397\,
            I => \N__49314\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__49394\,
            I => \N__49311\
        );

    \I__10545\ : InMux
    port map (
            O => \N__49393\,
            I => \N__49304\
        );

    \I__10544\ : InMux
    port map (
            O => \N__49392\,
            I => \N__49304\
        );

    \I__10543\ : InMux
    port map (
            O => \N__49391\,
            I => \N__49304\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__49386\,
            I => \N__49299\
        );

    \I__10541\ : LocalMux
    port map (
            O => \N__49383\,
            I => \N__49299\
        );

    \I__10540\ : InMux
    port map (
            O => \N__49382\,
            I => \N__49292\
        );

    \I__10539\ : InMux
    port map (
            O => \N__49381\,
            I => \N__49292\
        );

    \I__10538\ : InMux
    port map (
            O => \N__49380\,
            I => \N__49292\
        );

    \I__10537\ : InMux
    port map (
            O => \N__49379\,
            I => \N__49289\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__49374\,
            I => \N__49280\
        );

    \I__10535\ : Span4Mux_h
    port map (
            O => \N__49371\,
            I => \N__49280\
        );

    \I__10534\ : Span4Mux_h
    port map (
            O => \N__49366\,
            I => \N__49280\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__49359\,
            I => \N__49280\
        );

    \I__10532\ : InMux
    port map (
            O => \N__49358\,
            I => \N__49275\
        );

    \I__10531\ : InMux
    port map (
            O => \N__49357\,
            I => \N__49275\
        );

    \I__10530\ : InMux
    port map (
            O => \N__49356\,
            I => \N__49266\
        );

    \I__10529\ : Span4Mux_h
    port map (
            O => \N__49353\,
            I => \N__49261\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__49348\,
            I => \N__49261\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__49345\,
            I => \N__49256\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__49340\,
            I => \N__49256\
        );

    \I__10525\ : LocalMux
    port map (
            O => \N__49337\,
            I => \N__49250\
        );

    \I__10524\ : InMux
    port map (
            O => \N__49336\,
            I => \N__49243\
        );

    \I__10523\ : InMux
    port map (
            O => \N__49335\,
            I => \N__49243\
        );

    \I__10522\ : InMux
    port map (
            O => \N__49334\,
            I => \N__49243\
        );

    \I__10521\ : InMux
    port map (
            O => \N__49333\,
            I => \N__49236\
        );

    \I__10520\ : InMux
    port map (
            O => \N__49332\,
            I => \N__49236\
        );

    \I__10519\ : InMux
    port map (
            O => \N__49331\,
            I => \N__49236\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__49326\,
            I => \N__49231\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__49323\,
            I => \N__49231\
        );

    \I__10516\ : InMux
    port map (
            O => \N__49322\,
            I => \N__49228\
        );

    \I__10515\ : InMux
    port map (
            O => \N__49321\,
            I => \N__49223\
        );

    \I__10514\ : InMux
    port map (
            O => \N__49320\,
            I => \N__49223\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__49317\,
            I => \N__49212\
        );

    \I__10512\ : Span4Mux_h
    port map (
            O => \N__49314\,
            I => \N__49212\
        );

    \I__10511\ : Span4Mux_h
    port map (
            O => \N__49311\,
            I => \N__49212\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__49304\,
            I => \N__49212\
        );

    \I__10509\ : Span4Mux_h
    port map (
            O => \N__49299\,
            I => \N__49212\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__49292\,
            I => \N__49207\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__49289\,
            I => \N__49207\
        );

    \I__10506\ : Span4Mux_v
    port map (
            O => \N__49280\,
            I => \N__49204\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__49275\,
            I => \N__49198\
        );

    \I__10504\ : InMux
    port map (
            O => \N__49274\,
            I => \N__49193\
        );

    \I__10503\ : InMux
    port map (
            O => \N__49273\,
            I => \N__49193\
        );

    \I__10502\ : InMux
    port map (
            O => \N__49272\,
            I => \N__49190\
        );

    \I__10501\ : InMux
    port map (
            O => \N__49271\,
            I => \N__49183\
        );

    \I__10500\ : InMux
    port map (
            O => \N__49270\,
            I => \N__49183\
        );

    \I__10499\ : InMux
    port map (
            O => \N__49269\,
            I => \N__49183\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__49266\,
            I => \N__49180\
        );

    \I__10497\ : Span4Mux_h
    port map (
            O => \N__49261\,
            I => \N__49176\
        );

    \I__10496\ : Span4Mux_h
    port map (
            O => \N__49256\,
            I => \N__49173\
        );

    \I__10495\ : InMux
    port map (
            O => \N__49255\,
            I => \N__49166\
        );

    \I__10494\ : InMux
    port map (
            O => \N__49254\,
            I => \N__49166\
        );

    \I__10493\ : InMux
    port map (
            O => \N__49253\,
            I => \N__49166\
        );

    \I__10492\ : Span4Mux_h
    port map (
            O => \N__49250\,
            I => \N__49161\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__49243\,
            I => \N__49161\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__49236\,
            I => \N__49156\
        );

    \I__10489\ : Span4Mux_v
    port map (
            O => \N__49231\,
            I => \N__49156\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__49228\,
            I => \N__49153\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__49223\,
            I => \N__49150\
        );

    \I__10486\ : Span4Mux_v
    port map (
            O => \N__49212\,
            I => \N__49145\
        );

    \I__10485\ : Span4Mux_h
    port map (
            O => \N__49207\,
            I => \N__49145\
        );

    \I__10484\ : Sp12to4
    port map (
            O => \N__49204\,
            I => \N__49141\
        );

    \I__10483\ : InMux
    port map (
            O => \N__49203\,
            I => \N__49136\
        );

    \I__10482\ : InMux
    port map (
            O => \N__49202\,
            I => \N__49136\
        );

    \I__10481\ : InMux
    port map (
            O => \N__49201\,
            I => \N__49133\
        );

    \I__10480\ : Span4Mux_v
    port map (
            O => \N__49198\,
            I => \N__49130\
        );

    \I__10479\ : LocalMux
    port map (
            O => \N__49193\,
            I => \N__49125\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__49190\,
            I => \N__49125\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__49183\,
            I => \N__49122\
        );

    \I__10476\ : Span4Mux_h
    port map (
            O => \N__49180\,
            I => \N__49119\
        );

    \I__10475\ : InMux
    port map (
            O => \N__49179\,
            I => \N__49116\
        );

    \I__10474\ : Sp12to4
    port map (
            O => \N__49176\,
            I => \N__49111\
        );

    \I__10473\ : Sp12to4
    port map (
            O => \N__49173\,
            I => \N__49111\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__49166\,
            I => \N__49104\
        );

    \I__10471\ : Span4Mux_v
    port map (
            O => \N__49161\,
            I => \N__49104\
        );

    \I__10470\ : Span4Mux_v
    port map (
            O => \N__49156\,
            I => \N__49104\
        );

    \I__10469\ : Span4Mux_h
    port map (
            O => \N__49153\,
            I => \N__49097\
        );

    \I__10468\ : Span4Mux_v
    port map (
            O => \N__49150\,
            I => \N__49097\
        );

    \I__10467\ : Span4Mux_h
    port map (
            O => \N__49145\,
            I => \N__49097\
        );

    \I__10466\ : InMux
    port map (
            O => \N__49144\,
            I => \N__49094\
        );

    \I__10465\ : Span12Mux_h
    port map (
            O => \N__49141\,
            I => \N__49087\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__49136\,
            I => \N__49087\
        );

    \I__10463\ : LocalMux
    port map (
            O => \N__49133\,
            I => \N__49087\
        );

    \I__10462\ : Span4Mux_h
    port map (
            O => \N__49130\,
            I => \N__49084\
        );

    \I__10461\ : Span12Mux_h
    port map (
            O => \N__49125\,
            I => \N__49081\
        );

    \I__10460\ : Span4Mux_h
    port map (
            O => \N__49122\,
            I => \N__49076\
        );

    \I__10459\ : Span4Mux_v
    port map (
            O => \N__49119\,
            I => \N__49076\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__49116\,
            I => \N__49071\
        );

    \I__10457\ : Span12Mux_v
    port map (
            O => \N__49111\,
            I => \N__49071\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__49104\,
            I => \N__49066\
        );

    \I__10455\ : Span4Mux_v
    port map (
            O => \N__49097\,
            I => \N__49066\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__49094\,
            I => \N__49061\
        );

    \I__10453\ : Span12Mux_v
    port map (
            O => \N__49087\,
            I => \N__49061\
        );

    \I__10452\ : Odrv4
    port map (
            O => \N__49084\,
            I => \FRAME_MATCHER_state_31_N_2976_2\
        );

    \I__10451\ : Odrv12
    port map (
            O => \N__49081\,
            I => \FRAME_MATCHER_state_31_N_2976_2\
        );

    \I__10450\ : Odrv4
    port map (
            O => \N__49076\,
            I => \FRAME_MATCHER_state_31_N_2976_2\
        );

    \I__10449\ : Odrv12
    port map (
            O => \N__49071\,
            I => \FRAME_MATCHER_state_31_N_2976_2\
        );

    \I__10448\ : Odrv4
    port map (
            O => \N__49066\,
            I => \FRAME_MATCHER_state_31_N_2976_2\
        );

    \I__10447\ : Odrv12
    port map (
            O => \N__49061\,
            I => \FRAME_MATCHER_state_31_N_2976_2\
        );

    \I__10446\ : InMux
    port map (
            O => \N__49048\,
            I => \N__49041\
        );

    \I__10445\ : CascadeMux
    port map (
            O => \N__49047\,
            I => \N__49037\
        );

    \I__10444\ : InMux
    port map (
            O => \N__49046\,
            I => \N__49030\
        );

    \I__10443\ : InMux
    port map (
            O => \N__49045\,
            I => \N__49030\
        );

    \I__10442\ : InMux
    port map (
            O => \N__49044\,
            I => \N__49030\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__49041\,
            I => \N__49027\
        );

    \I__10440\ : InMux
    port map (
            O => \N__49040\,
            I => \N__49014\
        );

    \I__10439\ : InMux
    port map (
            O => \N__49037\,
            I => \N__49009\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__49030\,
            I => \N__48994\
        );

    \I__10437\ : Span4Mux_v
    port map (
            O => \N__49027\,
            I => \N__48994\
        );

    \I__10436\ : InMux
    port map (
            O => \N__49026\,
            I => \N__48987\
        );

    \I__10435\ : InMux
    port map (
            O => \N__49025\,
            I => \N__48987\
        );

    \I__10434\ : InMux
    port map (
            O => \N__49024\,
            I => \N__48987\
        );

    \I__10433\ : InMux
    port map (
            O => \N__49023\,
            I => \N__48982\
        );

    \I__10432\ : InMux
    port map (
            O => \N__49022\,
            I => \N__48982\
        );

    \I__10431\ : InMux
    port map (
            O => \N__49021\,
            I => \N__48971\
        );

    \I__10430\ : InMux
    port map (
            O => \N__49020\,
            I => \N__48965\
        );

    \I__10429\ : InMux
    port map (
            O => \N__49019\,
            I => \N__48962\
        );

    \I__10428\ : InMux
    port map (
            O => \N__49018\,
            I => \N__48957\
        );

    \I__10427\ : InMux
    port map (
            O => \N__49017\,
            I => \N__48957\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__49014\,
            I => \N__48954\
        );

    \I__10425\ : InMux
    port map (
            O => \N__49013\,
            I => \N__48950\
        );

    \I__10424\ : InMux
    port map (
            O => \N__49012\,
            I => \N__48940\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__49009\,
            I => \N__48935\
        );

    \I__10422\ : InMux
    port map (
            O => \N__49008\,
            I => \N__48928\
        );

    \I__10421\ : InMux
    port map (
            O => \N__49007\,
            I => \N__48928\
        );

    \I__10420\ : InMux
    port map (
            O => \N__49006\,
            I => \N__48923\
        );

    \I__10419\ : InMux
    port map (
            O => \N__49005\,
            I => \N__48923\
        );

    \I__10418\ : InMux
    port map (
            O => \N__49004\,
            I => \N__48916\
        );

    \I__10417\ : InMux
    port map (
            O => \N__49003\,
            I => \N__48916\
        );

    \I__10416\ : InMux
    port map (
            O => \N__49002\,
            I => \N__48916\
        );

    \I__10415\ : InMux
    port map (
            O => \N__49001\,
            I => \N__48909\
        );

    \I__10414\ : InMux
    port map (
            O => \N__49000\,
            I => \N__48909\
        );

    \I__10413\ : InMux
    port map (
            O => \N__48999\,
            I => \N__48909\
        );

    \I__10412\ : Span4Mux_v
    port map (
            O => \N__48994\,
            I => \N__48904\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__48987\,
            I => \N__48904\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__48982\,
            I => \N__48901\
        );

    \I__10409\ : CascadeMux
    port map (
            O => \N__48981\,
            I => \N__48898\
        );

    \I__10408\ : InMux
    port map (
            O => \N__48980\,
            I => \N__48892\
        );

    \I__10407\ : InMux
    port map (
            O => \N__48979\,
            I => \N__48877\
        );

    \I__10406\ : InMux
    port map (
            O => \N__48978\,
            I => \N__48877\
        );

    \I__10405\ : InMux
    port map (
            O => \N__48977\,
            I => \N__48877\
        );

    \I__10404\ : InMux
    port map (
            O => \N__48976\,
            I => \N__48877\
        );

    \I__10403\ : InMux
    port map (
            O => \N__48975\,
            I => \N__48872\
        );

    \I__10402\ : InMux
    port map (
            O => \N__48974\,
            I => \N__48872\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__48971\,
            I => \N__48869\
        );

    \I__10400\ : InMux
    port map (
            O => \N__48970\,
            I => \N__48864\
        );

    \I__10399\ : InMux
    port map (
            O => \N__48969\,
            I => \N__48864\
        );

    \I__10398\ : InMux
    port map (
            O => \N__48968\,
            I => \N__48861\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__48965\,
            I => \N__48858\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__48962\,
            I => \N__48851\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__48957\,
            I => \N__48851\
        );

    \I__10394\ : Span4Mux_h
    port map (
            O => \N__48954\,
            I => \N__48851\
        );

    \I__10393\ : CascadeMux
    port map (
            O => \N__48953\,
            I => \N__48848\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__48950\,
            I => \N__48841\
        );

    \I__10391\ : InMux
    port map (
            O => \N__48949\,
            I => \N__48834\
        );

    \I__10390\ : InMux
    port map (
            O => \N__48948\,
            I => \N__48834\
        );

    \I__10389\ : InMux
    port map (
            O => \N__48947\,
            I => \N__48834\
        );

    \I__10388\ : InMux
    port map (
            O => \N__48946\,
            I => \N__48830\
        );

    \I__10387\ : InMux
    port map (
            O => \N__48945\,
            I => \N__48827\
        );

    \I__10386\ : InMux
    port map (
            O => \N__48944\,
            I => \N__48822\
        );

    \I__10385\ : InMux
    port map (
            O => \N__48943\,
            I => \N__48822\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__48940\,
            I => \N__48819\
        );

    \I__10383\ : InMux
    port map (
            O => \N__48939\,
            I => \N__48814\
        );

    \I__10382\ : InMux
    port map (
            O => \N__48938\,
            I => \N__48814\
        );

    \I__10381\ : Span4Mux_v
    port map (
            O => \N__48935\,
            I => \N__48811\
        );

    \I__10380\ : InMux
    port map (
            O => \N__48934\,
            I => \N__48806\
        );

    \I__10379\ : InMux
    port map (
            O => \N__48933\,
            I => \N__48806\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__48928\,
            I => \N__48801\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__48923\,
            I => \N__48801\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__48916\,
            I => \N__48792\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__48909\,
            I => \N__48792\
        );

    \I__10374\ : Span4Mux_h
    port map (
            O => \N__48904\,
            I => \N__48792\
        );

    \I__10373\ : Span4Mux_h
    port map (
            O => \N__48901\,
            I => \N__48792\
        );

    \I__10372\ : InMux
    port map (
            O => \N__48898\,
            I => \N__48789\
        );

    \I__10371\ : InMux
    port map (
            O => \N__48897\,
            I => \N__48783\
        );

    \I__10370\ : InMux
    port map (
            O => \N__48896\,
            I => \N__48783\
        );

    \I__10369\ : InMux
    port map (
            O => \N__48895\,
            I => \N__48780\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__48892\,
            I => \N__48777\
        );

    \I__10367\ : InMux
    port map (
            O => \N__48891\,
            I => \N__48770\
        );

    \I__10366\ : InMux
    port map (
            O => \N__48890\,
            I => \N__48770\
        );

    \I__10365\ : InMux
    port map (
            O => \N__48889\,
            I => \N__48770\
        );

    \I__10364\ : InMux
    port map (
            O => \N__48888\,
            I => \N__48763\
        );

    \I__10363\ : InMux
    port map (
            O => \N__48887\,
            I => \N__48763\
        );

    \I__10362\ : InMux
    port map (
            O => \N__48886\,
            I => \N__48763\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__48877\,
            I => \N__48754\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__48872\,
            I => \N__48754\
        );

    \I__10359\ : Span4Mux_h
    port map (
            O => \N__48869\,
            I => \N__48754\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__48864\,
            I => \N__48754\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__48861\,
            I => \N__48747\
        );

    \I__10356\ : Span4Mux_h
    port map (
            O => \N__48858\,
            I => \N__48747\
        );

    \I__10355\ : Span4Mux_v
    port map (
            O => \N__48851\,
            I => \N__48747\
        );

    \I__10354\ : InMux
    port map (
            O => \N__48848\,
            I => \N__48744\
        );

    \I__10353\ : InMux
    port map (
            O => \N__48847\,
            I => \N__48728\
        );

    \I__10352\ : InMux
    port map (
            O => \N__48846\,
            I => \N__48728\
        );

    \I__10351\ : InMux
    port map (
            O => \N__48845\,
            I => \N__48723\
        );

    \I__10350\ : InMux
    port map (
            O => \N__48844\,
            I => \N__48723\
        );

    \I__10349\ : Span4Mux_h
    port map (
            O => \N__48841\,
            I => \N__48720\
        );

    \I__10348\ : LocalMux
    port map (
            O => \N__48834\,
            I => \N__48717\
        );

    \I__10347\ : InMux
    port map (
            O => \N__48833\,
            I => \N__48714\
        );

    \I__10346\ : LocalMux
    port map (
            O => \N__48830\,
            I => \N__48709\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__48827\,
            I => \N__48709\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__48822\,
            I => \N__48706\
        );

    \I__10343\ : Span4Mux_h
    port map (
            O => \N__48819\,
            I => \N__48703\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__48814\,
            I => \N__48698\
        );

    \I__10341\ : Span4Mux_v
    port map (
            O => \N__48811\,
            I => \N__48698\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__48806\,
            I => \N__48690\
        );

    \I__10339\ : Span4Mux_h
    port map (
            O => \N__48801\,
            I => \N__48690\
        );

    \I__10338\ : Span4Mux_v
    port map (
            O => \N__48792\,
            I => \N__48690\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__48789\,
            I => \N__48687\
        );

    \I__10336\ : InMux
    port map (
            O => \N__48788\,
            I => \N__48684\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__48783\,
            I => \N__48681\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__48780\,
            I => \N__48676\
        );

    \I__10333\ : Span4Mux_v
    port map (
            O => \N__48777\,
            I => \N__48676\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__48770\,
            I => \N__48667\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__48763\,
            I => \N__48667\
        );

    \I__10330\ : Span4Mux_v
    port map (
            O => \N__48754\,
            I => \N__48667\
        );

    \I__10329\ : Span4Mux_v
    port map (
            O => \N__48747\,
            I => \N__48667\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__48744\,
            I => \N__48664\
        );

    \I__10327\ : InMux
    port map (
            O => \N__48743\,
            I => \N__48659\
        );

    \I__10326\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48659\
        );

    \I__10325\ : InMux
    port map (
            O => \N__48741\,
            I => \N__48656\
        );

    \I__10324\ : InMux
    port map (
            O => \N__48740\,
            I => \N__48647\
        );

    \I__10323\ : InMux
    port map (
            O => \N__48739\,
            I => \N__48647\
        );

    \I__10322\ : InMux
    port map (
            O => \N__48738\,
            I => \N__48647\
        );

    \I__10321\ : InMux
    port map (
            O => \N__48737\,
            I => \N__48647\
        );

    \I__10320\ : InMux
    port map (
            O => \N__48736\,
            I => \N__48642\
        );

    \I__10319\ : InMux
    port map (
            O => \N__48735\,
            I => \N__48642\
        );

    \I__10318\ : InMux
    port map (
            O => \N__48734\,
            I => \N__48637\
        );

    \I__10317\ : InMux
    port map (
            O => \N__48733\,
            I => \N__48637\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__48728\,
            I => \N__48632\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__48723\,
            I => \N__48632\
        );

    \I__10314\ : Span4Mux_v
    port map (
            O => \N__48720\,
            I => \N__48629\
        );

    \I__10313\ : Span12Mux_s11_v
    port map (
            O => \N__48717\,
            I => \N__48626\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__48714\,
            I => \N__48615\
        );

    \I__10311\ : Span4Mux_h
    port map (
            O => \N__48709\,
            I => \N__48615\
        );

    \I__10310\ : Span4Mux_h
    port map (
            O => \N__48706\,
            I => \N__48615\
        );

    \I__10309\ : Span4Mux_h
    port map (
            O => \N__48703\,
            I => \N__48615\
        );

    \I__10308\ : Span4Mux_h
    port map (
            O => \N__48698\,
            I => \N__48615\
        );

    \I__10307\ : InMux
    port map (
            O => \N__48697\,
            I => \N__48612\
        );

    \I__10306\ : Span4Mux_h
    port map (
            O => \N__48690\,
            I => \N__48605\
        );

    \I__10305\ : Span4Mux_h
    port map (
            O => \N__48687\,
            I => \N__48605\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__48684\,
            I => \N__48605\
        );

    \I__10303\ : Span4Mux_h
    port map (
            O => \N__48681\,
            I => \N__48596\
        );

    \I__10302\ : Span4Mux_v
    port map (
            O => \N__48676\,
            I => \N__48596\
        );

    \I__10301\ : Span4Mux_h
    port map (
            O => \N__48667\,
            I => \N__48596\
        );

    \I__10300\ : Span4Mux_h
    port map (
            O => \N__48664\,
            I => \N__48596\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__48659\,
            I => n22661
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__48656\,
            I => n22661
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__48647\,
            I => n22661
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__48642\,
            I => n22661
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__48637\,
            I => n22661
        );

    \I__10294\ : Odrv12
    port map (
            O => \N__48632\,
            I => n22661
        );

    \I__10293\ : Odrv4
    port map (
            O => \N__48629\,
            I => n22661
        );

    \I__10292\ : Odrv12
    port map (
            O => \N__48626\,
            I => n22661
        );

    \I__10291\ : Odrv4
    port map (
            O => \N__48615\,
            I => n22661
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__48612\,
            I => n22661
        );

    \I__10289\ : Odrv4
    port map (
            O => \N__48605\,
            I => n22661
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__48596\,
            I => n22661
        );

    \I__10287\ : CascadeMux
    port map (
            O => \N__48571\,
            I => \N__48567\
        );

    \I__10286\ : CascadeMux
    port map (
            O => \N__48570\,
            I => \N__48563\
        );

    \I__10285\ : InMux
    port map (
            O => \N__48567\,
            I => \N__48559\
        );

    \I__10284\ : CascadeMux
    port map (
            O => \N__48566\,
            I => \N__48554\
        );

    \I__10283\ : InMux
    port map (
            O => \N__48563\,
            I => \N__48548\
        );

    \I__10282\ : InMux
    port map (
            O => \N__48562\,
            I => \N__48545\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__48559\,
            I => \N__48542\
        );

    \I__10280\ : InMux
    port map (
            O => \N__48558\,
            I => \N__48537\
        );

    \I__10279\ : InMux
    port map (
            O => \N__48557\,
            I => \N__48537\
        );

    \I__10278\ : InMux
    port map (
            O => \N__48554\,
            I => \N__48534\
        );

    \I__10277\ : InMux
    port map (
            O => \N__48553\,
            I => \N__48530\
        );

    \I__10276\ : InMux
    port map (
            O => \N__48552\,
            I => \N__48527\
        );

    \I__10275\ : InMux
    port map (
            O => \N__48551\,
            I => \N__48524\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__48548\,
            I => \N__48519\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__48545\,
            I => \N__48519\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__48542\,
            I => \N__48516\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__48537\,
            I => \N__48511\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__48534\,
            I => \N__48511\
        );

    \I__10269\ : InMux
    port map (
            O => \N__48533\,
            I => \N__48508\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__48530\,
            I => \N__48503\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__48527\,
            I => \N__48503\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__48524\,
            I => \N__48498\
        );

    \I__10265\ : Span4Mux_h
    port map (
            O => \N__48519\,
            I => \N__48498\
        );

    \I__10264\ : Span4Mux_h
    port map (
            O => \N__48516\,
            I => \N__48493\
        );

    \I__10263\ : Span4Mux_h
    port map (
            O => \N__48511\,
            I => \N__48493\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__48508\,
            I => encoder0_position_30
        );

    \I__10261\ : Odrv4
    port map (
            O => \N__48503\,
            I => encoder0_position_30
        );

    \I__10260\ : Odrv4
    port map (
            O => \N__48498\,
            I => encoder0_position_30
        );

    \I__10259\ : Odrv4
    port map (
            O => \N__48493\,
            I => encoder0_position_30
        );

    \I__10258\ : InMux
    port map (
            O => \N__48484\,
            I => \N__48481\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__48481\,
            I => \N__48477\
        );

    \I__10256\ : InMux
    port map (
            O => \N__48480\,
            I => \N__48474\
        );

    \I__10255\ : Span4Mux_h
    port map (
            O => \N__48477\,
            I => \N__48471\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__48474\,
            I => data_out_frame_6_6
        );

    \I__10253\ : Odrv4
    port map (
            O => \N__48471\,
            I => data_out_frame_6_6
        );

    \I__10252\ : CascadeMux
    port map (
            O => \N__48466\,
            I => \N__48463\
        );

    \I__10251\ : InMux
    port map (
            O => \N__48463\,
            I => \N__48460\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__48460\,
            I => \N__48457\
        );

    \I__10249\ : Span4Mux_v
    port map (
            O => \N__48457\,
            I => \N__48454\
        );

    \I__10248\ : Odrv4
    port map (
            O => \N__48454\,
            I => \c0.n6_adj_4241\
        );

    \I__10247\ : InMux
    port map (
            O => \N__48451\,
            I => \N__48445\
        );

    \I__10246\ : InMux
    port map (
            O => \N__48450\,
            I => \N__48442\
        );

    \I__10245\ : InMux
    port map (
            O => \N__48449\,
            I => \N__48437\
        );

    \I__10244\ : InMux
    port map (
            O => \N__48448\,
            I => \N__48437\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__48445\,
            I => \N__48434\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__48442\,
            I => \N__48431\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__48437\,
            I => \N__48428\
        );

    \I__10240\ : Span4Mux_h
    port map (
            O => \N__48434\,
            I => \N__48425\
        );

    \I__10239\ : Span4Mux_v
    port map (
            O => \N__48431\,
            I => \N__48420\
        );

    \I__10238\ : Span4Mux_h
    port map (
            O => \N__48428\,
            I => \N__48420\
        );

    \I__10237\ : Odrv4
    port map (
            O => \N__48425\,
            I => \c0.n13086\
        );

    \I__10236\ : Odrv4
    port map (
            O => \N__48420\,
            I => \c0.n13086\
        );

    \I__10235\ : CascadeMux
    port map (
            O => \N__48415\,
            I => \N__48411\
        );

    \I__10234\ : InMux
    port map (
            O => \N__48414\,
            I => \N__48405\
        );

    \I__10233\ : InMux
    port map (
            O => \N__48411\,
            I => \N__48405\
        );

    \I__10232\ : CascadeMux
    port map (
            O => \N__48410\,
            I => \N__48402\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__48405\,
            I => \N__48398\
        );

    \I__10230\ : InMux
    port map (
            O => \N__48402\,
            I => \N__48393\
        );

    \I__10229\ : InMux
    port map (
            O => \N__48401\,
            I => \N__48393\
        );

    \I__10228\ : Odrv12
    port map (
            O => \N__48398\,
            I => \c0.data_in_frame_8_5\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__48393\,
            I => \c0.data_in_frame_8_5\
        );

    \I__10226\ : CascadeMux
    port map (
            O => \N__48388\,
            I => \c0.n22415_cascade_\
        );

    \I__10225\ : CascadeMux
    port map (
            O => \N__48385\,
            I => \N__48380\
        );

    \I__10224\ : InMux
    port map (
            O => \N__48384\,
            I => \N__48375\
        );

    \I__10223\ : InMux
    port map (
            O => \N__48383\,
            I => \N__48375\
        );

    \I__10222\ : InMux
    port map (
            O => \N__48380\,
            I => \N__48372\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__48375\,
            I => \N__48369\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__48372\,
            I => \c0.data_in_frame_10_5\
        );

    \I__10219\ : Odrv4
    port map (
            O => \N__48369\,
            I => \c0.data_in_frame_10_5\
        );

    \I__10218\ : InMux
    port map (
            O => \N__48364\,
            I => \N__48361\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__48361\,
            I => \N__48358\
        );

    \I__10216\ : Odrv12
    port map (
            O => \N__48358\,
            I => \c0.n35\
        );

    \I__10215\ : CascadeMux
    port map (
            O => \N__48355\,
            I => \c0.n13771_cascade_\
        );

    \I__10214\ : InMux
    port map (
            O => \N__48352\,
            I => \N__48346\
        );

    \I__10213\ : InMux
    port map (
            O => \N__48351\,
            I => \N__48346\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__48346\,
            I => \c0.n22239\
        );

    \I__10211\ : CascadeMux
    port map (
            O => \N__48343\,
            I => \c0.n4_cascade_\
        );

    \I__10210\ : InMux
    port map (
            O => \N__48340\,
            I => \N__48337\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__48337\,
            I => \c0.n37\
        );

    \I__10208\ : InMux
    port map (
            O => \N__48334\,
            I => \N__48331\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__48331\,
            I => \N__48328\
        );

    \I__10206\ : Span4Mux_h
    port map (
            O => \N__48328\,
            I => \N__48325\
        );

    \I__10205\ : Odrv4
    port map (
            O => \N__48325\,
            I => \c0.n6_adj_4220\
        );

    \I__10204\ : CascadeMux
    port map (
            O => \N__48322\,
            I => \N__48318\
        );

    \I__10203\ : CascadeMux
    port map (
            O => \N__48321\,
            I => \N__48314\
        );

    \I__10202\ : InMux
    port map (
            O => \N__48318\,
            I => \N__48311\
        );

    \I__10201\ : CascadeMux
    port map (
            O => \N__48317\,
            I => \N__48308\
        );

    \I__10200\ : InMux
    port map (
            O => \N__48314\,
            I => \N__48305\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__48311\,
            I => \N__48302\
        );

    \I__10198\ : InMux
    port map (
            O => \N__48308\,
            I => \N__48299\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__48305\,
            I => \c0.data_in_frame_8_3\
        );

    \I__10196\ : Odrv12
    port map (
            O => \N__48302\,
            I => \c0.data_in_frame_8_3\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__48299\,
            I => \c0.data_in_frame_8_3\
        );

    \I__10194\ : InMux
    port map (
            O => \N__48292\,
            I => \N__48289\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__48289\,
            I => \c0.n13652\
        );

    \I__10192\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48283\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__48283\,
            I => \c0.n13771\
        );

    \I__10190\ : InMux
    port map (
            O => \N__48280\,
            I => \N__48274\
        );

    \I__10189\ : InMux
    port map (
            O => \N__48279\,
            I => \N__48274\
        );

    \I__10188\ : LocalMux
    port map (
            O => \N__48274\,
            I => \c0.data_in_frame_10_3\
        );

    \I__10187\ : CascadeMux
    port map (
            O => \N__48271\,
            I => \N__48268\
        );

    \I__10186\ : InMux
    port map (
            O => \N__48268\,
            I => \N__48265\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__48265\,
            I => \c0.n21964\
        );

    \I__10184\ : InMux
    port map (
            O => \N__48262\,
            I => \N__48259\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__48259\,
            I => \N__48256\
        );

    \I__10182\ : Span4Mux_h
    port map (
            O => \N__48256\,
            I => \N__48252\
        );

    \I__10181\ : InMux
    port map (
            O => \N__48255\,
            I => \N__48249\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__48252\,
            I => \c0.n22280\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__48249\,
            I => \c0.n22280\
        );

    \I__10178\ : CascadeMux
    port map (
            O => \N__48244\,
            I => \c0.n21964_cascade_\
        );

    \I__10177\ : InMux
    port map (
            O => \N__48241\,
            I => \N__48237\
        );

    \I__10176\ : InMux
    port map (
            O => \N__48240\,
            I => \N__48234\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__48237\,
            I => \N__48229\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__48234\,
            I => \N__48226\
        );

    \I__10173\ : InMux
    port map (
            O => \N__48233\,
            I => \N__48221\
        );

    \I__10172\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48221\
        );

    \I__10171\ : Span4Mux_h
    port map (
            O => \N__48229\,
            I => \N__48216\
        );

    \I__10170\ : Span4Mux_h
    port map (
            O => \N__48226\,
            I => \N__48216\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__48221\,
            I => \N__48213\
        );

    \I__10168\ : Odrv4
    port map (
            O => \N__48216\,
            I => \c0.n14113\
        );

    \I__10167\ : Odrv4
    port map (
            O => \N__48213\,
            I => \c0.n14113\
        );

    \I__10166\ : CascadeMux
    port map (
            O => \N__48208\,
            I => \N__48205\
        );

    \I__10165\ : InMux
    port map (
            O => \N__48205\,
            I => \N__48201\
        );

    \I__10164\ : CascadeMux
    port map (
            O => \N__48204\,
            I => \N__48198\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__48201\,
            I => \N__48193\
        );

    \I__10162\ : InMux
    port map (
            O => \N__48198\,
            I => \N__48190\
        );

    \I__10161\ : InMux
    port map (
            O => \N__48197\,
            I => \N__48185\
        );

    \I__10160\ : InMux
    port map (
            O => \N__48196\,
            I => \N__48185\
        );

    \I__10159\ : Span4Mux_h
    port map (
            O => \N__48193\,
            I => \N__48182\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__48190\,
            I => \N__48177\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__48185\,
            I => \N__48177\
        );

    \I__10156\ : Odrv4
    port map (
            O => \N__48182\,
            I => \c0.data_in_frame_2_5\
        );

    \I__10155\ : Odrv4
    port map (
            O => \N__48177\,
            I => \c0.data_in_frame_2_5\
        );

    \I__10154\ : CascadeMux
    port map (
            O => \N__48172\,
            I => \N__48165\
        );

    \I__10153\ : CascadeMux
    port map (
            O => \N__48171\,
            I => \N__48162\
        );

    \I__10152\ : CascadeMux
    port map (
            O => \N__48170\,
            I => \N__48159\
        );

    \I__10151\ : CascadeMux
    port map (
            O => \N__48169\,
            I => \N__48155\
        );

    \I__10150\ : CascadeMux
    port map (
            O => \N__48168\,
            I => \N__48150\
        );

    \I__10149\ : InMux
    port map (
            O => \N__48165\,
            I => \N__48145\
        );

    \I__10148\ : InMux
    port map (
            O => \N__48162\,
            I => \N__48145\
        );

    \I__10147\ : InMux
    port map (
            O => \N__48159\,
            I => \N__48140\
        );

    \I__10146\ : InMux
    port map (
            O => \N__48158\,
            I => \N__48140\
        );

    \I__10145\ : InMux
    port map (
            O => \N__48155\,
            I => \N__48134\
        );

    \I__10144\ : InMux
    port map (
            O => \N__48154\,
            I => \N__48134\
        );

    \I__10143\ : CascadeMux
    port map (
            O => \N__48153\,
            I => \N__48131\
        );

    \I__10142\ : InMux
    port map (
            O => \N__48150\,
            I => \N__48128\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__48145\,
            I => \N__48125\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__48140\,
            I => \N__48122\
        );

    \I__10139\ : InMux
    port map (
            O => \N__48139\,
            I => \N__48119\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__48134\,
            I => \N__48116\
        );

    \I__10137\ : InMux
    port map (
            O => \N__48131\,
            I => \N__48113\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__48128\,
            I => \N__48108\
        );

    \I__10135\ : Span4Mux_v
    port map (
            O => \N__48125\,
            I => \N__48108\
        );

    \I__10134\ : Span4Mux_h
    port map (
            O => \N__48122\,
            I => \N__48101\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__48119\,
            I => \N__48101\
        );

    \I__10132\ : Span4Mux_v
    port map (
            O => \N__48116\,
            I => \N__48101\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__48113\,
            I => \c0.data_in_frame_0_3\
        );

    \I__10130\ : Odrv4
    port map (
            O => \N__48108\,
            I => \c0.data_in_frame_0_3\
        );

    \I__10129\ : Odrv4
    port map (
            O => \N__48101\,
            I => \c0.data_in_frame_0_3\
        );

    \I__10128\ : CascadeMux
    port map (
            O => \N__48094\,
            I => \N__48091\
        );

    \I__10127\ : InMux
    port map (
            O => \N__48091\,
            I => \N__48081\
        );

    \I__10126\ : InMux
    port map (
            O => \N__48090\,
            I => \N__48081\
        );

    \I__10125\ : InMux
    port map (
            O => \N__48089\,
            I => \N__48081\
        );

    \I__10124\ : InMux
    port map (
            O => \N__48088\,
            I => \N__48078\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__48081\,
            I => \N__48075\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__48078\,
            I => \N__48072\
        );

    \I__10121\ : Span4Mux_v
    port map (
            O => \N__48075\,
            I => \N__48069\
        );

    \I__10120\ : Span4Mux_v
    port map (
            O => \N__48072\,
            I => \N__48066\
        );

    \I__10119\ : Span4Mux_h
    port map (
            O => \N__48069\,
            I => \N__48063\
        );

    \I__10118\ : Odrv4
    port map (
            O => \N__48066\,
            I => \c0.n13398\
        );

    \I__10117\ : Odrv4
    port map (
            O => \N__48063\,
            I => \c0.n13398\
        );

    \I__10116\ : InMux
    port map (
            O => \N__48058\,
            I => \N__48055\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__48055\,
            I => \N__48052\
        );

    \I__10114\ : Span4Mux_v
    port map (
            O => \N__48052\,
            I => \N__48049\
        );

    \I__10113\ : Span4Mux_h
    port map (
            O => \N__48049\,
            I => \N__48043\
        );

    \I__10112\ : InMux
    port map (
            O => \N__48048\,
            I => \N__48040\
        );

    \I__10111\ : CascadeMux
    port map (
            O => \N__48047\,
            I => \N__48037\
        );

    \I__10110\ : InMux
    port map (
            O => \N__48046\,
            I => \N__48034\
        );

    \I__10109\ : Span4Mux_v
    port map (
            O => \N__48043\,
            I => \N__48029\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__48040\,
            I => \N__48029\
        );

    \I__10107\ : InMux
    port map (
            O => \N__48037\,
            I => \N__48023\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__48034\,
            I => \N__48018\
        );

    \I__10105\ : Span4Mux_h
    port map (
            O => \N__48029\,
            I => \N__48018\
        );

    \I__10104\ : InMux
    port map (
            O => \N__48028\,
            I => \N__48015\
        );

    \I__10103\ : InMux
    port map (
            O => \N__48027\,
            I => \N__48010\
        );

    \I__10102\ : InMux
    port map (
            O => \N__48026\,
            I => \N__48010\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__48023\,
            I => data_in_frame_1_3
        );

    \I__10100\ : Odrv4
    port map (
            O => \N__48018\,
            I => data_in_frame_1_3
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__48015\,
            I => data_in_frame_1_3
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__48010\,
            I => data_in_frame_1_3
        );

    \I__10097\ : InMux
    port map (
            O => \N__48001\,
            I => \N__47998\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__47998\,
            I => \N__47994\
        );

    \I__10095\ : InMux
    port map (
            O => \N__47997\,
            I => \N__47989\
        );

    \I__10094\ : Span4Mux_h
    port map (
            O => \N__47994\,
            I => \N__47986\
        );

    \I__10093\ : InMux
    port map (
            O => \N__47993\,
            I => \N__47983\
        );

    \I__10092\ : InMux
    port map (
            O => \N__47992\,
            I => \N__47980\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__47989\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10090\ : Odrv4
    port map (
            O => \N__47986\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__47983\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__47980\,
            I => \c0.data_in_frame_3_5\
        );

    \I__10087\ : CascadeMux
    port map (
            O => \N__47971\,
            I => \c0.n13398_cascade_\
        );

    \I__10086\ : InMux
    port map (
            O => \N__47968\,
            I => \N__47962\
        );

    \I__10085\ : InMux
    port map (
            O => \N__47967\,
            I => \N__47962\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__47962\,
            I => \N__47959\
        );

    \I__10083\ : Odrv4
    port map (
            O => \N__47959\,
            I => \c0.n13852\
        );

    \I__10082\ : InMux
    port map (
            O => \N__47956\,
            I => \N__47953\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__47953\,
            I => \N__47950\
        );

    \I__10080\ : Span4Mux_h
    port map (
            O => \N__47950\,
            I => \N__47946\
        );

    \I__10079\ : InMux
    port map (
            O => \N__47949\,
            I => \N__47943\
        );

    \I__10078\ : Odrv4
    port map (
            O => \N__47946\,
            I => \c0.n21794\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__47943\,
            I => \c0.n21794\
        );

    \I__10076\ : InMux
    port map (
            O => \N__47938\,
            I => \N__47934\
        );

    \I__10075\ : CascadeMux
    port map (
            O => \N__47937\,
            I => \N__47931\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__47934\,
            I => \N__47927\
        );

    \I__10073\ : InMux
    port map (
            O => \N__47931\,
            I => \N__47924\
        );

    \I__10072\ : InMux
    port map (
            O => \N__47930\,
            I => \N__47921\
        );

    \I__10071\ : Span4Mux_h
    port map (
            O => \N__47927\,
            I => \N__47918\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__47924\,
            I => \c0.data_in_frame_8_2\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__47921\,
            I => \c0.data_in_frame_8_2\
        );

    \I__10068\ : Odrv4
    port map (
            O => \N__47918\,
            I => \c0.data_in_frame_8_2\
        );

    \I__10067\ : CascadeMux
    port map (
            O => \N__47911\,
            I => \c0.n21794_cascade_\
        );

    \I__10066\ : InMux
    port map (
            O => \N__47908\,
            I => \N__47903\
        );

    \I__10065\ : CascadeMux
    port map (
            O => \N__47907\,
            I => \N__47898\
        );

    \I__10064\ : InMux
    port map (
            O => \N__47906\,
            I => \N__47895\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__47903\,
            I => \N__47892\
        );

    \I__10062\ : InMux
    port map (
            O => \N__47902\,
            I => \N__47889\
        );

    \I__10061\ : InMux
    port map (
            O => \N__47901\,
            I => \N__47884\
        );

    \I__10060\ : InMux
    port map (
            O => \N__47898\,
            I => \N__47884\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__47895\,
            I => \N__47880\
        );

    \I__10058\ : Span4Mux_v
    port map (
            O => \N__47892\,
            I => \N__47877\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__47889\,
            I => \N__47874\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__47884\,
            I => \N__47871\
        );

    \I__10055\ : InMux
    port map (
            O => \N__47883\,
            I => \N__47868\
        );

    \I__10054\ : Sp12to4
    port map (
            O => \N__47880\,
            I => \N__47865\
        );

    \I__10053\ : Span4Mux_v
    port map (
            O => \N__47877\,
            I => \N__47860\
        );

    \I__10052\ : Span4Mux_v
    port map (
            O => \N__47874\,
            I => \N__47860\
        );

    \I__10051\ : Span4Mux_h
    port map (
            O => \N__47871\,
            I => \N__47857\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__47868\,
            I => \c0.data_in_frame_5_7\
        );

    \I__10049\ : Odrv12
    port map (
            O => \N__47865\,
            I => \c0.data_in_frame_5_7\
        );

    \I__10048\ : Odrv4
    port map (
            O => \N__47860\,
            I => \c0.data_in_frame_5_7\
        );

    \I__10047\ : Odrv4
    port map (
            O => \N__47857\,
            I => \c0.data_in_frame_5_7\
        );

    \I__10046\ : CascadeMux
    port map (
            O => \N__47848\,
            I => \c0.n6_adj_4257_cascade_\
        );

    \I__10045\ : InMux
    port map (
            O => \N__47845\,
            I => \N__47841\
        );

    \I__10044\ : InMux
    port map (
            O => \N__47844\,
            I => \N__47838\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__47841\,
            I => \N__47835\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__47838\,
            I => \N__47830\
        );

    \I__10041\ : Span4Mux_h
    port map (
            O => \N__47835\,
            I => \N__47830\
        );

    \I__10040\ : Odrv4
    port map (
            O => \N__47830\,
            I => \c0.n21825\
        );

    \I__10039\ : InMux
    port map (
            O => \N__47827\,
            I => \N__47824\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__47824\,
            I => \N__47820\
        );

    \I__10037\ : InMux
    port map (
            O => \N__47823\,
            I => \N__47817\
        );

    \I__10036\ : Span4Mux_h
    port map (
            O => \N__47820\,
            I => \N__47814\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__47817\,
            I => \c0.data_in_frame_9_5\
        );

    \I__10034\ : Odrv4
    port map (
            O => \N__47814\,
            I => \c0.data_in_frame_9_5\
        );

    \I__10033\ : CascadeMux
    port map (
            O => \N__47809\,
            I => \c0.n8_adj_4254_cascade_\
        );

    \I__10032\ : InMux
    port map (
            O => \N__47806\,
            I => \N__47803\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__47803\,
            I => \N__47799\
        );

    \I__10030\ : InMux
    port map (
            O => \N__47802\,
            I => \N__47796\
        );

    \I__10029\ : Span4Mux_h
    port map (
            O => \N__47799\,
            I => \N__47793\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__47796\,
            I => \c0.n4_adj_4255\
        );

    \I__10027\ : Odrv4
    port map (
            O => \N__47793\,
            I => \c0.n4_adj_4255\
        );

    \I__10026\ : CascadeMux
    port map (
            O => \N__47788\,
            I => \N__47784\
        );

    \I__10025\ : CascadeMux
    port map (
            O => \N__47787\,
            I => \N__47781\
        );

    \I__10024\ : InMux
    port map (
            O => \N__47784\,
            I => \N__47778\
        );

    \I__10023\ : InMux
    port map (
            O => \N__47781\,
            I => \N__47775\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__47778\,
            I => \N__47772\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__47775\,
            I => \c0.data_in_frame_5_5\
        );

    \I__10020\ : Odrv4
    port map (
            O => \N__47772\,
            I => \c0.data_in_frame_5_5\
        );

    \I__10019\ : CascadeMux
    port map (
            O => \N__47767\,
            I => \N__47763\
        );

    \I__10018\ : InMux
    port map (
            O => \N__47766\,
            I => \N__47759\
        );

    \I__10017\ : InMux
    port map (
            O => \N__47763\,
            I => \N__47755\
        );

    \I__10016\ : InMux
    port map (
            O => \N__47762\,
            I => \N__47752\
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47749\
        );

    \I__10014\ : InMux
    port map (
            O => \N__47758\,
            I => \N__47746\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__47755\,
            I => \c0.data_in_frame_3_1\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__47752\,
            I => \c0.data_in_frame_3_1\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__47749\,
            I => \c0.data_in_frame_3_1\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__47746\,
            I => \c0.data_in_frame_3_1\
        );

    \I__10009\ : InMux
    port map (
            O => \N__47737\,
            I => \N__47733\
        );

    \I__10008\ : CascadeMux
    port map (
            O => \N__47736\,
            I => \N__47730\
        );

    \I__10007\ : LocalMux
    port map (
            O => \N__47733\,
            I => \N__47727\
        );

    \I__10006\ : InMux
    port map (
            O => \N__47730\,
            I => \N__47722\
        );

    \I__10005\ : Span4Mux_h
    port map (
            O => \N__47727\,
            I => \N__47719\
        );

    \I__10004\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47714\
        );

    \I__10003\ : InMux
    port map (
            O => \N__47725\,
            I => \N__47714\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__47722\,
            I => \c0.data_in_frame_3_2\
        );

    \I__10001\ : Odrv4
    port map (
            O => \N__47719\,
            I => \c0.data_in_frame_3_2\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__47714\,
            I => \c0.data_in_frame_3_2\
        );

    \I__9999\ : InMux
    port map (
            O => \N__47707\,
            I => \N__47704\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__47704\,
            I => \c0.n6_adj_4395\
        );

    \I__9997\ : InMux
    port map (
            O => \N__47701\,
            I => \N__47697\
        );

    \I__9996\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47694\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__47697\,
            I => \N__47690\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__47694\,
            I => \N__47685\
        );

    \I__9993\ : CascadeMux
    port map (
            O => \N__47693\,
            I => \N__47681\
        );

    \I__9992\ : Span4Mux_h
    port map (
            O => \N__47690\,
            I => \N__47678\
        );

    \I__9991\ : CascadeMux
    port map (
            O => \N__47689\,
            I => \N__47675\
        );

    \I__9990\ : CascadeMux
    port map (
            O => \N__47688\,
            I => \N__47672\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__47685\,
            I => \N__47669\
        );

    \I__9988\ : InMux
    port map (
            O => \N__47684\,
            I => \N__47664\
        );

    \I__9987\ : InMux
    port map (
            O => \N__47681\,
            I => \N__47664\
        );

    \I__9986\ : Span4Mux_v
    port map (
            O => \N__47678\,
            I => \N__47661\
        );

    \I__9985\ : InMux
    port map (
            O => \N__47675\,
            I => \N__47656\
        );

    \I__9984\ : InMux
    port map (
            O => \N__47672\,
            I => \N__47656\
        );

    \I__9983\ : Span4Mux_v
    port map (
            O => \N__47669\,
            I => \N__47651\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__47664\,
            I => \N__47651\
        );

    \I__9981\ : Odrv4
    port map (
            O => \N__47661\,
            I => data_in_frame_1_1
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__47656\,
            I => data_in_frame_1_1
        );

    \I__9979\ : Odrv4
    port map (
            O => \N__47651\,
            I => data_in_frame_1_1
        );

    \I__9978\ : InMux
    port map (
            O => \N__47644\,
            I => \N__47641\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__47641\,
            I => \N__47637\
        );

    \I__9976\ : InMux
    port map (
            O => \N__47640\,
            I => \N__47634\
        );

    \I__9975\ : Span4Mux_v
    port map (
            O => \N__47637\,
            I => \N__47628\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__47634\,
            I => \N__47625\
        );

    \I__9973\ : InMux
    port map (
            O => \N__47633\,
            I => \N__47620\
        );

    \I__9972\ : InMux
    port map (
            O => \N__47632\,
            I => \N__47617\
        );

    \I__9971\ : InMux
    port map (
            O => \N__47631\,
            I => \N__47612\
        );

    \I__9970\ : Span4Mux_v
    port map (
            O => \N__47628\,
            I => \N__47607\
        );

    \I__9969\ : Span4Mux_h
    port map (
            O => \N__47625\,
            I => \N__47607\
        );

    \I__9968\ : InMux
    port map (
            O => \N__47624\,
            I => \N__47604\
        );

    \I__9967\ : InMux
    port map (
            O => \N__47623\,
            I => \N__47601\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__47620\,
            I => \N__47596\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__47617\,
            I => \N__47596\
        );

    \I__9964\ : InMux
    port map (
            O => \N__47616\,
            I => \N__47591\
        );

    \I__9963\ : InMux
    port map (
            O => \N__47615\,
            I => \N__47591\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__47612\,
            I => data_in_frame_1_5
        );

    \I__9961\ : Odrv4
    port map (
            O => \N__47607\,
            I => data_in_frame_1_5
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__47604\,
            I => data_in_frame_1_5
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__47601\,
            I => data_in_frame_1_5
        );

    \I__9958\ : Odrv4
    port map (
            O => \N__47596\,
            I => data_in_frame_1_5
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__47591\,
            I => data_in_frame_1_5
        );

    \I__9956\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47575\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__47575\,
            I => \N__47572\
        );

    \I__9954\ : Span4Mux_h
    port map (
            O => \N__47572\,
            I => \N__47569\
        );

    \I__9953\ : Odrv4
    port map (
            O => \N__47569\,
            I => \c0.n21986\
        );

    \I__9952\ : CascadeMux
    port map (
            O => \N__47566\,
            I => \c0.n13848_cascade_\
        );

    \I__9951\ : InMux
    port map (
            O => \N__47563\,
            I => \N__47560\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__47560\,
            I => \N__47557\
        );

    \I__9949\ : Span4Mux_h
    port map (
            O => \N__47557\,
            I => \N__47554\
        );

    \I__9948\ : Span4Mux_v
    port map (
            O => \N__47554\,
            I => \N__47551\
        );

    \I__9947\ : Odrv4
    port map (
            O => \N__47551\,
            I => \c0.n13_adj_4405\
        );

    \I__9946\ : InMux
    port map (
            O => \N__47548\,
            I => \N__47544\
        );

    \I__9945\ : CascadeMux
    port map (
            O => \N__47547\,
            I => \N__47541\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__47544\,
            I => \N__47536\
        );

    \I__9943\ : InMux
    port map (
            O => \N__47541\,
            I => \N__47529\
        );

    \I__9942\ : InMux
    port map (
            O => \N__47540\,
            I => \N__47529\
        );

    \I__9941\ : InMux
    port map (
            O => \N__47539\,
            I => \N__47529\
        );

    \I__9940\ : Odrv4
    port map (
            O => \N__47536\,
            I => \c0.data_in_frame_2_7\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__47529\,
            I => \c0.data_in_frame_2_7\
        );

    \I__9938\ : CascadeMux
    port map (
            O => \N__47524\,
            I => \N__47519\
        );

    \I__9937\ : CascadeMux
    port map (
            O => \N__47523\,
            I => \N__47516\
        );

    \I__9936\ : CascadeMux
    port map (
            O => \N__47522\,
            I => \N__47513\
        );

    \I__9935\ : InMux
    port map (
            O => \N__47519\,
            I => \N__47510\
        );

    \I__9934\ : InMux
    port map (
            O => \N__47516\,
            I => \N__47505\
        );

    \I__9933\ : InMux
    port map (
            O => \N__47513\,
            I => \N__47502\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__47510\,
            I => \N__47497\
        );

    \I__9931\ : InMux
    port map (
            O => \N__47509\,
            I => \N__47494\
        );

    \I__9930\ : CascadeMux
    port map (
            O => \N__47508\,
            I => \N__47490\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__47505\,
            I => \N__47487\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__47502\,
            I => \N__47484\
        );

    \I__9927\ : InMux
    port map (
            O => \N__47501\,
            I => \N__47479\
        );

    \I__9926\ : InMux
    port map (
            O => \N__47500\,
            I => \N__47479\
        );

    \I__9925\ : Span4Mux_h
    port map (
            O => \N__47497\,
            I => \N__47476\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__47494\,
            I => \N__47473\
        );

    \I__9923\ : InMux
    port map (
            O => \N__47493\,
            I => \N__47468\
        );

    \I__9922\ : InMux
    port map (
            O => \N__47490\,
            I => \N__47468\
        );

    \I__9921\ : Odrv4
    port map (
            O => \N__47487\,
            I => \c0.data_in_frame_0_7\
        );

    \I__9920\ : Odrv4
    port map (
            O => \N__47484\,
            I => \c0.data_in_frame_0_7\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__47479\,
            I => \c0.data_in_frame_0_7\
        );

    \I__9918\ : Odrv4
    port map (
            O => \N__47476\,
            I => \c0.data_in_frame_0_7\
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__47473\,
            I => \c0.data_in_frame_0_7\
        );

    \I__9916\ : LocalMux
    port map (
            O => \N__47468\,
            I => \c0.data_in_frame_0_7\
        );

    \I__9915\ : InMux
    port map (
            O => \N__47455\,
            I => \N__47451\
        );

    \I__9914\ : InMux
    port map (
            O => \N__47454\,
            I => \N__47447\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__47451\,
            I => \N__47443\
        );

    \I__9912\ : InMux
    port map (
            O => \N__47450\,
            I => \N__47440\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__47447\,
            I => \N__47437\
        );

    \I__9910\ : InMux
    port map (
            O => \N__47446\,
            I => \N__47434\
        );

    \I__9909\ : Span4Mux_v
    port map (
            O => \N__47443\,
            I => \N__47431\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__47440\,
            I => \c0.data_in_frame_8_4\
        );

    \I__9907\ : Odrv4
    port map (
            O => \N__47437\,
            I => \c0.data_in_frame_8_4\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__47434\,
            I => \c0.data_in_frame_8_4\
        );

    \I__9905\ : Odrv4
    port map (
            O => \N__47431\,
            I => \c0.data_in_frame_8_4\
        );

    \I__9904\ : CascadeMux
    port map (
            O => \N__47422\,
            I => \c0.n21861_cascade_\
        );

    \I__9903\ : InMux
    port map (
            O => \N__47419\,
            I => \N__47416\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__47416\,
            I => \c0.n6_adj_4258\
        );

    \I__9901\ : SRMux
    port map (
            O => \N__47413\,
            I => \N__47410\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__47410\,
            I => \N__47407\
        );

    \I__9899\ : Span4Mux_s2_v
    port map (
            O => \N__47407\,
            I => \N__47404\
        );

    \I__9898\ : Odrv4
    port map (
            O => \N__47404\,
            I => \c0.n3_adj_4474\
        );

    \I__9897\ : CascadeMux
    port map (
            O => \N__47401\,
            I => \N__47398\
        );

    \I__9896\ : InMux
    port map (
            O => \N__47398\,
            I => \N__47395\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__47395\,
            I => \N__47392\
        );

    \I__9894\ : Span4Mux_v
    port map (
            O => \N__47392\,
            I => \N__47388\
        );

    \I__9893\ : CascadeMux
    port map (
            O => \N__47391\,
            I => \N__47385\
        );

    \I__9892\ : Span4Mux_v
    port map (
            O => \N__47388\,
            I => \N__47381\
        );

    \I__9891\ : InMux
    port map (
            O => \N__47385\,
            I => \N__47377\
        );

    \I__9890\ : InMux
    port map (
            O => \N__47384\,
            I => \N__47374\
        );

    \I__9889\ : Span4Mux_h
    port map (
            O => \N__47381\,
            I => \N__47371\
        );

    \I__9888\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47368\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__47377\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__47374\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__9885\ : Odrv4
    port map (
            O => \N__47371\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__47368\,
            I => \c0.FRAME_MATCHER_i_5\
        );

    \I__9883\ : CascadeMux
    port map (
            O => \N__47359\,
            I => \N__47356\
        );

    \I__9882\ : InMux
    port map (
            O => \N__47356\,
            I => \N__47352\
        );

    \I__9881\ : InMux
    port map (
            O => \N__47355\,
            I => \N__47349\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__47352\,
            I => \N__47342\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__47349\,
            I => \N__47342\
        );

    \I__9878\ : InMux
    port map (
            O => \N__47348\,
            I => \N__47339\
        );

    \I__9877\ : InMux
    port map (
            O => \N__47347\,
            I => \N__47336\
        );

    \I__9876\ : Span4Mux_v
    port map (
            O => \N__47342\,
            I => \N__47333\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__47339\,
            I => \N__47326\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__47336\,
            I => \N__47326\
        );

    \I__9873\ : Span4Mux_v
    port map (
            O => \N__47333\,
            I => \N__47326\
        );

    \I__9872\ : Odrv4
    port map (
            O => \N__47326\,
            I => \c0.FRAME_MATCHER_i_6\
        );

    \I__9871\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47317\
        );

    \I__9870\ : CascadeMux
    port map (
            O => \N__47322\,
            I => \N__47314\
        );

    \I__9869\ : CascadeMux
    port map (
            O => \N__47321\,
            I => \N__47311\
        );

    \I__9868\ : InMux
    port map (
            O => \N__47320\,
            I => \N__47308\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__47317\,
            I => \N__47305\
        );

    \I__9866\ : InMux
    port map (
            O => \N__47314\,
            I => \N__47300\
        );

    \I__9865\ : InMux
    port map (
            O => \N__47311\,
            I => \N__47300\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__47308\,
            I => \N__47297\
        );

    \I__9863\ : Span4Mux_h
    port map (
            O => \N__47305\,
            I => \N__47294\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__47300\,
            I => \N__47291\
        );

    \I__9861\ : Span4Mux_h
    port map (
            O => \N__47297\,
            I => \N__47288\
        );

    \I__9860\ : Span4Mux_h
    port map (
            O => \N__47294\,
            I => \N__47283\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__47291\,
            I => \N__47283\
        );

    \I__9858\ : Span4Mux_v
    port map (
            O => \N__47288\,
            I => \N__47280\
        );

    \I__9857\ : Span4Mux_v
    port map (
            O => \N__47283\,
            I => \N__47277\
        );

    \I__9856\ : Span4Mux_v
    port map (
            O => \N__47280\,
            I => \N__47274\
        );

    \I__9855\ : Span4Mux_v
    port map (
            O => \N__47277\,
            I => \N__47271\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__47274\,
            I => \c0.n11_adj_4326\
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__47271\,
            I => \c0.n11_adj_4326\
        );

    \I__9852\ : InMux
    port map (
            O => \N__47266\,
            I => \N__47263\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__47263\,
            I => \N__47260\
        );

    \I__9850\ : Span4Mux_h
    port map (
            O => \N__47260\,
            I => \N__47257\
        );

    \I__9849\ : Odrv4
    port map (
            O => \N__47257\,
            I => \c0.n10_adj_4399\
        );

    \I__9848\ : InMux
    port map (
            O => \N__47254\,
            I => \N__47250\
        );

    \I__9847\ : InMux
    port map (
            O => \N__47253\,
            I => \N__47247\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__47250\,
            I => \N__47243\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__47247\,
            I => \N__47240\
        );

    \I__9844\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47236\
        );

    \I__9843\ : Span4Mux_h
    port map (
            O => \N__47243\,
            I => \N__47233\
        );

    \I__9842\ : Span4Mux_h
    port map (
            O => \N__47240\,
            I => \N__47230\
        );

    \I__9841\ : InMux
    port map (
            O => \N__47239\,
            I => \N__47227\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__47236\,
            I => \c0.n13033\
        );

    \I__9839\ : Odrv4
    port map (
            O => \N__47233\,
            I => \c0.n13033\
        );

    \I__9838\ : Odrv4
    port map (
            O => \N__47230\,
            I => \c0.n13033\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__47227\,
            I => \c0.n13033\
        );

    \I__9836\ : IoInMux
    port map (
            O => \N__47218\,
            I => \N__47203\
        );

    \I__9835\ : CascadeMux
    port map (
            O => \N__47217\,
            I => \N__47199\
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__47216\,
            I => \N__47195\
        );

    \I__9833\ : CascadeMux
    port map (
            O => \N__47215\,
            I => \N__47191\
        );

    \I__9832\ : CascadeMux
    port map (
            O => \N__47214\,
            I => \N__47186\
        );

    \I__9831\ : CascadeMux
    port map (
            O => \N__47213\,
            I => \N__47182\
        );

    \I__9830\ : CascadeMux
    port map (
            O => \N__47212\,
            I => \N__47178\
        );

    \I__9829\ : CascadeMux
    port map (
            O => \N__47211\,
            I => \N__47173\
        );

    \I__9828\ : CascadeMux
    port map (
            O => \N__47210\,
            I => \N__47169\
        );

    \I__9827\ : CascadeMux
    port map (
            O => \N__47209\,
            I => \N__47165\
        );

    \I__9826\ : CascadeMux
    port map (
            O => \N__47208\,
            I => \N__47160\
        );

    \I__9825\ : CascadeMux
    port map (
            O => \N__47207\,
            I => \N__47156\
        );

    \I__9824\ : CascadeMux
    port map (
            O => \N__47206\,
            I => \N__47152\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__47203\,
            I => \N__47136\
        );

    \I__9822\ : InMux
    port map (
            O => \N__47202\,
            I => \N__47121\
        );

    \I__9821\ : InMux
    port map (
            O => \N__47199\,
            I => \N__47121\
        );

    \I__9820\ : InMux
    port map (
            O => \N__47198\,
            I => \N__47121\
        );

    \I__9819\ : InMux
    port map (
            O => \N__47195\,
            I => \N__47121\
        );

    \I__9818\ : InMux
    port map (
            O => \N__47194\,
            I => \N__47121\
        );

    \I__9817\ : InMux
    port map (
            O => \N__47191\,
            I => \N__47121\
        );

    \I__9816\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47121\
        );

    \I__9815\ : InMux
    port map (
            O => \N__47189\,
            I => \N__47106\
        );

    \I__9814\ : InMux
    port map (
            O => \N__47186\,
            I => \N__47106\
        );

    \I__9813\ : InMux
    port map (
            O => \N__47185\,
            I => \N__47106\
        );

    \I__9812\ : InMux
    port map (
            O => \N__47182\,
            I => \N__47106\
        );

    \I__9811\ : InMux
    port map (
            O => \N__47181\,
            I => \N__47106\
        );

    \I__9810\ : InMux
    port map (
            O => \N__47178\,
            I => \N__47106\
        );

    \I__9809\ : InMux
    port map (
            O => \N__47177\,
            I => \N__47106\
        );

    \I__9808\ : InMux
    port map (
            O => \N__47176\,
            I => \N__47091\
        );

    \I__9807\ : InMux
    port map (
            O => \N__47173\,
            I => \N__47091\
        );

    \I__9806\ : InMux
    port map (
            O => \N__47172\,
            I => \N__47091\
        );

    \I__9805\ : InMux
    port map (
            O => \N__47169\,
            I => \N__47091\
        );

    \I__9804\ : InMux
    port map (
            O => \N__47168\,
            I => \N__47091\
        );

    \I__9803\ : InMux
    port map (
            O => \N__47165\,
            I => \N__47091\
        );

    \I__9802\ : InMux
    port map (
            O => \N__47164\,
            I => \N__47091\
        );

    \I__9801\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47076\
        );

    \I__9800\ : InMux
    port map (
            O => \N__47160\,
            I => \N__47076\
        );

    \I__9799\ : InMux
    port map (
            O => \N__47159\,
            I => \N__47076\
        );

    \I__9798\ : InMux
    port map (
            O => \N__47156\,
            I => \N__47076\
        );

    \I__9797\ : InMux
    port map (
            O => \N__47155\,
            I => \N__47076\
        );

    \I__9796\ : InMux
    port map (
            O => \N__47152\,
            I => \N__47076\
        );

    \I__9795\ : InMux
    port map (
            O => \N__47151\,
            I => \N__47076\
        );

    \I__9794\ : CascadeMux
    port map (
            O => \N__47150\,
            I => \N__47072\
        );

    \I__9793\ : CascadeMux
    port map (
            O => \N__47149\,
            I => \N__47068\
        );

    \I__9792\ : CascadeMux
    port map (
            O => \N__47148\,
            I => \N__47064\
        );

    \I__9791\ : CascadeMux
    port map (
            O => \N__47147\,
            I => \N__47059\
        );

    \I__9790\ : CascadeMux
    port map (
            O => \N__47146\,
            I => \N__47055\
        );

    \I__9789\ : CascadeMux
    port map (
            O => \N__47145\,
            I => \N__47051\
        );

    \I__9788\ : CascadeMux
    port map (
            O => \N__47144\,
            I => \N__47046\
        );

    \I__9787\ : CascadeMux
    port map (
            O => \N__47143\,
            I => \N__47042\
        );

    \I__9786\ : CascadeMux
    port map (
            O => \N__47142\,
            I => \N__47038\
        );

    \I__9785\ : CascadeMux
    port map (
            O => \N__47141\,
            I => \N__47033\
        );

    \I__9784\ : CascadeMux
    port map (
            O => \N__47140\,
            I => \N__47029\
        );

    \I__9783\ : CascadeMux
    port map (
            O => \N__47139\,
            I => \N__47025\
        );

    \I__9782\ : IoSpan4Mux
    port map (
            O => \N__47136\,
            I => \N__47003\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__47121\,
            I => \N__47003\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__47106\,
            I => \N__47003\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__47091\,
            I => \N__47003\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__47076\,
            I => \N__47000\
        );

    \I__9777\ : InMux
    port map (
            O => \N__47075\,
            I => \N__46985\
        );

    \I__9776\ : InMux
    port map (
            O => \N__47072\,
            I => \N__46985\
        );

    \I__9775\ : InMux
    port map (
            O => \N__47071\,
            I => \N__46985\
        );

    \I__9774\ : InMux
    port map (
            O => \N__47068\,
            I => \N__46985\
        );

    \I__9773\ : InMux
    port map (
            O => \N__47067\,
            I => \N__46985\
        );

    \I__9772\ : InMux
    port map (
            O => \N__47064\,
            I => \N__46985\
        );

    \I__9771\ : InMux
    port map (
            O => \N__47063\,
            I => \N__46985\
        );

    \I__9770\ : InMux
    port map (
            O => \N__47062\,
            I => \N__46970\
        );

    \I__9769\ : InMux
    port map (
            O => \N__47059\,
            I => \N__46970\
        );

    \I__9768\ : InMux
    port map (
            O => \N__47058\,
            I => \N__46970\
        );

    \I__9767\ : InMux
    port map (
            O => \N__47055\,
            I => \N__46970\
        );

    \I__9766\ : InMux
    port map (
            O => \N__47054\,
            I => \N__46970\
        );

    \I__9765\ : InMux
    port map (
            O => \N__47051\,
            I => \N__46970\
        );

    \I__9764\ : InMux
    port map (
            O => \N__47050\,
            I => \N__46970\
        );

    \I__9763\ : InMux
    port map (
            O => \N__47049\,
            I => \N__46955\
        );

    \I__9762\ : InMux
    port map (
            O => \N__47046\,
            I => \N__46955\
        );

    \I__9761\ : InMux
    port map (
            O => \N__47045\,
            I => \N__46955\
        );

    \I__9760\ : InMux
    port map (
            O => \N__47042\,
            I => \N__46955\
        );

    \I__9759\ : InMux
    port map (
            O => \N__47041\,
            I => \N__46955\
        );

    \I__9758\ : InMux
    port map (
            O => \N__47038\,
            I => \N__46955\
        );

    \I__9757\ : InMux
    port map (
            O => \N__47037\,
            I => \N__46955\
        );

    \I__9756\ : InMux
    port map (
            O => \N__47036\,
            I => \N__46940\
        );

    \I__9755\ : InMux
    port map (
            O => \N__47033\,
            I => \N__46940\
        );

    \I__9754\ : InMux
    port map (
            O => \N__47032\,
            I => \N__46940\
        );

    \I__9753\ : InMux
    port map (
            O => \N__47029\,
            I => \N__46940\
        );

    \I__9752\ : InMux
    port map (
            O => \N__47028\,
            I => \N__46940\
        );

    \I__9751\ : InMux
    port map (
            O => \N__47025\,
            I => \N__46940\
        );

    \I__9750\ : InMux
    port map (
            O => \N__47024\,
            I => \N__46940\
        );

    \I__9749\ : CascadeMux
    port map (
            O => \N__47023\,
            I => \N__46936\
        );

    \I__9748\ : CascadeMux
    port map (
            O => \N__47022\,
            I => \N__46932\
        );

    \I__9747\ : CascadeMux
    port map (
            O => \N__47021\,
            I => \N__46928\
        );

    \I__9746\ : CascadeMux
    port map (
            O => \N__47020\,
            I => \N__46923\
        );

    \I__9745\ : CascadeMux
    port map (
            O => \N__47019\,
            I => \N__46919\
        );

    \I__9744\ : CascadeMux
    port map (
            O => \N__47018\,
            I => \N__46915\
        );

    \I__9743\ : CascadeMux
    port map (
            O => \N__47017\,
            I => \N__46910\
        );

    \I__9742\ : CascadeMux
    port map (
            O => \N__47016\,
            I => \N__46906\
        );

    \I__9741\ : CascadeMux
    port map (
            O => \N__47015\,
            I => \N__46902\
        );

    \I__9740\ : CascadeMux
    port map (
            O => \N__47014\,
            I => \N__46897\
        );

    \I__9739\ : CascadeMux
    port map (
            O => \N__47013\,
            I => \N__46893\
        );

    \I__9738\ : CascadeMux
    port map (
            O => \N__47012\,
            I => \N__46889\
        );

    \I__9737\ : Span4Mux_s3_v
    port map (
            O => \N__47003\,
            I => \N__46865\
        );

    \I__9736\ : Span4Mux_h
    port map (
            O => \N__47000\,
            I => \N__46865\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__46985\,
            I => \N__46865\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__46970\,
            I => \N__46865\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__46955\,
            I => \N__46865\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__46940\,
            I => \N__46862\
        );

    \I__9731\ : InMux
    port map (
            O => \N__46939\,
            I => \N__46847\
        );

    \I__9730\ : InMux
    port map (
            O => \N__46936\,
            I => \N__46847\
        );

    \I__9729\ : InMux
    port map (
            O => \N__46935\,
            I => \N__46847\
        );

    \I__9728\ : InMux
    port map (
            O => \N__46932\,
            I => \N__46847\
        );

    \I__9727\ : InMux
    port map (
            O => \N__46931\,
            I => \N__46847\
        );

    \I__9726\ : InMux
    port map (
            O => \N__46928\,
            I => \N__46847\
        );

    \I__9725\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46847\
        );

    \I__9724\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46832\
        );

    \I__9723\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46832\
        );

    \I__9722\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46832\
        );

    \I__9721\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46832\
        );

    \I__9720\ : InMux
    port map (
            O => \N__46918\,
            I => \N__46832\
        );

    \I__9719\ : InMux
    port map (
            O => \N__46915\,
            I => \N__46832\
        );

    \I__9718\ : InMux
    port map (
            O => \N__46914\,
            I => \N__46832\
        );

    \I__9717\ : InMux
    port map (
            O => \N__46913\,
            I => \N__46817\
        );

    \I__9716\ : InMux
    port map (
            O => \N__46910\,
            I => \N__46817\
        );

    \I__9715\ : InMux
    port map (
            O => \N__46909\,
            I => \N__46817\
        );

    \I__9714\ : InMux
    port map (
            O => \N__46906\,
            I => \N__46817\
        );

    \I__9713\ : InMux
    port map (
            O => \N__46905\,
            I => \N__46817\
        );

    \I__9712\ : InMux
    port map (
            O => \N__46902\,
            I => \N__46817\
        );

    \I__9711\ : InMux
    port map (
            O => \N__46901\,
            I => \N__46817\
        );

    \I__9710\ : InMux
    port map (
            O => \N__46900\,
            I => \N__46802\
        );

    \I__9709\ : InMux
    port map (
            O => \N__46897\,
            I => \N__46802\
        );

    \I__9708\ : InMux
    port map (
            O => \N__46896\,
            I => \N__46802\
        );

    \I__9707\ : InMux
    port map (
            O => \N__46893\,
            I => \N__46802\
        );

    \I__9706\ : InMux
    port map (
            O => \N__46892\,
            I => \N__46802\
        );

    \I__9705\ : InMux
    port map (
            O => \N__46889\,
            I => \N__46802\
        );

    \I__9704\ : InMux
    port map (
            O => \N__46888\,
            I => \N__46802\
        );

    \I__9703\ : CascadeMux
    port map (
            O => \N__46887\,
            I => \N__46798\
        );

    \I__9702\ : CascadeMux
    port map (
            O => \N__46886\,
            I => \N__46794\
        );

    \I__9701\ : CascadeMux
    port map (
            O => \N__46885\,
            I => \N__46790\
        );

    \I__9700\ : CascadeMux
    port map (
            O => \N__46884\,
            I => \N__46785\
        );

    \I__9699\ : CascadeMux
    port map (
            O => \N__46883\,
            I => \N__46781\
        );

    \I__9698\ : CascadeMux
    port map (
            O => \N__46882\,
            I => \N__46777\
        );

    \I__9697\ : CascadeMux
    port map (
            O => \N__46881\,
            I => \N__46772\
        );

    \I__9696\ : CascadeMux
    port map (
            O => \N__46880\,
            I => \N__46768\
        );

    \I__9695\ : CascadeMux
    port map (
            O => \N__46879\,
            I => \N__46764\
        );

    \I__9694\ : CascadeMux
    port map (
            O => \N__46878\,
            I => \N__46759\
        );

    \I__9693\ : CascadeMux
    port map (
            O => \N__46877\,
            I => \N__46755\
        );

    \I__9692\ : CascadeMux
    port map (
            O => \N__46876\,
            I => \N__46751\
        );

    \I__9691\ : Span4Mux_v
    port map (
            O => \N__46865\,
            I => \N__46730\
        );

    \I__9690\ : Span4Mux_h
    port map (
            O => \N__46862\,
            I => \N__46730\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__46847\,
            I => \N__46730\
        );

    \I__9688\ : LocalMux
    port map (
            O => \N__46832\,
            I => \N__46730\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__46817\,
            I => \N__46730\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__46802\,
            I => \N__46727\
        );

    \I__9685\ : InMux
    port map (
            O => \N__46801\,
            I => \N__46712\
        );

    \I__9684\ : InMux
    port map (
            O => \N__46798\,
            I => \N__46712\
        );

    \I__9683\ : InMux
    port map (
            O => \N__46797\,
            I => \N__46712\
        );

    \I__9682\ : InMux
    port map (
            O => \N__46794\,
            I => \N__46712\
        );

    \I__9681\ : InMux
    port map (
            O => \N__46793\,
            I => \N__46712\
        );

    \I__9680\ : InMux
    port map (
            O => \N__46790\,
            I => \N__46712\
        );

    \I__9679\ : InMux
    port map (
            O => \N__46789\,
            I => \N__46712\
        );

    \I__9678\ : InMux
    port map (
            O => \N__46788\,
            I => \N__46697\
        );

    \I__9677\ : InMux
    port map (
            O => \N__46785\,
            I => \N__46697\
        );

    \I__9676\ : InMux
    port map (
            O => \N__46784\,
            I => \N__46697\
        );

    \I__9675\ : InMux
    port map (
            O => \N__46781\,
            I => \N__46697\
        );

    \I__9674\ : InMux
    port map (
            O => \N__46780\,
            I => \N__46697\
        );

    \I__9673\ : InMux
    port map (
            O => \N__46777\,
            I => \N__46697\
        );

    \I__9672\ : InMux
    port map (
            O => \N__46776\,
            I => \N__46697\
        );

    \I__9671\ : InMux
    port map (
            O => \N__46775\,
            I => \N__46682\
        );

    \I__9670\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46682\
        );

    \I__9669\ : InMux
    port map (
            O => \N__46771\,
            I => \N__46682\
        );

    \I__9668\ : InMux
    port map (
            O => \N__46768\,
            I => \N__46682\
        );

    \I__9667\ : InMux
    port map (
            O => \N__46767\,
            I => \N__46682\
        );

    \I__9666\ : InMux
    port map (
            O => \N__46764\,
            I => \N__46682\
        );

    \I__9665\ : InMux
    port map (
            O => \N__46763\,
            I => \N__46682\
        );

    \I__9664\ : InMux
    port map (
            O => \N__46762\,
            I => \N__46667\
        );

    \I__9663\ : InMux
    port map (
            O => \N__46759\,
            I => \N__46667\
        );

    \I__9662\ : InMux
    port map (
            O => \N__46758\,
            I => \N__46667\
        );

    \I__9661\ : InMux
    port map (
            O => \N__46755\,
            I => \N__46667\
        );

    \I__9660\ : InMux
    port map (
            O => \N__46754\,
            I => \N__46667\
        );

    \I__9659\ : InMux
    port map (
            O => \N__46751\,
            I => \N__46667\
        );

    \I__9658\ : InMux
    port map (
            O => \N__46750\,
            I => \N__46667\
        );

    \I__9657\ : CascadeMux
    port map (
            O => \N__46749\,
            I => \N__46663\
        );

    \I__9656\ : CascadeMux
    port map (
            O => \N__46748\,
            I => \N__46659\
        );

    \I__9655\ : CascadeMux
    port map (
            O => \N__46747\,
            I => \N__46655\
        );

    \I__9654\ : CascadeMux
    port map (
            O => \N__46746\,
            I => \N__46650\
        );

    \I__9653\ : CascadeMux
    port map (
            O => \N__46745\,
            I => \N__46646\
        );

    \I__9652\ : CascadeMux
    port map (
            O => \N__46744\,
            I => \N__46642\
        );

    \I__9651\ : CascadeMux
    port map (
            O => \N__46743\,
            I => \N__46637\
        );

    \I__9650\ : CascadeMux
    port map (
            O => \N__46742\,
            I => \N__46633\
        );

    \I__9649\ : CascadeMux
    port map (
            O => \N__46741\,
            I => \N__46629\
        );

    \I__9648\ : Span4Mux_v
    port map (
            O => \N__46730\,
            I => \N__46603\
        );

    \I__9647\ : Span4Mux_h
    port map (
            O => \N__46727\,
            I => \N__46603\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__46712\,
            I => \N__46603\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__46697\,
            I => \N__46603\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__46682\,
            I => \N__46603\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__46667\,
            I => \N__46603\
        );

    \I__9642\ : InMux
    port map (
            O => \N__46666\,
            I => \N__46588\
        );

    \I__9641\ : InMux
    port map (
            O => \N__46663\,
            I => \N__46588\
        );

    \I__9640\ : InMux
    port map (
            O => \N__46662\,
            I => \N__46588\
        );

    \I__9639\ : InMux
    port map (
            O => \N__46659\,
            I => \N__46588\
        );

    \I__9638\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46588\
        );

    \I__9637\ : InMux
    port map (
            O => \N__46655\,
            I => \N__46588\
        );

    \I__9636\ : InMux
    port map (
            O => \N__46654\,
            I => \N__46588\
        );

    \I__9635\ : InMux
    port map (
            O => \N__46653\,
            I => \N__46573\
        );

    \I__9634\ : InMux
    port map (
            O => \N__46650\,
            I => \N__46573\
        );

    \I__9633\ : InMux
    port map (
            O => \N__46649\,
            I => \N__46573\
        );

    \I__9632\ : InMux
    port map (
            O => \N__46646\,
            I => \N__46573\
        );

    \I__9631\ : InMux
    port map (
            O => \N__46645\,
            I => \N__46573\
        );

    \I__9630\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46573\
        );

    \I__9629\ : InMux
    port map (
            O => \N__46641\,
            I => \N__46573\
        );

    \I__9628\ : InMux
    port map (
            O => \N__46640\,
            I => \N__46558\
        );

    \I__9627\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46558\
        );

    \I__9626\ : InMux
    port map (
            O => \N__46636\,
            I => \N__46558\
        );

    \I__9625\ : InMux
    port map (
            O => \N__46633\,
            I => \N__46558\
        );

    \I__9624\ : InMux
    port map (
            O => \N__46632\,
            I => \N__46558\
        );

    \I__9623\ : InMux
    port map (
            O => \N__46629\,
            I => \N__46558\
        );

    \I__9622\ : InMux
    port map (
            O => \N__46628\,
            I => \N__46558\
        );

    \I__9621\ : CascadeMux
    port map (
            O => \N__46627\,
            I => \N__46554\
        );

    \I__9620\ : CascadeMux
    port map (
            O => \N__46626\,
            I => \N__46550\
        );

    \I__9619\ : CascadeMux
    port map (
            O => \N__46625\,
            I => \N__46546\
        );

    \I__9618\ : CascadeMux
    port map (
            O => \N__46624\,
            I => \N__46541\
        );

    \I__9617\ : CascadeMux
    port map (
            O => \N__46623\,
            I => \N__46537\
        );

    \I__9616\ : CascadeMux
    port map (
            O => \N__46622\,
            I => \N__46533\
        );

    \I__9615\ : CascadeMux
    port map (
            O => \N__46621\,
            I => \N__46504\
        );

    \I__9614\ : CascadeMux
    port map (
            O => \N__46620\,
            I => \N__46500\
        );

    \I__9613\ : CascadeMux
    port map (
            O => \N__46619\,
            I => \N__46496\
        );

    \I__9612\ : CascadeMux
    port map (
            O => \N__46618\,
            I => \N__46488\
        );

    \I__9611\ : CascadeMux
    port map (
            O => \N__46617\,
            I => \N__46484\
        );

    \I__9610\ : CascadeMux
    port map (
            O => \N__46616\,
            I => \N__46480\
        );

    \I__9609\ : Span4Mux_v
    port map (
            O => \N__46603\,
            I => \N__46470\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__46588\,
            I => \N__46470\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__46573\,
            I => \N__46470\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__46558\,
            I => \N__46470\
        );

    \I__9605\ : InMux
    port map (
            O => \N__46557\,
            I => \N__46455\
        );

    \I__9604\ : InMux
    port map (
            O => \N__46554\,
            I => \N__46455\
        );

    \I__9603\ : InMux
    port map (
            O => \N__46553\,
            I => \N__46455\
        );

    \I__9602\ : InMux
    port map (
            O => \N__46550\,
            I => \N__46455\
        );

    \I__9601\ : InMux
    port map (
            O => \N__46549\,
            I => \N__46455\
        );

    \I__9600\ : InMux
    port map (
            O => \N__46546\,
            I => \N__46455\
        );

    \I__9599\ : InMux
    port map (
            O => \N__46545\,
            I => \N__46455\
        );

    \I__9598\ : InMux
    port map (
            O => \N__46544\,
            I => \N__46440\
        );

    \I__9597\ : InMux
    port map (
            O => \N__46541\,
            I => \N__46440\
        );

    \I__9596\ : InMux
    port map (
            O => \N__46540\,
            I => \N__46440\
        );

    \I__9595\ : InMux
    port map (
            O => \N__46537\,
            I => \N__46440\
        );

    \I__9594\ : InMux
    port map (
            O => \N__46536\,
            I => \N__46440\
        );

    \I__9593\ : InMux
    port map (
            O => \N__46533\,
            I => \N__46440\
        );

    \I__9592\ : InMux
    port map (
            O => \N__46532\,
            I => \N__46440\
        );

    \I__9591\ : InMux
    port map (
            O => \N__46531\,
            I => \N__46433\
        );

    \I__9590\ : InMux
    port map (
            O => \N__46530\,
            I => \N__46433\
        );

    \I__9589\ : InMux
    port map (
            O => \N__46529\,
            I => \N__46433\
        );

    \I__9588\ : InMux
    port map (
            O => \N__46528\,
            I => \N__46424\
        );

    \I__9587\ : InMux
    port map (
            O => \N__46527\,
            I => \N__46424\
        );

    \I__9586\ : InMux
    port map (
            O => \N__46526\,
            I => \N__46424\
        );

    \I__9585\ : InMux
    port map (
            O => \N__46525\,
            I => \N__46424\
        );

    \I__9584\ : InMux
    port map (
            O => \N__46524\,
            I => \N__46417\
        );

    \I__9583\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46417\
        );

    \I__9582\ : InMux
    port map (
            O => \N__46522\,
            I => \N__46417\
        );

    \I__9581\ : InMux
    port map (
            O => \N__46521\,
            I => \N__46408\
        );

    \I__9580\ : InMux
    port map (
            O => \N__46520\,
            I => \N__46408\
        );

    \I__9579\ : InMux
    port map (
            O => \N__46519\,
            I => \N__46408\
        );

    \I__9578\ : InMux
    port map (
            O => \N__46518\,
            I => \N__46408\
        );

    \I__9577\ : InMux
    port map (
            O => \N__46517\,
            I => \N__46401\
        );

    \I__9576\ : InMux
    port map (
            O => \N__46516\,
            I => \N__46401\
        );

    \I__9575\ : InMux
    port map (
            O => \N__46515\,
            I => \N__46401\
        );

    \I__9574\ : InMux
    port map (
            O => \N__46514\,
            I => \N__46392\
        );

    \I__9573\ : InMux
    port map (
            O => \N__46513\,
            I => \N__46392\
        );

    \I__9572\ : InMux
    port map (
            O => \N__46512\,
            I => \N__46392\
        );

    \I__9571\ : InMux
    port map (
            O => \N__46511\,
            I => \N__46392\
        );

    \I__9570\ : CascadeMux
    port map (
            O => \N__46510\,
            I => \N__46388\
        );

    \I__9569\ : CascadeMux
    port map (
            O => \N__46509\,
            I => \N__46384\
        );

    \I__9568\ : CascadeMux
    port map (
            O => \N__46508\,
            I => \N__46380\
        );

    \I__9567\ : InMux
    port map (
            O => \N__46507\,
            I => \N__46364\
        );

    \I__9566\ : InMux
    port map (
            O => \N__46504\,
            I => \N__46364\
        );

    \I__9565\ : InMux
    port map (
            O => \N__46503\,
            I => \N__46364\
        );

    \I__9564\ : InMux
    port map (
            O => \N__46500\,
            I => \N__46364\
        );

    \I__9563\ : InMux
    port map (
            O => \N__46499\,
            I => \N__46364\
        );

    \I__9562\ : InMux
    port map (
            O => \N__46496\,
            I => \N__46364\
        );

    \I__9561\ : InMux
    port map (
            O => \N__46495\,
            I => \N__46364\
        );

    \I__9560\ : CascadeMux
    port map (
            O => \N__46494\,
            I => \N__46360\
        );

    \I__9559\ : CascadeMux
    port map (
            O => \N__46493\,
            I => \N__46356\
        );

    \I__9558\ : CascadeMux
    port map (
            O => \N__46492\,
            I => \N__46352\
        );

    \I__9557\ : InMux
    port map (
            O => \N__46491\,
            I => \N__46336\
        );

    \I__9556\ : InMux
    port map (
            O => \N__46488\,
            I => \N__46336\
        );

    \I__9555\ : InMux
    port map (
            O => \N__46487\,
            I => \N__46336\
        );

    \I__9554\ : InMux
    port map (
            O => \N__46484\,
            I => \N__46336\
        );

    \I__9553\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46336\
        );

    \I__9552\ : InMux
    port map (
            O => \N__46480\,
            I => \N__46336\
        );

    \I__9551\ : InMux
    port map (
            O => \N__46479\,
            I => \N__46336\
        );

    \I__9550\ : Span4Mux_v
    port map (
            O => \N__46470\,
            I => \N__46329\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__46455\,
            I => \N__46329\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__46440\,
            I => \N__46329\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__46433\,
            I => \N__46316\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__46424\,
            I => \N__46316\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__46417\,
            I => \N__46316\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__46408\,
            I => \N__46316\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__46401\,
            I => \N__46316\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__46392\,
            I => \N__46316\
        );

    \I__9541\ : InMux
    port map (
            O => \N__46391\,
            I => \N__46301\
        );

    \I__9540\ : InMux
    port map (
            O => \N__46388\,
            I => \N__46301\
        );

    \I__9539\ : InMux
    port map (
            O => \N__46387\,
            I => \N__46301\
        );

    \I__9538\ : InMux
    port map (
            O => \N__46384\,
            I => \N__46301\
        );

    \I__9537\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46301\
        );

    \I__9536\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46301\
        );

    \I__9535\ : InMux
    port map (
            O => \N__46379\,
            I => \N__46301\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__46364\,
            I => \N__46298\
        );

    \I__9533\ : InMux
    port map (
            O => \N__46363\,
            I => \N__46283\
        );

    \I__9532\ : InMux
    port map (
            O => \N__46360\,
            I => \N__46283\
        );

    \I__9531\ : InMux
    port map (
            O => \N__46359\,
            I => \N__46283\
        );

    \I__9530\ : InMux
    port map (
            O => \N__46356\,
            I => \N__46283\
        );

    \I__9529\ : InMux
    port map (
            O => \N__46355\,
            I => \N__46283\
        );

    \I__9528\ : InMux
    port map (
            O => \N__46352\,
            I => \N__46283\
        );

    \I__9527\ : InMux
    port map (
            O => \N__46351\,
            I => \N__46283\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__46336\,
            I => \N__46259\
        );

    \I__9525\ : Span4Mux_v
    port map (
            O => \N__46329\,
            I => \N__46252\
        );

    \I__9524\ : Span4Mux_v
    port map (
            O => \N__46316\,
            I => \N__46252\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__46301\,
            I => \N__46252\
        );

    \I__9522\ : Span4Mux_v
    port map (
            O => \N__46298\,
            I => \N__46247\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__46283\,
            I => \N__46247\
        );

    \I__9520\ : InMux
    port map (
            O => \N__46282\,
            I => \N__46240\
        );

    \I__9519\ : InMux
    port map (
            O => \N__46281\,
            I => \N__46240\
        );

    \I__9518\ : InMux
    port map (
            O => \N__46280\,
            I => \N__46240\
        );

    \I__9517\ : InMux
    port map (
            O => \N__46279\,
            I => \N__46231\
        );

    \I__9516\ : InMux
    port map (
            O => \N__46278\,
            I => \N__46231\
        );

    \I__9515\ : InMux
    port map (
            O => \N__46277\,
            I => \N__46231\
        );

    \I__9514\ : InMux
    port map (
            O => \N__46276\,
            I => \N__46231\
        );

    \I__9513\ : InMux
    port map (
            O => \N__46275\,
            I => \N__46224\
        );

    \I__9512\ : InMux
    port map (
            O => \N__46274\,
            I => \N__46224\
        );

    \I__9511\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46224\
        );

    \I__9510\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46215\
        );

    \I__9509\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46215\
        );

    \I__9508\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46215\
        );

    \I__9507\ : InMux
    port map (
            O => \N__46269\,
            I => \N__46215\
        );

    \I__9506\ : InMux
    port map (
            O => \N__46268\,
            I => \N__46208\
        );

    \I__9505\ : InMux
    port map (
            O => \N__46267\,
            I => \N__46208\
        );

    \I__9504\ : InMux
    port map (
            O => \N__46266\,
            I => \N__46208\
        );

    \I__9503\ : InMux
    port map (
            O => \N__46265\,
            I => \N__46199\
        );

    \I__9502\ : InMux
    port map (
            O => \N__46264\,
            I => \N__46199\
        );

    \I__9501\ : InMux
    port map (
            O => \N__46263\,
            I => \N__46199\
        );

    \I__9500\ : InMux
    port map (
            O => \N__46262\,
            I => \N__46199\
        );

    \I__9499\ : Odrv4
    port map (
            O => \N__46259\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9498\ : Odrv4
    port map (
            O => \N__46252\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9497\ : Odrv4
    port map (
            O => \N__46247\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__46240\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__46231\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__46224\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__46215\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__46208\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__46199\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9490\ : InMux
    port map (
            O => \N__46180\,
            I => \bfn_19_32_0_\
        );

    \I__9489\ : CascadeMux
    port map (
            O => \N__46177\,
            I => \N__46171\
        );

    \I__9488\ : InMux
    port map (
            O => \N__46176\,
            I => \N__46168\
        );

    \I__9487\ : CascadeMux
    port map (
            O => \N__46175\,
            I => \N__46165\
        );

    \I__9486\ : CascadeMux
    port map (
            O => \N__46174\,
            I => \N__46162\
        );

    \I__9485\ : InMux
    port map (
            O => \N__46171\,
            I => \N__46159\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__46168\,
            I => \N__46155\
        );

    \I__9483\ : InMux
    port map (
            O => \N__46165\,
            I => \N__46152\
        );

    \I__9482\ : InMux
    port map (
            O => \N__46162\,
            I => \N__46149\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__46159\,
            I => \N__46144\
        );

    \I__9480\ : InMux
    port map (
            O => \N__46158\,
            I => \N__46141\
        );

    \I__9479\ : Span4Mux_v
    port map (
            O => \N__46155\,
            I => \N__46138\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__46152\,
            I => \N__46135\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__46149\,
            I => \N__46132\
        );

    \I__9476\ : InMux
    port map (
            O => \N__46148\,
            I => \N__46129\
        );

    \I__9475\ : InMux
    port map (
            O => \N__46147\,
            I => \N__46126\
        );

    \I__9474\ : Span4Mux_h
    port map (
            O => \N__46144\,
            I => \N__46121\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__46141\,
            I => \N__46121\
        );

    \I__9472\ : Span4Mux_h
    port map (
            O => \N__46138\,
            I => \N__46116\
        );

    \I__9471\ : Span4Mux_v
    port map (
            O => \N__46135\,
            I => \N__46116\
        );

    \I__9470\ : Span4Mux_h
    port map (
            O => \N__46132\,
            I => \N__46113\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__46129\,
            I => \N__46110\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__46126\,
            I => \N__46104\
        );

    \I__9467\ : Span4Mux_h
    port map (
            O => \N__46121\,
            I => \N__46104\
        );

    \I__9466\ : Span4Mux_h
    port map (
            O => \N__46116\,
            I => \N__46099\
        );

    \I__9465\ : Span4Mux_v
    port map (
            O => \N__46113\,
            I => \N__46099\
        );

    \I__9464\ : Span12Mux_h
    port map (
            O => \N__46110\,
            I => \N__46096\
        );

    \I__9463\ : InMux
    port map (
            O => \N__46109\,
            I => \N__46093\
        );

    \I__9462\ : Sp12to4
    port map (
            O => \N__46104\,
            I => \N__46090\
        );

    \I__9461\ : Span4Mux_v
    port map (
            O => \N__46099\,
            I => \N__46087\
        );

    \I__9460\ : Span12Mux_v
    port map (
            O => \N__46096\,
            I => \N__46084\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__46093\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__9458\ : Odrv12
    port map (
            O => \N__46090\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__46087\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__9456\ : Odrv12
    port map (
            O => \N__46084\,
            I => \c0.FRAME_MATCHER_i_31\
        );

    \I__9455\ : SRMux
    port map (
            O => \N__46075\,
            I => \N__46072\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__46072\,
            I => \N__46069\
        );

    \I__9453\ : Span4Mux_s1_v
    port map (
            O => \N__46069\,
            I => \N__46066\
        );

    \I__9452\ : Span4Mux_v
    port map (
            O => \N__46066\,
            I => \N__46063\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__46063\,
            I => \c0.n3_adj_4421\
        );

    \I__9450\ : SRMux
    port map (
            O => \N__46060\,
            I => \N__46057\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__46057\,
            I => \c0.n3_adj_4475\
        );

    \I__9448\ : InMux
    port map (
            O => \N__46054\,
            I => \N__46051\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__46051\,
            I => \N__46045\
        );

    \I__9446\ : InMux
    port map (
            O => \N__46050\,
            I => \N__46040\
        );

    \I__9445\ : InMux
    port map (
            O => \N__46049\,
            I => \N__46040\
        );

    \I__9444\ : InMux
    port map (
            O => \N__46048\,
            I => \N__46036\
        );

    \I__9443\ : Span4Mux_h
    port map (
            O => \N__46045\,
            I => \N__46031\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__46040\,
            I => \N__46031\
        );

    \I__9441\ : InMux
    port map (
            O => \N__46039\,
            I => \N__46027\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__46036\,
            I => \N__46024\
        );

    \I__9439\ : Span4Mux_v
    port map (
            O => \N__46031\,
            I => \N__46021\
        );

    \I__9438\ : InMux
    port map (
            O => \N__46030\,
            I => \N__46018\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__46027\,
            I => \N__46015\
        );

    \I__9436\ : Span4Mux_v
    port map (
            O => \N__46024\,
            I => \N__46011\
        );

    \I__9435\ : Span4Mux_v
    port map (
            O => \N__46021\,
            I => \N__46006\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__46018\,
            I => \N__46006\
        );

    \I__9433\ : Span4Mux_h
    port map (
            O => \N__46015\,
            I => \N__46003\
        );

    \I__9432\ : CascadeMux
    port map (
            O => \N__46014\,
            I => \N__46000\
        );

    \I__9431\ : Span4Mux_v
    port map (
            O => \N__46011\,
            I => \N__45996\
        );

    \I__9430\ : Span4Mux_h
    port map (
            O => \N__46006\,
            I => \N__45993\
        );

    \I__9429\ : Sp12to4
    port map (
            O => \N__46003\,
            I => \N__45990\
        );

    \I__9428\ : InMux
    port map (
            O => \N__46000\,
            I => \N__45987\
        );

    \I__9427\ : InMux
    port map (
            O => \N__45999\,
            I => \N__45984\
        );

    \I__9426\ : Span4Mux_v
    port map (
            O => \N__45996\,
            I => \N__45981\
        );

    \I__9425\ : Span4Mux_v
    port map (
            O => \N__45993\,
            I => \N__45978\
        );

    \I__9424\ : Span12Mux_v
    port map (
            O => \N__45990\,
            I => \N__45975\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__45987\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__45984\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__9421\ : Odrv4
    port map (
            O => \N__45981\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__9420\ : Odrv4
    port map (
            O => \N__45978\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__9419\ : Odrv12
    port map (
            O => \N__45975\,
            I => \c0.FRAME_MATCHER_i_3\
        );

    \I__9418\ : SRMux
    port map (
            O => \N__45964\,
            I => \N__45961\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__45961\,
            I => \N__45958\
        );

    \I__9416\ : Odrv4
    port map (
            O => \N__45958\,
            I => \c0.n3_adj_4472\
        );

    \I__9415\ : SRMux
    port map (
            O => \N__45955\,
            I => \N__45952\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__45952\,
            I => \N__45949\
        );

    \I__9413\ : Span4Mux_s3_v
    port map (
            O => \N__45949\,
            I => \N__45946\
        );

    \I__9412\ : Odrv4
    port map (
            O => \N__45946\,
            I => \c0.n3_adj_4428\
        );

    \I__9411\ : InMux
    port map (
            O => \N__45943\,
            I => \N__45937\
        );

    \I__9410\ : InMux
    port map (
            O => \N__45942\,
            I => \N__45937\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__45937\,
            I => \N__45933\
        );

    \I__9408\ : InMux
    port map (
            O => \N__45936\,
            I => \N__45930\
        );

    \I__9407\ : Span4Mux_v
    port map (
            O => \N__45933\,
            I => \N__45927\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__45930\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__9405\ : Odrv4
    port map (
            O => \N__45927\,
            I => \c0.FRAME_MATCHER_i_30\
        );

    \I__9404\ : InMux
    port map (
            O => \N__45922\,
            I => \bfn_19_31_0_\
        );

    \I__9403\ : SRMux
    port map (
            O => \N__45919\,
            I => \N__45916\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__45916\,
            I => \N__45913\
        );

    \I__9401\ : Span4Mux_v
    port map (
            O => \N__45913\,
            I => \N__45910\
        );

    \I__9400\ : Odrv4
    port map (
            O => \N__45910\,
            I => \c0.n3_adj_4426\
        );

    \I__9399\ : InMux
    port map (
            O => \N__45907\,
            I => \bfn_19_29_0_\
        );

    \I__9398\ : InMux
    port map (
            O => \N__45904\,
            I => \N__45900\
        );

    \I__9397\ : InMux
    port map (
            O => \N__45903\,
            I => \N__45897\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__45900\,
            I => \N__45891\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__45897\,
            I => \N__45891\
        );

    \I__9394\ : InMux
    port map (
            O => \N__45896\,
            I => \N__45888\
        );

    \I__9393\ : Span4Mux_v
    port map (
            O => \N__45891\,
            I => \N__45885\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__45888\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__45885\,
            I => \c0.FRAME_MATCHER_i_29\
        );

    \I__9390\ : InMux
    port map (
            O => \N__45880\,
            I => \bfn_19_30_0_\
        );

    \I__9389\ : InMux
    port map (
            O => \N__45877\,
            I => \N__45873\
        );

    \I__9388\ : CascadeMux
    port map (
            O => \N__45876\,
            I => \N__45870\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__45873\,
            I => \N__45866\
        );

    \I__9386\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45863\
        );

    \I__9385\ : InMux
    port map (
            O => \N__45869\,
            I => \N__45860\
        );

    \I__9384\ : Sp12to4
    port map (
            O => \N__45866\,
            I => \N__45857\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__45863\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__45860\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__9381\ : Odrv12
    port map (
            O => \N__45857\,
            I => \c0.FRAME_MATCHER_i_27\
        );

    \I__9380\ : InMux
    port map (
            O => \N__45850\,
            I => \bfn_19_28_0_\
        );

    \I__9379\ : SRMux
    port map (
            O => \N__45847\,
            I => \N__45844\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__45844\,
            I => \N__45841\
        );

    \I__9377\ : Odrv4
    port map (
            O => \N__45841\,
            I => \c0.n3_adj_4432\
        );

    \I__9376\ : InMux
    port map (
            O => \N__45838\,
            I => \N__45834\
        );

    \I__9375\ : CascadeMux
    port map (
            O => \N__45837\,
            I => \N__45831\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__45834\,
            I => \N__45827\
        );

    \I__9373\ : InMux
    port map (
            O => \N__45831\,
            I => \N__45824\
        );

    \I__9372\ : InMux
    port map (
            O => \N__45830\,
            I => \N__45821\
        );

    \I__9371\ : Span4Mux_v
    port map (
            O => \N__45827\,
            I => \N__45818\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__45824\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__45821\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__9368\ : Odrv4
    port map (
            O => \N__45818\,
            I => \c0.FRAME_MATCHER_i_26\
        );

    \I__9367\ : InMux
    port map (
            O => \N__45811\,
            I => \bfn_19_27_0_\
        );

    \I__9366\ : SRMux
    port map (
            O => \N__45808\,
            I => \N__45805\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__45805\,
            I => \c0.n3_adj_4433\
        );

    \I__9364\ : CascadeMux
    port map (
            O => \N__45802\,
            I => \N__45799\
        );

    \I__9363\ : InMux
    port map (
            O => \N__45799\,
            I => \N__45795\
        );

    \I__9362\ : CascadeMux
    port map (
            O => \N__45798\,
            I => \N__45792\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__45795\,
            I => \N__45788\
        );

    \I__9360\ : InMux
    port map (
            O => \N__45792\,
            I => \N__45785\
        );

    \I__9359\ : InMux
    port map (
            O => \N__45791\,
            I => \N__45782\
        );

    \I__9358\ : Span4Mux_v
    port map (
            O => \N__45788\,
            I => \N__45779\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__45785\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__45782\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__9355\ : Odrv4
    port map (
            O => \N__45779\,
            I => \c0.FRAME_MATCHER_i_25\
        );

    \I__9354\ : InMux
    port map (
            O => \N__45772\,
            I => \bfn_19_26_0_\
        );

    \I__9353\ : SRMux
    port map (
            O => \N__45769\,
            I => \N__45766\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__45766\,
            I => \N__45763\
        );

    \I__9351\ : Odrv4
    port map (
            O => \N__45763\,
            I => \c0.n3_adj_4434\
        );

    \I__9350\ : CascadeMux
    port map (
            O => \N__45760\,
            I => \N__45756\
        );

    \I__9349\ : CascadeMux
    port map (
            O => \N__45759\,
            I => \N__45753\
        );

    \I__9348\ : InMux
    port map (
            O => \N__45756\,
            I => \N__45750\
        );

    \I__9347\ : InMux
    port map (
            O => \N__45753\,
            I => \N__45746\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__45750\,
            I => \N__45743\
        );

    \I__9345\ : InMux
    port map (
            O => \N__45749\,
            I => \N__45740\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__45746\,
            I => \N__45737\
        );

    \I__9343\ : Odrv4
    port map (
            O => \N__45743\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__45740\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__9341\ : Odrv4
    port map (
            O => \N__45737\,
            I => \c0.FRAME_MATCHER_i_24\
        );

    \I__9340\ : InMux
    port map (
            O => \N__45730\,
            I => \bfn_19_25_0_\
        );

    \I__9339\ : SRMux
    port map (
            O => \N__45727\,
            I => \N__45724\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__45724\,
            I => \N__45721\
        );

    \I__9337\ : Span4Mux_h
    port map (
            O => \N__45721\,
            I => \N__45718\
        );

    \I__9336\ : Odrv4
    port map (
            O => \N__45718\,
            I => \c0.n3_adj_4435\
        );

    \I__9335\ : InMux
    port map (
            O => \N__45715\,
            I => \N__45711\
        );

    \I__9334\ : CascadeMux
    port map (
            O => \N__45714\,
            I => \N__45708\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__45711\,
            I => \N__45704\
        );

    \I__9332\ : InMux
    port map (
            O => \N__45708\,
            I => \N__45701\
        );

    \I__9331\ : InMux
    port map (
            O => \N__45707\,
            I => \N__45698\
        );

    \I__9330\ : Span4Mux_h
    port map (
            O => \N__45704\,
            I => \N__45695\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__45701\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__9328\ : LocalMux
    port map (
            O => \N__45698\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__45695\,
            I => \c0.FRAME_MATCHER_i_23\
        );

    \I__9326\ : InMux
    port map (
            O => \N__45688\,
            I => \bfn_19_24_0_\
        );

    \I__9325\ : SRMux
    port map (
            O => \N__45685\,
            I => \N__45682\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__45682\,
            I => \N__45679\
        );

    \I__9323\ : Odrv12
    port map (
            O => \N__45679\,
            I => \c0.n3_adj_4436\
        );

    \I__9322\ : InMux
    port map (
            O => \N__45676\,
            I => \N__45671\
        );

    \I__9321\ : InMux
    port map (
            O => \N__45675\,
            I => \N__45668\
        );

    \I__9320\ : InMux
    port map (
            O => \N__45674\,
            I => \N__45665\
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__45671\,
            I => \N__45662\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__45668\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__45665\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__9316\ : Odrv4
    port map (
            O => \N__45662\,
            I => \c0.FRAME_MATCHER_i_22\
        );

    \I__9315\ : InMux
    port map (
            O => \N__45655\,
            I => \bfn_19_23_0_\
        );

    \I__9314\ : SRMux
    port map (
            O => \N__45652\,
            I => \N__45649\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__45649\,
            I => \N__45646\
        );

    \I__9312\ : Span4Mux_h
    port map (
            O => \N__45646\,
            I => \N__45643\
        );

    \I__9311\ : Odrv4
    port map (
            O => \N__45643\,
            I => \c0.n3_adj_4438\
        );

    \I__9310\ : CascadeMux
    port map (
            O => \N__45640\,
            I => \N__45637\
        );

    \I__9309\ : InMux
    port map (
            O => \N__45637\,
            I => \N__45634\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__45634\,
            I => \N__45631\
        );

    \I__9307\ : Span4Mux_h
    port map (
            O => \N__45631\,
            I => \N__45626\
        );

    \I__9306\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45623\
        );

    \I__9305\ : InMux
    port map (
            O => \N__45629\,
            I => \N__45620\
        );

    \I__9304\ : Odrv4
    port map (
            O => \N__45626\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__45623\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__45620\,
            I => \c0.FRAME_MATCHER_i_21\
        );

    \I__9301\ : InMux
    port map (
            O => \N__45613\,
            I => \bfn_19_22_0_\
        );

    \I__9300\ : SRMux
    port map (
            O => \N__45610\,
            I => \N__45607\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__45607\,
            I => \N__45604\
        );

    \I__9298\ : Odrv4
    port map (
            O => \N__45604\,
            I => \c0.n3_adj_4440\
        );

    \I__9297\ : SRMux
    port map (
            O => \N__45601\,
            I => \N__45598\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__45598\,
            I => \N__45595\
        );

    \I__9295\ : Span4Mux_h
    port map (
            O => \N__45595\,
            I => \N__45592\
        );

    \I__9294\ : Span4Mux_h
    port map (
            O => \N__45592\,
            I => \N__45589\
        );

    \I__9293\ : Odrv4
    port map (
            O => \N__45589\,
            I => \c0.n3_adj_4444\
        );

    \I__9292\ : InMux
    port map (
            O => \N__45586\,
            I => \bfn_19_21_0_\
        );

    \I__9291\ : CascadeMux
    port map (
            O => \N__45583\,
            I => \N__45580\
        );

    \I__9290\ : InMux
    port map (
            O => \N__45580\,
            I => \N__45576\
        );

    \I__9289\ : InMux
    port map (
            O => \N__45579\,
            I => \N__45573\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__45576\,
            I => \N__45570\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__45573\,
            I => \N__45566\
        );

    \I__9286\ : Span4Mux_h
    port map (
            O => \N__45570\,
            I => \N__45563\
        );

    \I__9285\ : InMux
    port map (
            O => \N__45569\,
            I => \N__45560\
        );

    \I__9284\ : Span4Mux_h
    port map (
            O => \N__45566\,
            I => \N__45557\
        );

    \I__9283\ : Odrv4
    port map (
            O => \N__45563\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__45560\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__9281\ : Odrv4
    port map (
            O => \N__45557\,
            I => \c0.FRAME_MATCHER_i_18\
        );

    \I__9280\ : InMux
    port map (
            O => \N__45550\,
            I => \bfn_19_19_0_\
        );

    \I__9279\ : SRMux
    port map (
            O => \N__45547\,
            I => \N__45544\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__45544\,
            I => \N__45541\
        );

    \I__9277\ : Span4Mux_v
    port map (
            O => \N__45541\,
            I => \N__45538\
        );

    \I__9276\ : Odrv4
    port map (
            O => \N__45538\,
            I => \c0.n3_adj_4446\
        );

    \I__9275\ : CascadeMux
    port map (
            O => \N__45535\,
            I => \N__45531\
        );

    \I__9274\ : InMux
    port map (
            O => \N__45534\,
            I => \N__45528\
        );

    \I__9273\ : InMux
    port map (
            O => \N__45531\,
            I => \N__45525\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__45528\,
            I => \N__45521\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__45525\,
            I => \N__45518\
        );

    \I__9270\ : InMux
    port map (
            O => \N__45524\,
            I => \N__45515\
        );

    \I__9269\ : Span4Mux_v
    port map (
            O => \N__45521\,
            I => \N__45512\
        );

    \I__9268\ : Odrv4
    port map (
            O => \N__45518\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__45515\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__9266\ : Odrv4
    port map (
            O => \N__45512\,
            I => \c0.FRAME_MATCHER_i_19\
        );

    \I__9265\ : InMux
    port map (
            O => \N__45505\,
            I => \bfn_19_20_0_\
        );

    \I__9264\ : CascadeMux
    port map (
            O => \N__45502\,
            I => \N__45499\
        );

    \I__9263\ : InMux
    port map (
            O => \N__45499\,
            I => \N__45495\
        );

    \I__9262\ : InMux
    port map (
            O => \N__45498\,
            I => \N__45492\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__45495\,
            I => \N__45488\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__45492\,
            I => \N__45485\
        );

    \I__9259\ : InMux
    port map (
            O => \N__45491\,
            I => \N__45482\
        );

    \I__9258\ : Span4Mux_v
    port map (
            O => \N__45488\,
            I => \N__45477\
        );

    \I__9257\ : Span4Mux_v
    port map (
            O => \N__45485\,
            I => \N__45477\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__45482\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__9255\ : Odrv4
    port map (
            O => \N__45477\,
            I => \c0.FRAME_MATCHER_i_17\
        );

    \I__9254\ : InMux
    port map (
            O => \N__45472\,
            I => \bfn_19_18_0_\
        );

    \I__9253\ : SRMux
    port map (
            O => \N__45469\,
            I => \N__45466\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__45466\,
            I => \N__45463\
        );

    \I__9251\ : Span4Mux_h
    port map (
            O => \N__45463\,
            I => \N__45460\
        );

    \I__9250\ : Span4Mux_v
    port map (
            O => \N__45460\,
            I => \N__45457\
        );

    \I__9249\ : Odrv4
    port map (
            O => \N__45457\,
            I => \c0.n3_adj_4448\
        );

    \I__9248\ : InMux
    port map (
            O => \N__45454\,
            I => \bfn_19_17_0_\
        );

    \I__9247\ : SRMux
    port map (
            O => \N__45451\,
            I => \N__45448\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__45448\,
            I => \N__45445\
        );

    \I__9245\ : Odrv12
    port map (
            O => \N__45445\,
            I => \c0.n3_adj_4450\
        );

    \I__9244\ : InMux
    port map (
            O => \N__45442\,
            I => \bfn_19_16_0_\
        );

    \I__9243\ : CascadeMux
    port map (
            O => \N__45439\,
            I => \N__45436\
        );

    \I__9242\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45432\
        );

    \I__9241\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45429\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__45432\,
            I => \N__45426\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__45429\,
            I => \N__45422\
        );

    \I__9238\ : Span4Mux_h
    port map (
            O => \N__45426\,
            I => \N__45419\
        );

    \I__9237\ : InMux
    port map (
            O => \N__45425\,
            I => \N__45416\
        );

    \I__9236\ : Span4Mux_v
    port map (
            O => \N__45422\,
            I => \N__45413\
        );

    \I__9235\ : Odrv4
    port map (
            O => \N__45419\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__45416\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__9233\ : Odrv4
    port map (
            O => \N__45413\,
            I => \c0.FRAME_MATCHER_i_14\
        );

    \I__9232\ : InMux
    port map (
            O => \N__45406\,
            I => \bfn_19_15_0_\
        );

    \I__9231\ : SRMux
    port map (
            O => \N__45403\,
            I => \N__45400\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__45400\,
            I => \N__45397\
        );

    \I__9229\ : Span4Mux_v
    port map (
            O => \N__45397\,
            I => \N__45394\
        );

    \I__9228\ : Sp12to4
    port map (
            O => \N__45394\,
            I => \N__45391\
        );

    \I__9227\ : Odrv12
    port map (
            O => \N__45391\,
            I => \c0.n3_adj_4453\
        );

    \I__9226\ : InMux
    port map (
            O => \N__45388\,
            I => \bfn_19_14_0_\
        );

    \I__9225\ : CascadeMux
    port map (
            O => \N__45385\,
            I => \N__45381\
        );

    \I__9224\ : CascadeMux
    port map (
            O => \N__45384\,
            I => \N__45378\
        );

    \I__9223\ : InMux
    port map (
            O => \N__45381\,
            I => \N__45375\
        );

    \I__9222\ : InMux
    port map (
            O => \N__45378\,
            I => \N__45372\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__45375\,
            I => \N__45369\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__45372\,
            I => \N__45366\
        );

    \I__9219\ : Span4Mux_h
    port map (
            O => \N__45369\,
            I => \N__45363\
        );

    \I__9218\ : Span4Mux_h
    port map (
            O => \N__45366\,
            I => \N__45359\
        );

    \I__9217\ : Span4Mux_v
    port map (
            O => \N__45363\,
            I => \N__45356\
        );

    \I__9216\ : InMux
    port map (
            O => \N__45362\,
            I => \N__45353\
        );

    \I__9215\ : Odrv4
    port map (
            O => \N__45359\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__9214\ : Odrv4
    port map (
            O => \N__45356\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__45353\,
            I => \c0.FRAME_MATCHER_i_12\
        );

    \I__9212\ : InMux
    port map (
            O => \N__45346\,
            I => \bfn_19_13_0_\
        );

    \I__9211\ : SRMux
    port map (
            O => \N__45343\,
            I => \N__45340\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__45340\,
            I => \N__45337\
        );

    \I__9209\ : Span4Mux_v
    port map (
            O => \N__45337\,
            I => \N__45334\
        );

    \I__9208\ : Odrv4
    port map (
            O => \N__45334\,
            I => \c0.n3_adj_4456\
        );

    \I__9207\ : InMux
    port map (
            O => \N__45331\,
            I => \N__45328\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__45328\,
            I => \N__45324\
        );

    \I__9205\ : InMux
    port map (
            O => \N__45327\,
            I => \N__45321\
        );

    \I__9204\ : Sp12to4
    port map (
            O => \N__45324\,
            I => \N__45318\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__45321\,
            I => \N__45315\
        );

    \I__9202\ : Span12Mux_h
    port map (
            O => \N__45318\,
            I => \N__45309\
        );

    \I__9201\ : Sp12to4
    port map (
            O => \N__45315\,
            I => \N__45309\
        );

    \I__9200\ : InMux
    port map (
            O => \N__45314\,
            I => \N__45306\
        );

    \I__9199\ : Odrv12
    port map (
            O => \N__45309\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__45306\,
            I => \c0.FRAME_MATCHER_i_11\
        );

    \I__9197\ : InMux
    port map (
            O => \N__45301\,
            I => \bfn_19_12_0_\
        );

    \I__9196\ : SRMux
    port map (
            O => \N__45298\,
            I => \N__45295\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__45295\,
            I => \N__45292\
        );

    \I__9194\ : Span4Mux_h
    port map (
            O => \N__45292\,
            I => \N__45289\
        );

    \I__9193\ : Span4Mux_v
    port map (
            O => \N__45289\,
            I => \N__45286\
        );

    \I__9192\ : Span4Mux_v
    port map (
            O => \N__45286\,
            I => \N__45283\
        );

    \I__9191\ : Odrv4
    port map (
            O => \N__45283\,
            I => \c0.n3_adj_4458\
        );

    \I__9190\ : CascadeMux
    port map (
            O => \N__45280\,
            I => \N__45276\
        );

    \I__9189\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45273\
        );

    \I__9188\ : InMux
    port map (
            O => \N__45276\,
            I => \N__45270\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__45273\,
            I => \N__45267\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__45270\,
            I => \N__45261\
        );

    \I__9185\ : Span4Mux_v
    port map (
            O => \N__45267\,
            I => \N__45261\
        );

    \I__9184\ : InMux
    port map (
            O => \N__45266\,
            I => \N__45258\
        );

    \I__9183\ : Sp12to4
    port map (
            O => \N__45261\,
            I => \N__45255\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__45258\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__9181\ : Odrv12
    port map (
            O => \N__45255\,
            I => \c0.FRAME_MATCHER_i_9\
        );

    \I__9180\ : InMux
    port map (
            O => \N__45250\,
            I => \bfn_19_10_0_\
        );

    \I__9179\ : SRMux
    port map (
            O => \N__45247\,
            I => \N__45244\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__45244\,
            I => \N__45241\
        );

    \I__9177\ : Span4Mux_v
    port map (
            O => \N__45241\,
            I => \N__45238\
        );

    \I__9176\ : Span4Mux_h
    port map (
            O => \N__45238\,
            I => \N__45235\
        );

    \I__9175\ : Odrv4
    port map (
            O => \N__45235\,
            I => \c0.n3_adj_4462\
        );

    \I__9174\ : InMux
    port map (
            O => \N__45232\,
            I => \bfn_19_11_0_\
        );

    \I__9173\ : InMux
    port map (
            O => \N__45229\,
            I => \N__45226\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__45226\,
            I => \N__45222\
        );

    \I__9171\ : InMux
    port map (
            O => \N__45225\,
            I => \N__45219\
        );

    \I__9170\ : Span4Mux_v
    port map (
            O => \N__45222\,
            I => \N__45216\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__45219\,
            I => \N__45212\
        );

    \I__9168\ : Span4Mux_v
    port map (
            O => \N__45216\,
            I => \N__45209\
        );

    \I__9167\ : InMux
    port map (
            O => \N__45215\,
            I => \N__45206\
        );

    \I__9166\ : Sp12to4
    port map (
            O => \N__45212\,
            I => \N__45203\
        );

    \I__9165\ : Odrv4
    port map (
            O => \N__45209\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__45206\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__9163\ : Odrv12
    port map (
            O => \N__45203\,
            I => \c0.FRAME_MATCHER_i_8\
        );

    \I__9162\ : InMux
    port map (
            O => \N__45196\,
            I => \bfn_19_9_0_\
        );

    \I__9161\ : SRMux
    port map (
            O => \N__45193\,
            I => \N__45190\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__45190\,
            I => \N__45187\
        );

    \I__9159\ : Span4Mux_h
    port map (
            O => \N__45187\,
            I => \N__45184\
        );

    \I__9158\ : Span4Mux_v
    port map (
            O => \N__45184\,
            I => \N__45181\
        );

    \I__9157\ : Odrv4
    port map (
            O => \N__45181\,
            I => \c0.n3_adj_4463\
        );

    \I__9156\ : InMux
    port map (
            O => \N__45178\,
            I => \N__45175\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__45175\,
            I => \N__45171\
        );

    \I__9154\ : InMux
    port map (
            O => \N__45174\,
            I => \N__45168\
        );

    \I__9153\ : Sp12to4
    port map (
            O => \N__45171\,
            I => \N__45165\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__45168\,
            I => \N__45162\
        );

    \I__9151\ : Span12Mux_h
    port map (
            O => \N__45165\,
            I => \N__45159\
        );

    \I__9150\ : Span4Mux_v
    port map (
            O => \N__45162\,
            I => \N__45156\
        );

    \I__9149\ : Span12Mux_v
    port map (
            O => \N__45159\,
            I => \N__45152\
        );

    \I__9148\ : Span4Mux_v
    port map (
            O => \N__45156\,
            I => \N__45149\
        );

    \I__9147\ : InMux
    port map (
            O => \N__45155\,
            I => \N__45146\
        );

    \I__9146\ : Odrv12
    port map (
            O => \N__45152\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__9145\ : Odrv4
    port map (
            O => \N__45149\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__45146\,
            I => \c0.FRAME_MATCHER_i_7\
        );

    \I__9143\ : InMux
    port map (
            O => \N__45139\,
            I => \bfn_19_8_0_\
        );

    \I__9142\ : SRMux
    port map (
            O => \N__45136\,
            I => \N__45133\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__45133\,
            I => \N__45130\
        );

    \I__9140\ : Sp12to4
    port map (
            O => \N__45130\,
            I => \N__45127\
        );

    \I__9139\ : Span12Mux_h
    port map (
            O => \N__45127\,
            I => \N__45124\
        );

    \I__9138\ : Span12Mux_v
    port map (
            O => \N__45124\,
            I => \N__45121\
        );

    \I__9137\ : Odrv12
    port map (
            O => \N__45121\,
            I => \c0.n3_adj_4465\
        );

    \I__9136\ : InMux
    port map (
            O => \N__45118\,
            I => \bfn_19_7_0_\
        );

    \I__9135\ : SRMux
    port map (
            O => \N__45115\,
            I => \N__45112\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__45112\,
            I => \N__45109\
        );

    \I__9133\ : Span4Mux_v
    port map (
            O => \N__45109\,
            I => \N__45106\
        );

    \I__9132\ : Span4Mux_v
    port map (
            O => \N__45106\,
            I => \N__45103\
        );

    \I__9131\ : Odrv4
    port map (
            O => \N__45103\,
            I => \c0.n3_adj_4467\
        );

    \I__9130\ : InMux
    port map (
            O => \N__45100\,
            I => \bfn_19_6_0_\
        );

    \I__9129\ : SRMux
    port map (
            O => \N__45097\,
            I => \N__45094\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__45094\,
            I => \N__45091\
        );

    \I__9127\ : Span4Mux_v
    port map (
            O => \N__45091\,
            I => \N__45088\
        );

    \I__9126\ : Odrv4
    port map (
            O => \N__45088\,
            I => \c0.n3_adj_4468\
        );

    \I__9125\ : CascadeMux
    port map (
            O => \N__45085\,
            I => \N__45082\
        );

    \I__9124\ : InMux
    port map (
            O => \N__45082\,
            I => \N__45078\
        );

    \I__9123\ : InMux
    port map (
            O => \N__45081\,
            I => \N__45074\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__45078\,
            I => \N__45070\
        );

    \I__9121\ : CascadeMux
    port map (
            O => \N__45077\,
            I => \N__45066\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__45074\,
            I => \N__45061\
        );

    \I__9119\ : InMux
    port map (
            O => \N__45073\,
            I => \N__45058\
        );

    \I__9118\ : Span4Mux_v
    port map (
            O => \N__45070\,
            I => \N__45055\
        );

    \I__9117\ : InMux
    port map (
            O => \N__45069\,
            I => \N__45052\
        );

    \I__9116\ : InMux
    port map (
            O => \N__45066\,
            I => \N__45049\
        );

    \I__9115\ : InMux
    port map (
            O => \N__45065\,
            I => \N__45044\
        );

    \I__9114\ : InMux
    port map (
            O => \N__45064\,
            I => \N__45044\
        );

    \I__9113\ : Span4Mux_h
    port map (
            O => \N__45061\,
            I => \N__45039\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__45058\,
            I => \N__45039\
        );

    \I__9111\ : Span4Mux_h
    port map (
            O => \N__45055\,
            I => \N__45034\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__45052\,
            I => \N__45034\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__45049\,
            I => \N__45027\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__45044\,
            I => \N__45027\
        );

    \I__9107\ : Span4Mux_v
    port map (
            O => \N__45039\,
            I => \N__45027\
        );

    \I__9106\ : Span4Mux_v
    port map (
            O => \N__45034\,
            I => \N__45022\
        );

    \I__9105\ : Span4Mux_v
    port map (
            O => \N__45027\,
            I => \N__45022\
        );

    \I__9104\ : Span4Mux_v
    port map (
            O => \N__45022\,
            I => \N__45019\
        );

    \I__9103\ : Span4Mux_v
    port map (
            O => \N__45019\,
            I => \N__45015\
        );

    \I__9102\ : InMux
    port map (
            O => \N__45018\,
            I => \N__45012\
        );

    \I__9101\ : Odrv4
    port map (
            O => \N__45015\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__45012\,
            I => \c0.FRAME_MATCHER_i_4\
        );

    \I__9099\ : InMux
    port map (
            O => \N__45007\,
            I => \bfn_19_5_0_\
        );

    \I__9098\ : SRMux
    port map (
            O => \N__45004\,
            I => \N__45001\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__45001\,
            I => \N__44998\
        );

    \I__9096\ : Span4Mux_v
    port map (
            O => \N__44998\,
            I => \N__44995\
        );

    \I__9095\ : Span4Mux_v
    port map (
            O => \N__44995\,
            I => \N__44992\
        );

    \I__9094\ : Span4Mux_v
    port map (
            O => \N__44992\,
            I => \N__44989\
        );

    \I__9093\ : Odrv4
    port map (
            O => \N__44989\,
            I => \c0.n3_adj_4470\
        );

    \I__9092\ : InMux
    port map (
            O => \N__44986\,
            I => \bfn_19_4_0_\
        );

    \I__9091\ : InMux
    port map (
            O => \N__44983\,
            I => \bfn_19_3_0_\
        );

    \I__9090\ : SRMux
    port map (
            O => \N__44980\,
            I => \N__44977\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__44977\,
            I => \N__44974\
        );

    \I__9088\ : Span4Mux_s2_v
    port map (
            O => \N__44974\,
            I => \N__44971\
        );

    \I__9087\ : Odrv4
    port map (
            O => \N__44971\,
            I => \c0.n3\
        );

    \I__9086\ : InMux
    port map (
            O => \N__44968\,
            I => \bfn_19_2_0_\
        );

    \I__9085\ : InMux
    port map (
            O => \N__44965\,
            I => \N__44962\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__44962\,
            I => \N__44959\
        );

    \I__9083\ : Span4Mux_h
    port map (
            O => \N__44959\,
            I => \N__44956\
        );

    \I__9082\ : Odrv4
    port map (
            O => \N__44956\,
            I => \c0.n29_adj_4382\
        );

    \I__9081\ : CascadeMux
    port map (
            O => \N__44953\,
            I => \N__44950\
        );

    \I__9080\ : InMux
    port map (
            O => \N__44950\,
            I => \N__44947\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__44947\,
            I => \N__44944\
        );

    \I__9078\ : Span4Mux_s1_v
    port map (
            O => \N__44944\,
            I => \N__44941\
        );

    \I__9077\ : Span4Mux_v
    port map (
            O => \N__44941\,
            I => \N__44938\
        );

    \I__9076\ : Span4Mux_h
    port map (
            O => \N__44938\,
            I => \N__44935\
        );

    \I__9075\ : Span4Mux_h
    port map (
            O => \N__44935\,
            I => \N__44932\
        );

    \I__9074\ : Odrv4
    port map (
            O => \N__44932\,
            I => \c0.n161\
        );

    \I__9073\ : InMux
    port map (
            O => \N__44929\,
            I => \N__44926\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__44926\,
            I => \N__44922\
        );

    \I__9071\ : InMux
    port map (
            O => \N__44925\,
            I => \N__44918\
        );

    \I__9070\ : Span4Mux_h
    port map (
            O => \N__44922\,
            I => \N__44915\
        );

    \I__9069\ : InMux
    port map (
            O => \N__44921\,
            I => \N__44912\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__44918\,
            I => data_in_frame_22_1
        );

    \I__9067\ : Odrv4
    port map (
            O => \N__44915\,
            I => data_in_frame_22_1
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__44912\,
            I => data_in_frame_22_1
        );

    \I__9065\ : CascadeMux
    port map (
            O => \N__44905\,
            I => \c0.rx.n22611_cascade_\
        );

    \I__9064\ : CascadeMux
    port map (
            O => \N__44902\,
            I => \c0.rx.n8_cascade_\
        );

    \I__9063\ : CascadeMux
    port map (
            O => \N__44899\,
            I => \N__44895\
        );

    \I__9062\ : CascadeMux
    port map (
            O => \N__44898\,
            I => \N__44892\
        );

    \I__9061\ : InMux
    port map (
            O => \N__44895\,
            I => \N__44889\
        );

    \I__9060\ : InMux
    port map (
            O => \N__44892\,
            I => \N__44886\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__44889\,
            I => \c0.data_in_frame_29_2\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__44886\,
            I => \c0.data_in_frame_29_2\
        );

    \I__9057\ : InMux
    port map (
            O => \N__44881\,
            I => \N__44877\
        );

    \I__9056\ : InMux
    port map (
            O => \N__44880\,
            I => \N__44874\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__44877\,
            I => \N__44871\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__44874\,
            I => \c0.data_in_frame_29_1\
        );

    \I__9053\ : Odrv12
    port map (
            O => \N__44871\,
            I => \c0.data_in_frame_29_1\
        );

    \I__9052\ : CascadeMux
    port map (
            O => \N__44866\,
            I => \c0.n23388_cascade_\
        );

    \I__9051\ : InMux
    port map (
            O => \N__44863\,
            I => \N__44860\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__44860\,
            I => \c0.n30_adj_4299\
        );

    \I__9049\ : CascadeMux
    port map (
            O => \N__44857\,
            I => \c0.n15_adj_4376_cascade_\
        );

    \I__9048\ : InMux
    port map (
            O => \N__44854\,
            I => \N__44851\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__44851\,
            I => \N__44848\
        );

    \I__9046\ : Odrv12
    port map (
            O => \N__44848\,
            I => \c0.n17_adj_4378\
        );

    \I__9045\ : CascadeMux
    port map (
            O => \N__44845\,
            I => \c0.n18_adj_4379_cascade_\
        );

    \I__9044\ : InMux
    port map (
            O => \N__44842\,
            I => \N__44839\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__44839\,
            I => \c0.n27_adj_4383\
        );

    \I__9042\ : CascadeMux
    port map (
            O => \N__44836\,
            I => \c0.n30_adj_4380_cascade_\
        );

    \I__9041\ : InMux
    port map (
            O => \N__44833\,
            I => \N__44830\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__44830\,
            I => \N__44827\
        );

    \I__9039\ : Span4Mux_v
    port map (
            O => \N__44827\,
            I => \N__44824\
        );

    \I__9038\ : Odrv4
    port map (
            O => \N__44824\,
            I => \c0.n28_adj_4381\
        );

    \I__9037\ : InMux
    port map (
            O => \N__44821\,
            I => \N__44818\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__44818\,
            I => \N__44814\
        );

    \I__9035\ : InMux
    port map (
            O => \N__44817\,
            I => \N__44811\
        );

    \I__9034\ : Odrv4
    port map (
            O => \N__44814\,
            I => \c0.n13000\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__44811\,
            I => \c0.n13000\
        );

    \I__9032\ : CascadeMux
    port map (
            O => \N__44806\,
            I => \c0.n10_adj_4286_cascade_\
        );

    \I__9031\ : CascadeMux
    port map (
            O => \N__44803\,
            I => \N__44799\
        );

    \I__9030\ : InMux
    port map (
            O => \N__44802\,
            I => \N__44794\
        );

    \I__9029\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44794\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__44794\,
            I => \c0.data_in_frame_28_2\
        );

    \I__9027\ : CascadeMux
    port map (
            O => \N__44791\,
            I => \N__44787\
        );

    \I__9026\ : InMux
    port map (
            O => \N__44790\,
            I => \N__44784\
        );

    \I__9025\ : InMux
    port map (
            O => \N__44787\,
            I => \N__44781\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__44784\,
            I => \N__44778\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__44781\,
            I => \c0.data_in_frame_29_0\
        );

    \I__9022\ : Odrv4
    port map (
            O => \N__44778\,
            I => \c0.data_in_frame_29_0\
        );

    \I__9021\ : InMux
    port map (
            O => \N__44773\,
            I => \N__44770\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__44770\,
            I => \N__44767\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__44767\,
            I => \N__44764\
        );

    \I__9018\ : Span4Mux_v
    port map (
            O => \N__44764\,
            I => \N__44761\
        );

    \I__9017\ : Span4Mux_v
    port map (
            O => \N__44761\,
            I => \N__44758\
        );

    \I__9016\ : Odrv4
    port map (
            O => \N__44758\,
            I => \c0.n17600\
        );

    \I__9015\ : CascadeMux
    port map (
            O => \N__44755\,
            I => \c0.n19_cascade_\
        );

    \I__9014\ : InMux
    port map (
            O => \N__44752\,
            I => \N__44749\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__44749\,
            I => \c0.n23389\
        );

    \I__9012\ : CascadeMux
    port map (
            O => \N__44746\,
            I => \c0.n32_adj_4295_cascade_\
        );

    \I__9011\ : InMux
    port map (
            O => \N__44743\,
            I => \N__44740\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__44740\,
            I => \N__44737\
        );

    \I__9009\ : Odrv4
    port map (
            O => \N__44737\,
            I => \c0.n23523\
        );

    \I__9008\ : InMux
    port map (
            O => \N__44734\,
            I => \N__44731\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__44731\,
            I => \c0.n34\
        );

    \I__9006\ : InMux
    port map (
            O => \N__44728\,
            I => \N__44725\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__44725\,
            I => \N__44720\
        );

    \I__9004\ : InMux
    port map (
            O => \N__44724\,
            I => \N__44715\
        );

    \I__9003\ : InMux
    port map (
            O => \N__44723\,
            I => \N__44715\
        );

    \I__9002\ : Odrv4
    port map (
            O => \N__44720\,
            I => \c0.n17790\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__44715\,
            I => \c0.n17790\
        );

    \I__9000\ : InMux
    port map (
            O => \N__44710\,
            I => \N__44707\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__44707\,
            I => \N__44704\
        );

    \I__8998\ : Span4Mux_v
    port map (
            O => \N__44704\,
            I => \N__44699\
        );

    \I__8997\ : CascadeMux
    port map (
            O => \N__44703\,
            I => \N__44692\
        );

    \I__8996\ : InMux
    port map (
            O => \N__44702\,
            I => \N__44689\
        );

    \I__8995\ : Span4Mux_v
    port map (
            O => \N__44699\,
            I => \N__44686\
        );

    \I__8994\ : InMux
    port map (
            O => \N__44698\,
            I => \N__44683\
        );

    \I__8993\ : InMux
    port map (
            O => \N__44697\,
            I => \N__44678\
        );

    \I__8992\ : InMux
    port map (
            O => \N__44696\,
            I => \N__44678\
        );

    \I__8991\ : InMux
    port map (
            O => \N__44695\,
            I => \N__44673\
        );

    \I__8990\ : InMux
    port map (
            O => \N__44692\,
            I => \N__44673\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__44689\,
            I => data_in_frame_1_0
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__44686\,
            I => data_in_frame_1_0
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__44683\,
            I => data_in_frame_1_0
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__44678\,
            I => data_in_frame_1_0
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__44673\,
            I => data_in_frame_1_0
        );

    \I__8984\ : CascadeMux
    port map (
            O => \N__44662\,
            I => \N__44656\
        );

    \I__8983\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44650\
        );

    \I__8982\ : InMux
    port map (
            O => \N__44660\,
            I => \N__44647\
        );

    \I__8981\ : InMux
    port map (
            O => \N__44659\,
            I => \N__44644\
        );

    \I__8980\ : InMux
    port map (
            O => \N__44656\,
            I => \N__44637\
        );

    \I__8979\ : InMux
    port map (
            O => \N__44655\,
            I => \N__44637\
        );

    \I__8978\ : InMux
    port map (
            O => \N__44654\,
            I => \N__44637\
        );

    \I__8977\ : InMux
    port map (
            O => \N__44653\,
            I => \N__44634\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__44650\,
            I => n23726
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__44647\,
            I => n23726
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__44644\,
            I => n23726
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__44637\,
            I => n23726
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__44634\,
            I => n23726
        );

    \I__8971\ : CascadeMux
    port map (
            O => \N__44623\,
            I => \N__44620\
        );

    \I__8970\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44615\
        );

    \I__8969\ : InMux
    port map (
            O => \N__44619\,
            I => \N__44612\
        );

    \I__8968\ : CascadeMux
    port map (
            O => \N__44618\,
            I => \N__44609\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__44615\,
            I => \N__44603\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__44612\,
            I => \N__44600\
        );

    \I__8965\ : InMux
    port map (
            O => \N__44609\,
            I => \N__44597\
        );

    \I__8964\ : InMux
    port map (
            O => \N__44608\,
            I => \N__44592\
        );

    \I__8963\ : InMux
    port map (
            O => \N__44607\,
            I => \N__44592\
        );

    \I__8962\ : InMux
    port map (
            O => \N__44606\,
            I => \N__44588\
        );

    \I__8961\ : Span4Mux_v
    port map (
            O => \N__44603\,
            I => \N__44583\
        );

    \I__8960\ : Span4Mux_v
    port map (
            O => \N__44600\,
            I => \N__44583\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__44597\,
            I => \N__44578\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__44592\,
            I => \N__44578\
        );

    \I__8957\ : InMux
    port map (
            O => \N__44591\,
            I => \N__44575\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__44588\,
            I => \N__44572\
        );

    \I__8955\ : Span4Mux_h
    port map (
            O => \N__44583\,
            I => \N__44567\
        );

    \I__8954\ : Span4Mux_v
    port map (
            O => \N__44578\,
            I => \N__44567\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__44575\,
            I => control_mode_0
        );

    \I__8952\ : Odrv4
    port map (
            O => \N__44572\,
            I => control_mode_0
        );

    \I__8951\ : Odrv4
    port map (
            O => \N__44567\,
            I => control_mode_0
        );

    \I__8950\ : CascadeMux
    port map (
            O => \N__44560\,
            I => \N__44556\
        );

    \I__8949\ : InMux
    port map (
            O => \N__44559\,
            I => \N__44553\
        );

    \I__8948\ : InMux
    port map (
            O => \N__44556\,
            I => \N__44550\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__44553\,
            I => \c0.data_in_frame_29_4\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__44550\,
            I => \c0.data_in_frame_29_4\
        );

    \I__8945\ : CascadeMux
    port map (
            O => \N__44545\,
            I => \n4_cascade_\
        );

    \I__8944\ : CascadeMux
    port map (
            O => \N__44542\,
            I => \N__44538\
        );

    \I__8943\ : CascadeMux
    port map (
            O => \N__44541\,
            I => \N__44535\
        );

    \I__8942\ : InMux
    port map (
            O => \N__44538\,
            I => \N__44529\
        );

    \I__8941\ : InMux
    port map (
            O => \N__44535\,
            I => \N__44529\
        );

    \I__8940\ : InMux
    port map (
            O => \N__44534\,
            I => \N__44526\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__44529\,
            I => \N__44523\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__44526\,
            I => \c0.data_in_frame_4_6\
        );

    \I__8937\ : Odrv12
    port map (
            O => \N__44523\,
            I => \c0.data_in_frame_4_6\
        );

    \I__8936\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44515\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__44515\,
            I => \N__44512\
        );

    \I__8934\ : Odrv4
    port map (
            O => \N__44512\,
            I => n4
        );

    \I__8933\ : CascadeMux
    port map (
            O => \N__44509\,
            I => \c0.n21758_cascade_\
        );

    \I__8932\ : CascadeMux
    port map (
            O => \N__44506\,
            I => \N__44502\
        );

    \I__8931\ : CascadeMux
    port map (
            O => \N__44505\,
            I => \N__44499\
        );

    \I__8930\ : InMux
    port map (
            O => \N__44502\,
            I => \N__44496\
        );

    \I__8929\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44493\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__44496\,
            I => \N__44488\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__44493\,
            I => \N__44485\
        );

    \I__8926\ : InMux
    port map (
            O => \N__44492\,
            I => \N__44480\
        );

    \I__8925\ : InMux
    port map (
            O => \N__44491\,
            I => \N__44480\
        );

    \I__8924\ : Odrv4
    port map (
            O => \N__44488\,
            I => \c0.data_in_frame_2_4\
        );

    \I__8923\ : Odrv12
    port map (
            O => \N__44485\,
            I => \c0.data_in_frame_2_4\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__44480\,
            I => \c0.data_in_frame_2_4\
        );

    \I__8921\ : CascadeMux
    port map (
            O => \N__44473\,
            I => \N__44470\
        );

    \I__8920\ : InMux
    port map (
            O => \N__44470\,
            I => \N__44465\
        );

    \I__8919\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44462\
        );

    \I__8918\ : InMux
    port map (
            O => \N__44468\,
            I => \N__44459\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__44465\,
            I => \N__44454\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__44462\,
            I => \N__44454\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__44459\,
            I => \c0.data_in_frame_5_0\
        );

    \I__8914\ : Odrv4
    port map (
            O => \N__44454\,
            I => \c0.data_in_frame_5_0\
        );

    \I__8913\ : InMux
    port map (
            O => \N__44449\,
            I => \N__44445\
        );

    \I__8912\ : CascadeMux
    port map (
            O => \N__44448\,
            I => \N__44440\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__44445\,
            I => \N__44437\
        );

    \I__8910\ : InMux
    port map (
            O => \N__44444\,
            I => \N__44432\
        );

    \I__8909\ : InMux
    port map (
            O => \N__44443\,
            I => \N__44432\
        );

    \I__8908\ : InMux
    port map (
            O => \N__44440\,
            I => \N__44429\
        );

    \I__8907\ : Sp12to4
    port map (
            O => \N__44437\,
            I => \N__44424\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__44432\,
            I => \N__44424\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__44429\,
            I => \c0.data_in_frame_2_0\
        );

    \I__8904\ : Odrv12
    port map (
            O => \N__44424\,
            I => \c0.data_in_frame_2_0\
        );

    \I__8903\ : InMux
    port map (
            O => \N__44419\,
            I => \N__44416\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__44416\,
            I => \N__44412\
        );

    \I__8901\ : InMux
    port map (
            O => \N__44415\,
            I => \N__44409\
        );

    \I__8900\ : Span4Mux_v
    port map (
            O => \N__44412\,
            I => \N__44406\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__44409\,
            I => data_in_frame_6_1
        );

    \I__8898\ : Odrv4
    port map (
            O => \N__44406\,
            I => data_in_frame_6_1
        );

    \I__8897\ : InMux
    port map (
            O => \N__44401\,
            I => \N__44395\
        );

    \I__8896\ : InMux
    port map (
            O => \N__44400\,
            I => \N__44388\
        );

    \I__8895\ : InMux
    port map (
            O => \N__44399\,
            I => \N__44388\
        );

    \I__8894\ : InMux
    port map (
            O => \N__44398\,
            I => \N__44388\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__44395\,
            I => \c0.data_in_frame_4_7\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__44388\,
            I => \c0.data_in_frame_4_7\
        );

    \I__8891\ : CascadeMux
    port map (
            O => \N__44383\,
            I => \N__44380\
        );

    \I__8890\ : InMux
    port map (
            O => \N__44380\,
            I => \N__44375\
        );

    \I__8889\ : InMux
    port map (
            O => \N__44379\,
            I => \N__44372\
        );

    \I__8888\ : InMux
    port map (
            O => \N__44378\,
            I => \N__44369\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__44375\,
            I => \c0.data_in_frame_5_1\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__44372\,
            I => \c0.data_in_frame_5_1\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__44369\,
            I => \c0.data_in_frame_5_1\
        );

    \I__8884\ : InMux
    port map (
            O => \N__44362\,
            I => \N__44356\
        );

    \I__8883\ : InMux
    port map (
            O => \N__44361\,
            I => \N__44356\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__44356\,
            I => \N__44352\
        );

    \I__8881\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44349\
        );

    \I__8880\ : Odrv12
    port map (
            O => \N__44352\,
            I => \c0.n21992\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__44349\,
            I => \c0.n21992\
        );

    \I__8878\ : CascadeMux
    port map (
            O => \N__44344\,
            I => \N__44340\
        );

    \I__8877\ : CascadeMux
    port map (
            O => \N__44343\,
            I => \N__44337\
        );

    \I__8876\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44333\
        );

    \I__8875\ : InMux
    port map (
            O => \N__44337\,
            I => \N__44330\
        );

    \I__8874\ : InMux
    port map (
            O => \N__44336\,
            I => \N__44327\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__44333\,
            I => \c0.data_in_frame_2_2\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__44330\,
            I => \c0.data_in_frame_2_2\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__44327\,
            I => \c0.data_in_frame_2_2\
        );

    \I__8870\ : CascadeMux
    port map (
            O => \N__44320\,
            I => \N__44317\
        );

    \I__8869\ : InMux
    port map (
            O => \N__44317\,
            I => \N__44314\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__44314\,
            I => \N__44311\
        );

    \I__8867\ : Span4Mux_v
    port map (
            O => \N__44311\,
            I => \N__44305\
        );

    \I__8866\ : InMux
    port map (
            O => \N__44310\,
            I => \N__44302\
        );

    \I__8865\ : CascadeMux
    port map (
            O => \N__44309\,
            I => \N__44299\
        );

    \I__8864\ : CascadeMux
    port map (
            O => \N__44308\,
            I => \N__44294\
        );

    \I__8863\ : Span4Mux_v
    port map (
            O => \N__44305\,
            I => \N__44287\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__44302\,
            I => \N__44287\
        );

    \I__8861\ : InMux
    port map (
            O => \N__44299\,
            I => \N__44282\
        );

    \I__8860\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44282\
        );

    \I__8859\ : InMux
    port map (
            O => \N__44297\,
            I => \N__44279\
        );

    \I__8858\ : InMux
    port map (
            O => \N__44294\,
            I => \N__44272\
        );

    \I__8857\ : InMux
    port map (
            O => \N__44293\,
            I => \N__44272\
        );

    \I__8856\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44272\
        );

    \I__8855\ : Odrv4
    port map (
            O => \N__44287\,
            I => data_in_frame_1_7
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__44282\,
            I => data_in_frame_1_7
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__44279\,
            I => data_in_frame_1_7
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__44272\,
            I => data_in_frame_1_7
        );

    \I__8851\ : InMux
    port map (
            O => \N__44263\,
            I => \N__44260\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__44260\,
            I => \c0.n39_adj_4406\
        );

    \I__8849\ : CascadeMux
    port map (
            O => \N__44257\,
            I => \N__44252\
        );

    \I__8848\ : InMux
    port map (
            O => \N__44256\,
            I => \N__44248\
        );

    \I__8847\ : InMux
    port map (
            O => \N__44255\,
            I => \N__44245\
        );

    \I__8846\ : InMux
    port map (
            O => \N__44252\,
            I => \N__44242\
        );

    \I__8845\ : InMux
    port map (
            O => \N__44251\,
            I => \N__44239\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__44248\,
            I => \N__44236\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__44245\,
            I => data_in_frame_6_7
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__44242\,
            I => data_in_frame_6_7
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__44239\,
            I => data_in_frame_6_7
        );

    \I__8840\ : Odrv4
    port map (
            O => \N__44236\,
            I => data_in_frame_6_7
        );

    \I__8839\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44224\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__44224\,
            I => \c0.n21882\
        );

    \I__8837\ : InMux
    port map (
            O => \N__44221\,
            I => \N__44217\
        );

    \I__8836\ : InMux
    port map (
            O => \N__44220\,
            I => \N__44214\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__44217\,
            I => \N__44211\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__44214\,
            I => \c0.n21928\
        );

    \I__8833\ : Odrv4
    port map (
            O => \N__44211\,
            I => \c0.n21928\
        );

    \I__8832\ : CascadeMux
    port map (
            O => \N__44206\,
            I => \c0.n14037_cascade_\
        );

    \I__8831\ : InMux
    port map (
            O => \N__44203\,
            I => \N__44200\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__44200\,
            I => \c0.n6_adj_4369\
        );

    \I__8829\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44194\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__44194\,
            I => \c0.n5_adj_4368\
        );

    \I__8827\ : InMux
    port map (
            O => \N__44191\,
            I => \N__44188\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__44188\,
            I => \c0.data_out_frame_29__7__N_1474\
        );

    \I__8825\ : CascadeMux
    port map (
            O => \N__44185\,
            I => \N__44182\
        );

    \I__8824\ : InMux
    port map (
            O => \N__44182\,
            I => \N__44178\
        );

    \I__8823\ : InMux
    port map (
            O => \N__44181\,
            I => \N__44175\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__44178\,
            I => \N__44172\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__44175\,
            I => data_in_frame_6_6
        );

    \I__8820\ : Odrv4
    port map (
            O => \N__44172\,
            I => data_in_frame_6_6
        );

    \I__8819\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44162\
        );

    \I__8818\ : InMux
    port map (
            O => \N__44166\,
            I => \N__44159\
        );

    \I__8817\ : InMux
    port map (
            O => \N__44165\,
            I => \N__44156\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__44162\,
            I => \N__44153\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__44159\,
            I => \N__44150\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__44156\,
            I => \N__44147\
        );

    \I__8813\ : Span4Mux_h
    port map (
            O => \N__44153\,
            I => \N__44142\
        );

    \I__8812\ : Span4Mux_v
    port map (
            O => \N__44150\,
            I => \N__44137\
        );

    \I__8811\ : Span4Mux_h
    port map (
            O => \N__44147\,
            I => \N__44137\
        );

    \I__8810\ : CascadeMux
    port map (
            O => \N__44146\,
            I => \N__44132\
        );

    \I__8809\ : InMux
    port map (
            O => \N__44145\,
            I => \N__44129\
        );

    \I__8808\ : Span4Mux_v
    port map (
            O => \N__44142\,
            I => \N__44126\
        );

    \I__8807\ : Span4Mux_v
    port map (
            O => \N__44137\,
            I => \N__44123\
        );

    \I__8806\ : InMux
    port map (
            O => \N__44136\,
            I => \N__44120\
        );

    \I__8805\ : InMux
    port map (
            O => \N__44135\,
            I => \N__44115\
        );

    \I__8804\ : InMux
    port map (
            O => \N__44132\,
            I => \N__44115\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__44129\,
            I => \c0.data_in_frame_0_2\
        );

    \I__8802\ : Odrv4
    port map (
            O => \N__44126\,
            I => \c0.data_in_frame_0_2\
        );

    \I__8801\ : Odrv4
    port map (
            O => \N__44123\,
            I => \c0.data_in_frame_0_2\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__44120\,
            I => \c0.data_in_frame_0_2\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__44115\,
            I => \c0.data_in_frame_0_2\
        );

    \I__8798\ : CascadeMux
    port map (
            O => \N__44104\,
            I => \N__44100\
        );

    \I__8797\ : InMux
    port map (
            O => \N__44103\,
            I => \N__44096\
        );

    \I__8796\ : InMux
    port map (
            O => \N__44100\,
            I => \N__44093\
        );

    \I__8795\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44090\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__44096\,
            I => \N__44087\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__44093\,
            I => \c0.data_in_frame_3_6\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__44090\,
            I => \c0.data_in_frame_3_6\
        );

    \I__8791\ : Odrv4
    port map (
            O => \N__44087\,
            I => \c0.data_in_frame_3_6\
        );

    \I__8790\ : InMux
    port map (
            O => \N__44080\,
            I => \N__44073\
        );

    \I__8789\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44073\
        );

    \I__8788\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44070\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__44073\,
            I => \c0.data_in_frame_4_1\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__44070\,
            I => \c0.data_in_frame_4_1\
        );

    \I__8785\ : InMux
    port map (
            O => \N__44065\,
            I => \N__44061\
        );

    \I__8784\ : InMux
    port map (
            O => \N__44064\,
            I => \N__44058\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__44061\,
            I => \c0.n22218\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__44058\,
            I => \c0.n22218\
        );

    \I__8781\ : CascadeMux
    port map (
            O => \N__44053\,
            I => \c0.n21928_cascade_\
        );

    \I__8780\ : InMux
    port map (
            O => \N__44050\,
            I => \N__44045\
        );

    \I__8779\ : CascadeMux
    port map (
            O => \N__44049\,
            I => \N__44042\
        );

    \I__8778\ : CascadeMux
    port map (
            O => \N__44048\,
            I => \N__44039\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__44045\,
            I => \N__44035\
        );

    \I__8776\ : InMux
    port map (
            O => \N__44042\,
            I => \N__44032\
        );

    \I__8775\ : InMux
    port map (
            O => \N__44039\,
            I => \N__44029\
        );

    \I__8774\ : InMux
    port map (
            O => \N__44038\,
            I => \N__44026\
        );

    \I__8773\ : Span4Mux_h
    port map (
            O => \N__44035\,
            I => \N__44021\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__44032\,
            I => \N__44021\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__44029\,
            I => \c0.data_in_frame_2_3\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__44026\,
            I => \c0.data_in_frame_2_3\
        );

    \I__8769\ : Odrv4
    port map (
            O => \N__44021\,
            I => \c0.data_in_frame_2_3\
        );

    \I__8768\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44009\
        );

    \I__8767\ : InMux
    port map (
            O => \N__44013\,
            I => \N__44006\
        );

    \I__8766\ : InMux
    port map (
            O => \N__44012\,
            I => \N__44003\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__44009\,
            I => \N__44000\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__44006\,
            I => \c0.n21791\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__44003\,
            I => \c0.n21791\
        );

    \I__8762\ : Odrv4
    port map (
            O => \N__44000\,
            I => \c0.n21791\
        );

    \I__8761\ : CascadeMux
    port map (
            O => \N__43993\,
            I => \c0.n21882_cascade_\
        );

    \I__8760\ : InMux
    port map (
            O => \N__43990\,
            I => \N__43987\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__43987\,
            I => \N__43984\
        );

    \I__8758\ : Span4Mux_v
    port map (
            O => \N__43984\,
            I => \N__43981\
        );

    \I__8757\ : Odrv4
    port map (
            O => \N__43981\,
            I => \c0.data_out_frame_0__7__N_2744\
        );

    \I__8756\ : CascadeMux
    port map (
            O => \N__43978\,
            I => \c0.data_out_frame_0__7__N_2744_cascade_\
        );

    \I__8755\ : CascadeMux
    port map (
            O => \N__43975\,
            I => \c0.n6_adj_4272_cascade_\
        );

    \I__8754\ : CascadeMux
    port map (
            O => \N__43972\,
            I => \N__43967\
        );

    \I__8753\ : InMux
    port map (
            O => \N__43971\,
            I => \N__43962\
        );

    \I__8752\ : InMux
    port map (
            O => \N__43970\,
            I => \N__43962\
        );

    \I__8751\ : InMux
    port map (
            O => \N__43967\,
            I => \N__43959\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__43962\,
            I => \N__43956\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__43959\,
            I => \c0.data_in_frame_3_7\
        );

    \I__8748\ : Odrv4
    port map (
            O => \N__43956\,
            I => \c0.data_in_frame_3_7\
        );

    \I__8747\ : InMux
    port map (
            O => \N__43951\,
            I => \N__43948\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__43948\,
            I => \c0.n21803\
        );

    \I__8745\ : InMux
    port map (
            O => \N__43945\,
            I => \N__43942\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__43942\,
            I => \N__43939\
        );

    \I__8743\ : Odrv12
    port map (
            O => \N__43939\,
            I => \c0.n18_adj_4370\
        );

    \I__8742\ : InMux
    port map (
            O => \N__43936\,
            I => \N__43933\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__43933\,
            I => \c0.n22194\
        );

    \I__8740\ : CascadeMux
    port map (
            O => \N__43930\,
            I => \c0.n21803_cascade_\
        );

    \I__8739\ : InMux
    port map (
            O => \N__43927\,
            I => \N__43924\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__43924\,
            I => \c0.n30_adj_4371\
        );

    \I__8737\ : InMux
    port map (
            O => \N__43921\,
            I => \N__43915\
        );

    \I__8736\ : InMux
    port map (
            O => \N__43920\,
            I => \N__43910\
        );

    \I__8735\ : InMux
    port map (
            O => \N__43919\,
            I => \N__43910\
        );

    \I__8734\ : InMux
    port map (
            O => \N__43918\,
            I => \N__43907\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__43915\,
            I => \N__43904\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__43910\,
            I => \N__43901\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__43907\,
            I => \N__43892\
        );

    \I__8730\ : Span4Mux_v
    port map (
            O => \N__43904\,
            I => \N__43892\
        );

    \I__8729\ : Span4Mux_h
    port map (
            O => \N__43901\,
            I => \N__43892\
        );

    \I__8728\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43889\
        );

    \I__8727\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43886\
        );

    \I__8726\ : Odrv4
    port map (
            O => \N__43892\,
            I => \c0.data_in_frame_0_1\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__43889\,
            I => \c0.data_in_frame_0_1\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__43886\,
            I => \c0.data_in_frame_0_1\
        );

    \I__8723\ : CascadeMux
    port map (
            O => \N__43879\,
            I => \N__43875\
        );

    \I__8722\ : InMux
    port map (
            O => \N__43878\,
            I => \N__43872\
        );

    \I__8721\ : InMux
    port map (
            O => \N__43875\,
            I => \N__43865\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__43872\,
            I => \N__43862\
        );

    \I__8719\ : InMux
    port map (
            O => \N__43871\,
            I => \N__43859\
        );

    \I__8718\ : InMux
    port map (
            O => \N__43870\,
            I => \N__43856\
        );

    \I__8717\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43851\
        );

    \I__8716\ : InMux
    port map (
            O => \N__43868\,
            I => \N__43851\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__43865\,
            I => \N__43848\
        );

    \I__8714\ : Odrv12
    port map (
            O => \N__43862\,
            I => \c0.data_in_frame_0_0\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__43859\,
            I => \c0.data_in_frame_0_0\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__43856\,
            I => \c0.data_in_frame_0_0\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__43851\,
            I => \c0.data_in_frame_0_0\
        );

    \I__8710\ : Odrv4
    port map (
            O => \N__43848\,
            I => \c0.data_in_frame_0_0\
        );

    \I__8709\ : CascadeMux
    port map (
            O => \N__43837\,
            I => \c0.n13376_cascade_\
        );

    \I__8708\ : InMux
    port map (
            O => \N__43834\,
            I => \N__43830\
        );

    \I__8707\ : InMux
    port map (
            O => \N__43833\,
            I => \N__43827\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__43830\,
            I => \c0.n13376\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__43827\,
            I => \c0.n13376\
        );

    \I__8704\ : InMux
    port map (
            O => \N__43822\,
            I => \N__43819\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__43819\,
            I => \N__43814\
        );

    \I__8702\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43811\
        );

    \I__8701\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43803\
        );

    \I__8700\ : Span4Mux_v
    port map (
            O => \N__43814\,
            I => \N__43800\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__43811\,
            I => \N__43797\
        );

    \I__8698\ : InMux
    port map (
            O => \N__43810\,
            I => \N__43794\
        );

    \I__8697\ : InMux
    port map (
            O => \N__43809\,
            I => \N__43791\
        );

    \I__8696\ : InMux
    port map (
            O => \N__43808\,
            I => \N__43784\
        );

    \I__8695\ : InMux
    port map (
            O => \N__43807\,
            I => \N__43784\
        );

    \I__8694\ : InMux
    port map (
            O => \N__43806\,
            I => \N__43784\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__43803\,
            I => data_in_frame_1_6
        );

    \I__8692\ : Odrv4
    port map (
            O => \N__43800\,
            I => data_in_frame_1_6
        );

    \I__8691\ : Odrv12
    port map (
            O => \N__43797\,
            I => data_in_frame_1_6
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__43794\,
            I => data_in_frame_1_6
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__43791\,
            I => data_in_frame_1_6
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__43784\,
            I => data_in_frame_1_6
        );

    \I__8687\ : InMux
    port map (
            O => \N__43771\,
            I => \N__43767\
        );

    \I__8686\ : InMux
    port map (
            O => \N__43770\,
            I => \N__43764\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__43767\,
            I => data_in_frame_6_2
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__43764\,
            I => data_in_frame_6_2
        );

    \I__8683\ : CascadeMux
    port map (
            O => \N__43759\,
            I => \c0.n13386_cascade_\
        );

    \I__8682\ : CascadeMux
    port map (
            O => \N__43756\,
            I => \N__43753\
        );

    \I__8681\ : InMux
    port map (
            O => \N__43753\,
            I => \N__43748\
        );

    \I__8680\ : InMux
    port map (
            O => \N__43752\,
            I => \N__43745\
        );

    \I__8679\ : InMux
    port map (
            O => \N__43751\,
            I => \N__43742\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__43748\,
            I => \c0.data_in_frame_4_4\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__43745\,
            I => \c0.data_in_frame_4_4\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__43742\,
            I => \c0.data_in_frame_4_4\
        );

    \I__8675\ : InMux
    port map (
            O => \N__43735\,
            I => \N__43732\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__43732\,
            I => \c0.n22261\
        );

    \I__8673\ : CascadeMux
    port map (
            O => \N__43729\,
            I => \N__43725\
        );

    \I__8672\ : InMux
    port map (
            O => \N__43728\,
            I => \N__43720\
        );

    \I__8671\ : InMux
    port map (
            O => \N__43725\,
            I => \N__43715\
        );

    \I__8670\ : InMux
    port map (
            O => \N__43724\,
            I => \N__43715\
        );

    \I__8669\ : InMux
    port map (
            O => \N__43723\,
            I => \N__43712\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__43720\,
            I => \c0.data_in_frame_2_1\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__43715\,
            I => \c0.data_in_frame_2_1\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__43712\,
            I => \c0.data_in_frame_2_1\
        );

    \I__8665\ : CascadeMux
    port map (
            O => \N__43705\,
            I => \c0.n22261_cascade_\
        );

    \I__8664\ : InMux
    port map (
            O => \N__43702\,
            I => \N__43699\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__43699\,
            I => \c0.n22320\
        );

    \I__8662\ : InMux
    port map (
            O => \N__43696\,
            I => \N__43693\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__43693\,
            I => \c0.n28_adj_4372\
        );

    \I__8660\ : InMux
    port map (
            O => \N__43690\,
            I => \N__43687\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__43687\,
            I => \c0.n22290\
        );

    \I__8658\ : CascadeMux
    port map (
            O => \N__43684\,
            I => \N__43681\
        );

    \I__8657\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43678\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__43678\,
            I => \c0.n22258\
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__43675\,
            I => \c0.n22258_cascade_\
        );

    \I__8654\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43669\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__43669\,
            I => \c0.n29_adj_4374\
        );

    \I__8652\ : CascadeMux
    port map (
            O => \N__43666\,
            I => \c0.n27_adj_4377_cascade_\
        );

    \I__8651\ : CascadeMux
    port map (
            O => \N__43663\,
            I => \c0.n14072_cascade_\
        );

    \I__8650\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43657\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__43657\,
            I => \c0.n14072\
        );

    \I__8648\ : CascadeMux
    port map (
            O => \N__43654\,
            I => \c0.n6_adj_4385_cascade_\
        );

    \I__8647\ : CascadeMux
    port map (
            O => \N__43651\,
            I => \c0.n21902_cascade_\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__43648\,
            I => \N__43645\
        );

    \I__8645\ : InMux
    port map (
            O => \N__43645\,
            I => \N__43639\
        );

    \I__8644\ : InMux
    port map (
            O => \N__43644\,
            I => \N__43639\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__43639\,
            I => \c0.data_in_frame_3_0\
        );

    \I__8642\ : InMux
    port map (
            O => \N__43636\,
            I => \N__43633\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__43633\,
            I => \c0.n21902\
        );

    \I__8640\ : CascadeMux
    port map (
            O => \N__43630\,
            I => \N__43626\
        );

    \I__8639\ : CascadeMux
    port map (
            O => \N__43629\,
            I => \N__43623\
        );

    \I__8638\ : InMux
    port map (
            O => \N__43626\,
            I => \N__43620\
        );

    \I__8637\ : InMux
    port map (
            O => \N__43623\,
            I => \N__43617\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__43620\,
            I => \c0.data_in_frame_5_2\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__43617\,
            I => \c0.data_in_frame_5_2\
        );

    \I__8634\ : CascadeMux
    port map (
            O => \N__43612\,
            I => \c0.n21879_cascade_\
        );

    \I__8633\ : CascadeMux
    port map (
            O => \N__43609\,
            I => \N__43606\
        );

    \I__8632\ : InMux
    port map (
            O => \N__43606\,
            I => \N__43599\
        );

    \I__8631\ : InMux
    port map (
            O => \N__43605\,
            I => \N__43599\
        );

    \I__8630\ : InMux
    port map (
            O => \N__43604\,
            I => \N__43596\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__43599\,
            I => \c0.data_in_frame_3_4\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__43596\,
            I => \c0.data_in_frame_3_4\
        );

    \I__8627\ : InMux
    port map (
            O => \N__43591\,
            I => \N__43588\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__43588\,
            I => \N__43585\
        );

    \I__8625\ : Odrv4
    port map (
            O => \N__43585\,
            I => \c0.n21957\
        );

    \I__8624\ : CascadeMux
    port map (
            O => \N__43582\,
            I => \c0.n21957_cascade_\
        );

    \I__8623\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43576\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__43576\,
            I => \c0.n22287\
        );

    \I__8621\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43564\
        );

    \I__8620\ : InMux
    port map (
            O => \N__43572\,
            I => \N__43564\
        );

    \I__8619\ : InMux
    port map (
            O => \N__43571\,
            I => \N__43564\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__43564\,
            I => \c0.data_in_frame_3_3\
        );

    \I__8617\ : CascadeMux
    port map (
            O => \N__43561\,
            I => \N__43558\
        );

    \I__8616\ : InMux
    port map (
            O => \N__43558\,
            I => \N__43552\
        );

    \I__8615\ : InMux
    port map (
            O => \N__43557\,
            I => \N__43552\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__43552\,
            I => \c0.data_in_frame_5_4\
        );

    \I__8613\ : InMux
    port map (
            O => \N__43549\,
            I => \N__43546\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__43546\,
            I => \N__43543\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__43543\,
            I => \c0.n23838\
        );

    \I__8610\ : InMux
    port map (
            O => \N__43540\,
            I => \N__43536\
        );

    \I__8609\ : InMux
    port map (
            O => \N__43539\,
            I => \N__43533\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__43536\,
            I => \N__43526\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__43533\,
            I => \N__43526\
        );

    \I__8606\ : InMux
    port map (
            O => \N__43532\,
            I => \N__43523\
        );

    \I__8605\ : InMux
    port map (
            O => \N__43531\,
            I => \N__43520\
        );

    \I__8604\ : Span4Mux_h
    port map (
            O => \N__43526\,
            I => \N__43517\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__43523\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__43520\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__8601\ : Odrv4
    port map (
            O => \N__43517\,
            I => \c0.FRAME_MATCHER_state_28\
        );

    \I__8600\ : SRMux
    port map (
            O => \N__43510\,
            I => \N__43507\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__43507\,
            I => \c0.n21378\
        );

    \I__8598\ : InMux
    port map (
            O => \N__43504\,
            I => \N__43499\
        );

    \I__8597\ : InMux
    port map (
            O => \N__43503\,
            I => \N__43496\
        );

    \I__8596\ : CascadeMux
    port map (
            O => \N__43502\,
            I => \N__43493\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__43499\,
            I => \N__43488\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__43496\,
            I => \N__43488\
        );

    \I__8593\ : InMux
    port map (
            O => \N__43493\,
            I => \N__43484\
        );

    \I__8592\ : Span4Mux_v
    port map (
            O => \N__43488\,
            I => \N__43481\
        );

    \I__8591\ : InMux
    port map (
            O => \N__43487\,
            I => \N__43478\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__43484\,
            I => \N__43475\
        );

    \I__8589\ : Span4Mux_h
    port map (
            O => \N__43481\,
            I => \N__43472\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__43478\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__8587\ : Odrv4
    port map (
            O => \N__43475\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__8586\ : Odrv4
    port map (
            O => \N__43472\,
            I => \c0.FRAME_MATCHER_state_31\
        );

    \I__8585\ : SRMux
    port map (
            O => \N__43465\,
            I => \N__43462\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__43462\,
            I => \N__43459\
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__43459\,
            I => \c0.n21332\
        );

    \I__8582\ : CascadeMux
    port map (
            O => \N__43456\,
            I => \N__43452\
        );

    \I__8581\ : InMux
    port map (
            O => \N__43455\,
            I => \N__43448\
        );

    \I__8580\ : InMux
    port map (
            O => \N__43452\,
            I => \N__43445\
        );

    \I__8579\ : InMux
    port map (
            O => \N__43451\,
            I => \N__43441\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__43448\,
            I => \N__43436\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__43445\,
            I => \N__43436\
        );

    \I__8576\ : InMux
    port map (
            O => \N__43444\,
            I => \N__43433\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__43441\,
            I => \N__43430\
        );

    \I__8574\ : Span4Mux_h
    port map (
            O => \N__43436\,
            I => \N__43427\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__43433\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__8572\ : Odrv12
    port map (
            O => \N__43430\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__8571\ : Odrv4
    port map (
            O => \N__43427\,
            I => \c0.FRAME_MATCHER_state_13\
        );

    \I__8570\ : SRMux
    port map (
            O => \N__43420\,
            I => \N__43417\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__43417\,
            I => \N__43414\
        );

    \I__8568\ : Odrv4
    port map (
            O => \N__43414\,
            I => \c0.n21354\
        );

    \I__8567\ : InMux
    port map (
            O => \N__43411\,
            I => \N__43407\
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__43410\,
            I => \N__43404\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__43407\,
            I => \N__43401\
        );

    \I__8564\ : InMux
    port map (
            O => \N__43404\,
            I => \N__43398\
        );

    \I__8563\ : Span4Mux_h
    port map (
            O => \N__43401\,
            I => \N__43395\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__43398\,
            I => \N__43388\
        );

    \I__8561\ : Span4Mux_v
    port map (
            O => \N__43395\,
            I => \N__43388\
        );

    \I__8560\ : InMux
    port map (
            O => \N__43394\,
            I => \N__43385\
        );

    \I__8559\ : InMux
    port map (
            O => \N__43393\,
            I => \N__43382\
        );

    \I__8558\ : Span4Mux_h
    port map (
            O => \N__43388\,
            I => \N__43379\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__43385\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__43382\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__8555\ : Odrv4
    port map (
            O => \N__43379\,
            I => \c0.FRAME_MATCHER_state_15\
        );

    \I__8554\ : SRMux
    port map (
            O => \N__43372\,
            I => \N__43369\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__43369\,
            I => \N__43366\
        );

    \I__8552\ : Odrv4
    port map (
            O => \N__43366\,
            I => \c0.n21358\
        );

    \I__8551\ : InMux
    port map (
            O => \N__43363\,
            I => \N__43358\
        );

    \I__8550\ : InMux
    port map (
            O => \N__43362\,
            I => \N__43353\
        );

    \I__8549\ : InMux
    port map (
            O => \N__43361\,
            I => \N__43353\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__43358\,
            I => \N__43350\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__43353\,
            I => \c0.n21734\
        );

    \I__8546\ : Odrv4
    port map (
            O => \N__43350\,
            I => \c0.n21734\
        );

    \I__8545\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43333\
        );

    \I__8544\ : InMux
    port map (
            O => \N__43344\,
            I => \N__43333\
        );

    \I__8543\ : InMux
    port map (
            O => \N__43343\,
            I => \N__43333\
        );

    \I__8542\ : InMux
    port map (
            O => \N__43342\,
            I => \N__43330\
        );

    \I__8541\ : InMux
    port map (
            O => \N__43341\,
            I => \N__43325\
        );

    \I__8540\ : InMux
    port map (
            O => \N__43340\,
            I => \N__43325\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__43333\,
            I => \N__43322\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__43330\,
            I => \N__43319\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__43325\,
            I => \N__43314\
        );

    \I__8536\ : Span4Mux_h
    port map (
            O => \N__43322\,
            I => \N__43314\
        );

    \I__8535\ : Span4Mux_h
    port map (
            O => \N__43319\,
            I => \N__43311\
        );

    \I__8534\ : Odrv4
    port map (
            O => \N__43314\,
            I => \c0.n13021\
        );

    \I__8533\ : Odrv4
    port map (
            O => \N__43311\,
            I => \c0.n13021\
        );

    \I__8532\ : CascadeMux
    port map (
            O => \N__43306\,
            I => \N__43303\
        );

    \I__8531\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43300\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__43300\,
            I => \N__43297\
        );

    \I__8529\ : Span4Mux_h
    port map (
            O => \N__43297\,
            I => \N__43294\
        );

    \I__8528\ : Odrv4
    port map (
            O => \N__43294\,
            I => \c0.n23965\
        );

    \I__8527\ : InMux
    port map (
            O => \N__43291\,
            I => \N__43287\
        );

    \I__8526\ : InMux
    port map (
            O => \N__43290\,
            I => \N__43284\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__43287\,
            I => \c0.n22575\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__43284\,
            I => \c0.n22575\
        );

    \I__8523\ : InMux
    port map (
            O => \N__43279\,
            I => \N__43276\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__43276\,
            I => \c0.n45_adj_4389\
        );

    \I__8521\ : CascadeMux
    port map (
            O => \N__43273\,
            I => \N__43270\
        );

    \I__8520\ : InMux
    port map (
            O => \N__43270\,
            I => \N__43251\
        );

    \I__8519\ : InMux
    port map (
            O => \N__43269\,
            I => \N__43251\
        );

    \I__8518\ : InMux
    port map (
            O => \N__43268\,
            I => \N__43251\
        );

    \I__8517\ : InMux
    port map (
            O => \N__43267\,
            I => \N__43246\
        );

    \I__8516\ : InMux
    port map (
            O => \N__43266\,
            I => \N__43246\
        );

    \I__8515\ : CascadeMux
    port map (
            O => \N__43265\,
            I => \N__43240\
        );

    \I__8514\ : InMux
    port map (
            O => \N__43264\,
            I => \N__43236\
        );

    \I__8513\ : InMux
    port map (
            O => \N__43263\,
            I => \N__43233\
        );

    \I__8512\ : InMux
    port map (
            O => \N__43262\,
            I => \N__43230\
        );

    \I__8511\ : InMux
    port map (
            O => \N__43261\,
            I => \N__43227\
        );

    \I__8510\ : InMux
    port map (
            O => \N__43260\,
            I => \N__43220\
        );

    \I__8509\ : InMux
    port map (
            O => \N__43259\,
            I => \N__43220\
        );

    \I__8508\ : InMux
    port map (
            O => \N__43258\,
            I => \N__43220\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__43251\,
            I => \N__43210\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__43246\,
            I => \N__43210\
        );

    \I__8505\ : InMux
    port map (
            O => \N__43245\,
            I => \N__43199\
        );

    \I__8504\ : InMux
    port map (
            O => \N__43244\,
            I => \N__43199\
        );

    \I__8503\ : InMux
    port map (
            O => \N__43243\,
            I => \N__43199\
        );

    \I__8502\ : InMux
    port map (
            O => \N__43240\,
            I => \N__43199\
        );

    \I__8501\ : InMux
    port map (
            O => \N__43239\,
            I => \N__43199\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__43236\,
            I => \N__43194\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__43233\,
            I => \N__43194\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__43230\,
            I => \N__43185\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__43227\,
            I => \N__43185\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__43220\,
            I => \N__43185\
        );

    \I__8495\ : InMux
    port map (
            O => \N__43219\,
            I => \N__43182\
        );

    \I__8494\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43179\
        );

    \I__8493\ : InMux
    port map (
            O => \N__43217\,
            I => \N__43176\
        );

    \I__8492\ : InMux
    port map (
            O => \N__43216\,
            I => \N__43172\
        );

    \I__8491\ : InMux
    port map (
            O => \N__43215\,
            I => \N__43166\
        );

    \I__8490\ : Span4Mux_v
    port map (
            O => \N__43210\,
            I => \N__43161\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__43199\,
            I => \N__43161\
        );

    \I__8488\ : Span4Mux_v
    port map (
            O => \N__43194\,
            I => \N__43158\
        );

    \I__8487\ : InMux
    port map (
            O => \N__43193\,
            I => \N__43151\
        );

    \I__8486\ : InMux
    port map (
            O => \N__43192\,
            I => \N__43148\
        );

    \I__8485\ : Span4Mux_v
    port map (
            O => \N__43185\,
            I => \N__43139\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__43182\,
            I => \N__43139\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__43179\,
            I => \N__43139\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__43176\,
            I => \N__43139\
        );

    \I__8481\ : InMux
    port map (
            O => \N__43175\,
            I => \N__43136\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__43172\,
            I => \N__43133\
        );

    \I__8479\ : InMux
    port map (
            O => \N__43171\,
            I => \N__43130\
        );

    \I__8478\ : InMux
    port map (
            O => \N__43170\,
            I => \N__43125\
        );

    \I__8477\ : InMux
    port map (
            O => \N__43169\,
            I => \N__43125\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__43166\,
            I => \N__43120\
        );

    \I__8475\ : Span4Mux_h
    port map (
            O => \N__43161\,
            I => \N__43120\
        );

    \I__8474\ : Sp12to4
    port map (
            O => \N__43158\,
            I => \N__43117\
        );

    \I__8473\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43112\
        );

    \I__8472\ : InMux
    port map (
            O => \N__43156\,
            I => \N__43112\
        );

    \I__8471\ : InMux
    port map (
            O => \N__43155\,
            I => \N__43106\
        );

    \I__8470\ : InMux
    port map (
            O => \N__43154\,
            I => \N__43103\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__43151\,
            I => \N__43096\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__43148\,
            I => \N__43096\
        );

    \I__8467\ : Span4Mux_h
    port map (
            O => \N__43139\,
            I => \N__43096\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__43136\,
            I => \N__43091\
        );

    \I__8465\ : Span4Mux_v
    port map (
            O => \N__43133\,
            I => \N__43091\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__43130\,
            I => \N__43080\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__43125\,
            I => \N__43080\
        );

    \I__8462\ : Sp12to4
    port map (
            O => \N__43120\,
            I => \N__43080\
        );

    \I__8461\ : Span12Mux_h
    port map (
            O => \N__43117\,
            I => \N__43080\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__43112\,
            I => \N__43080\
        );

    \I__8459\ : InMux
    port map (
            O => \N__43111\,
            I => \N__43072\
        );

    \I__8458\ : InMux
    port map (
            O => \N__43110\,
            I => \N__43072\
        );

    \I__8457\ : InMux
    port map (
            O => \N__43109\,
            I => \N__43072\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__43106\,
            I => \N__43067\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__43103\,
            I => \N__43067\
        );

    \I__8454\ : Span4Mux_v
    port map (
            O => \N__43096\,
            I => \N__43064\
        );

    \I__8453\ : Sp12to4
    port map (
            O => \N__43091\,
            I => \N__43059\
        );

    \I__8452\ : Span12Mux_v
    port map (
            O => \N__43080\,
            I => \N__43059\
        );

    \I__8451\ : InMux
    port map (
            O => \N__43079\,
            I => \N__43056\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__43072\,
            I => rx_data_ready
        );

    \I__8449\ : Odrv12
    port map (
            O => \N__43067\,
            I => rx_data_ready
        );

    \I__8448\ : Odrv4
    port map (
            O => \N__43064\,
            I => rx_data_ready
        );

    \I__8447\ : Odrv12
    port map (
            O => \N__43059\,
            I => rx_data_ready
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__43056\,
            I => rx_data_ready
        );

    \I__8445\ : InMux
    port map (
            O => \N__43045\,
            I => \N__43038\
        );

    \I__8444\ : InMux
    port map (
            O => \N__43044\,
            I => \N__43038\
        );

    \I__8443\ : InMux
    port map (
            O => \N__43043\,
            I => \N__43035\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__43038\,
            I => \N__43032\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__43035\,
            I => \N__43028\
        );

    \I__8440\ : Span4Mux_h
    port map (
            O => \N__43032\,
            I => \N__43025\
        );

    \I__8439\ : InMux
    port map (
            O => \N__43031\,
            I => \N__43022\
        );

    \I__8438\ : Span4Mux_v
    port map (
            O => \N__43028\,
            I => \N__43019\
        );

    \I__8437\ : Span4Mux_h
    port map (
            O => \N__43025\,
            I => \N__43016\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__43022\,
            I => data_in_3_1
        );

    \I__8435\ : Odrv4
    port map (
            O => \N__43019\,
            I => data_in_3_1
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__43016\,
            I => data_in_3_1
        );

    \I__8433\ : InMux
    port map (
            O => \N__43009\,
            I => \N__43004\
        );

    \I__8432\ : InMux
    port map (
            O => \N__43008\,
            I => \N__43001\
        );

    \I__8431\ : InMux
    port map (
            O => \N__43007\,
            I => \N__42998\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__43004\,
            I => \N__42995\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__43001\,
            I => \N__42990\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__42998\,
            I => \N__42990\
        );

    \I__8427\ : Odrv4
    port map (
            O => \N__42995\,
            I => \c0.n1\
        );

    \I__8426\ : Odrv12
    port map (
            O => \N__42990\,
            I => \c0.n1\
        );

    \I__8425\ : InMux
    port map (
            O => \N__42985\,
            I => \N__42982\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__42982\,
            I => \N__42979\
        );

    \I__8423\ : Span4Mux_v
    port map (
            O => \N__42979\,
            I => \N__42975\
        );

    \I__8422\ : InMux
    port map (
            O => \N__42978\,
            I => \N__42972\
        );

    \I__8421\ : Span4Mux_h
    port map (
            O => \N__42975\,
            I => \N__42966\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__42972\,
            I => \N__42966\
        );

    \I__8419\ : InMux
    port map (
            O => \N__42971\,
            I => \N__42963\
        );

    \I__8418\ : Sp12to4
    port map (
            O => \N__42966\,
            I => \N__42958\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__42963\,
            I => \N__42958\
        );

    \I__8416\ : Odrv12
    port map (
            O => \N__42958\,
            I => \c0.n19783\
        );

    \I__8415\ : InMux
    port map (
            O => \N__42955\,
            I => \N__42951\
        );

    \I__8414\ : InMux
    port map (
            O => \N__42954\,
            I => \N__42948\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__42951\,
            I => \N__42943\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__42948\,
            I => \N__42943\
        );

    \I__8411\ : Span4Mux_h
    port map (
            O => \N__42943\,
            I => \N__42940\
        );

    \I__8410\ : Odrv4
    port map (
            O => \N__42940\,
            I => \c0.n937\
        );

    \I__8409\ : InMux
    port map (
            O => \N__42937\,
            I => \N__42932\
        );

    \I__8408\ : CascadeMux
    port map (
            O => \N__42936\,
            I => \N__42929\
        );

    \I__8407\ : InMux
    port map (
            O => \N__42935\,
            I => \N__42925\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__42932\,
            I => \N__42922\
        );

    \I__8405\ : InMux
    port map (
            O => \N__42929\,
            I => \N__42919\
        );

    \I__8404\ : InMux
    port map (
            O => \N__42928\,
            I => \N__42916\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__42925\,
            I => \N__42913\
        );

    \I__8402\ : Span4Mux_h
    port map (
            O => \N__42922\,
            I => \N__42910\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__42919\,
            I => \N__42907\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__42916\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__8399\ : Odrv4
    port map (
            O => \N__42913\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__8398\ : Odrv4
    port map (
            O => \N__42910\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__8397\ : Odrv12
    port map (
            O => \N__42907\,
            I => \c0.FRAME_MATCHER_state_12\
        );

    \I__8396\ : SRMux
    port map (
            O => \N__42898\,
            I => \N__42895\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__42895\,
            I => \N__42892\
        );

    \I__8394\ : Span4Mux_h
    port map (
            O => \N__42892\,
            I => \N__42889\
        );

    \I__8393\ : Odrv4
    port map (
            O => \N__42889\,
            I => \c0.n21352\
        );

    \I__8392\ : CascadeMux
    port map (
            O => \N__42886\,
            I => \N__42881\
        );

    \I__8391\ : InMux
    port map (
            O => \N__42885\,
            I => \N__42877\
        );

    \I__8390\ : InMux
    port map (
            O => \N__42884\,
            I => \N__42874\
        );

    \I__8389\ : InMux
    port map (
            O => \N__42881\,
            I => \N__42871\
        );

    \I__8388\ : InMux
    port map (
            O => \N__42880\,
            I => \N__42867\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__42877\,
            I => \N__42864\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__42874\,
            I => \N__42859\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__42871\,
            I => \N__42859\
        );

    \I__8384\ : InMux
    port map (
            O => \N__42870\,
            I => \N__42856\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__42867\,
            I => \N__42853\
        );

    \I__8382\ : Span4Mux_v
    port map (
            O => \N__42864\,
            I => \N__42850\
        );

    \I__8381\ : Span4Mux_v
    port map (
            O => \N__42859\,
            I => \N__42847\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__42856\,
            I => \N__42844\
        );

    \I__8379\ : Odrv12
    port map (
            O => \N__42853\,
            I => \c0.n20_adj_4327\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__42850\,
            I => \c0.n20_adj_4327\
        );

    \I__8377\ : Odrv4
    port map (
            O => \N__42847\,
            I => \c0.n20_adj_4327\
        );

    \I__8376\ : Odrv12
    port map (
            O => \N__42844\,
            I => \c0.n20_adj_4327\
        );

    \I__8375\ : InMux
    port map (
            O => \N__42835\,
            I => \N__42830\
        );

    \I__8374\ : InMux
    port map (
            O => \N__42834\,
            I => \N__42827\
        );

    \I__8373\ : InMux
    port map (
            O => \N__42833\,
            I => \N__42822\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__42830\,
            I => \N__42819\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__42827\,
            I => \N__42816\
        );

    \I__8370\ : InMux
    port map (
            O => \N__42826\,
            I => \N__42813\
        );

    \I__8369\ : InMux
    port map (
            O => \N__42825\,
            I => \N__42810\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__42822\,
            I => \c0.n12992\
        );

    \I__8367\ : Odrv4
    port map (
            O => \N__42819\,
            I => \c0.n12992\
        );

    \I__8366\ : Odrv12
    port map (
            O => \N__42816\,
            I => \c0.n12992\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__42813\,
            I => \c0.n12992\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__42810\,
            I => \c0.n12992\
        );

    \I__8363\ : InMux
    port map (
            O => \N__42799\,
            I => \N__42782\
        );

    \I__8362\ : InMux
    port map (
            O => \N__42798\,
            I => \N__42779\
        );

    \I__8361\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42770\
        );

    \I__8360\ : InMux
    port map (
            O => \N__42796\,
            I => \N__42770\
        );

    \I__8359\ : InMux
    port map (
            O => \N__42795\,
            I => \N__42770\
        );

    \I__8358\ : InMux
    port map (
            O => \N__42794\,
            I => \N__42770\
        );

    \I__8357\ : InMux
    port map (
            O => \N__42793\,
            I => \N__42755\
        );

    \I__8356\ : InMux
    port map (
            O => \N__42792\,
            I => \N__42755\
        );

    \I__8355\ : InMux
    port map (
            O => \N__42791\,
            I => \N__42755\
        );

    \I__8354\ : InMux
    port map (
            O => \N__42790\,
            I => \N__42755\
        );

    \I__8353\ : InMux
    port map (
            O => \N__42789\,
            I => \N__42755\
        );

    \I__8352\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42752\
        );

    \I__8351\ : InMux
    port map (
            O => \N__42787\,
            I => \N__42745\
        );

    \I__8350\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42745\
        );

    \I__8349\ : InMux
    port map (
            O => \N__42785\,
            I => \N__42745\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__42782\,
            I => \N__42740\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__42779\,
            I => \N__42737\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__42770\,
            I => \N__42734\
        );

    \I__8345\ : InMux
    port map (
            O => \N__42769\,
            I => \N__42729\
        );

    \I__8344\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42729\
        );

    \I__8343\ : InMux
    port map (
            O => \N__42767\,
            I => \N__42724\
        );

    \I__8342\ : InMux
    port map (
            O => \N__42766\,
            I => \N__42724\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__42755\,
            I => \N__42721\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__42752\,
            I => \N__42716\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__42745\,
            I => \N__42716\
        );

    \I__8338\ : InMux
    port map (
            O => \N__42744\,
            I => \N__42711\
        );

    \I__8337\ : InMux
    port map (
            O => \N__42743\,
            I => \N__42711\
        );

    \I__8336\ : Span4Mux_v
    port map (
            O => \N__42740\,
            I => \N__42700\
        );

    \I__8335\ : Span4Mux_h
    port map (
            O => \N__42737\,
            I => \N__42693\
        );

    \I__8334\ : Span4Mux_h
    port map (
            O => \N__42734\,
            I => \N__42693\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__42729\,
            I => \N__42693\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__42724\,
            I => \N__42690\
        );

    \I__8331\ : Span4Mux_h
    port map (
            O => \N__42721\,
            I => \N__42687\
        );

    \I__8330\ : Span4Mux_v
    port map (
            O => \N__42716\,
            I => \N__42682\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__42711\,
            I => \N__42682\
        );

    \I__8328\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42675\
        );

    \I__8327\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42675\
        );

    \I__8326\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42675\
        );

    \I__8325\ : InMux
    port map (
            O => \N__42707\,
            I => \N__42664\
        );

    \I__8324\ : InMux
    port map (
            O => \N__42706\,
            I => \N__42664\
        );

    \I__8323\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42664\
        );

    \I__8322\ : InMux
    port map (
            O => \N__42704\,
            I => \N__42664\
        );

    \I__8321\ : InMux
    port map (
            O => \N__42703\,
            I => \N__42664\
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__42700\,
            I => \c0.n9668\
        );

    \I__8319\ : Odrv4
    port map (
            O => \N__42693\,
            I => \c0.n9668\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__42690\,
            I => \c0.n9668\
        );

    \I__8317\ : Odrv4
    port map (
            O => \N__42687\,
            I => \c0.n9668\
        );

    \I__8316\ : Odrv4
    port map (
            O => \N__42682\,
            I => \c0.n9668\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__42675\,
            I => \c0.n9668\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__42664\,
            I => \c0.n9668\
        );

    \I__8313\ : InMux
    port map (
            O => \N__42649\,
            I => \N__42646\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__42646\,
            I => \c0.n7_adj_4356\
        );

    \I__8311\ : InMux
    port map (
            O => \N__42643\,
            I => \N__42640\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__42640\,
            I => \N__42635\
        );

    \I__8309\ : InMux
    port map (
            O => \N__42639\,
            I => \N__42632\
        );

    \I__8308\ : InMux
    port map (
            O => \N__42638\,
            I => \N__42629\
        );

    \I__8307\ : Span4Mux_v
    port map (
            O => \N__42635\,
            I => \N__42624\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__42632\,
            I => \N__42624\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__42629\,
            I => \N__42621\
        );

    \I__8304\ : Odrv4
    port map (
            O => \N__42624\,
            I => \c0.n12876\
        );

    \I__8303\ : Odrv4
    port map (
            O => \N__42621\,
            I => \c0.n12876\
        );

    \I__8302\ : CascadeMux
    port map (
            O => \N__42616\,
            I => \N__42612\
        );

    \I__8301\ : InMux
    port map (
            O => \N__42615\,
            I => \N__42605\
        );

    \I__8300\ : InMux
    port map (
            O => \N__42612\,
            I => \N__42605\
        );

    \I__8299\ : InMux
    port map (
            O => \N__42611\,
            I => \N__42602\
        );

    \I__8298\ : InMux
    port map (
            O => \N__42610\,
            I => \N__42599\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__42605\,
            I => \N__42594\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__42602\,
            I => \N__42594\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__42599\,
            I => \c0.n21022\
        );

    \I__8294\ : Odrv4
    port map (
            O => \N__42594\,
            I => \c0.n21022\
        );

    \I__8293\ : InMux
    port map (
            O => \N__42589\,
            I => \N__42586\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__42586\,
            I => \N__42581\
        );

    \I__8291\ : InMux
    port map (
            O => \N__42585\,
            I => \N__42578\
        );

    \I__8290\ : InMux
    port map (
            O => \N__42584\,
            I => \N__42575\
        );

    \I__8289\ : Odrv4
    port map (
            O => \N__42581\,
            I => \c0.n12991\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__42578\,
            I => \c0.n12991\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__42575\,
            I => \c0.n12991\
        );

    \I__8286\ : InMux
    port map (
            O => \N__42568\,
            I => \N__42564\
        );

    \I__8285\ : CascadeMux
    port map (
            O => \N__42567\,
            I => \N__42561\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__42564\,
            I => \N__42558\
        );

    \I__8283\ : InMux
    port map (
            O => \N__42561\,
            I => \N__42555\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__42558\,
            I => \c0.n5024\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__42555\,
            I => \c0.n5024\
        );

    \I__8280\ : CascadeMux
    port map (
            O => \N__42550\,
            I => \c0.n5_adj_4342_cascade_\
        );

    \I__8279\ : InMux
    port map (
            O => \N__42547\,
            I => \N__42542\
        );

    \I__8278\ : InMux
    port map (
            O => \N__42546\,
            I => \N__42539\
        );

    \I__8277\ : CascadeMux
    port map (
            O => \N__42545\,
            I => \N__42535\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__42542\,
            I => \N__42532\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__42539\,
            I => \N__42529\
        );

    \I__8274\ : InMux
    port map (
            O => \N__42538\,
            I => \N__42524\
        );

    \I__8273\ : InMux
    port map (
            O => \N__42535\,
            I => \N__42524\
        );

    \I__8272\ : Span4Mux_v
    port map (
            O => \N__42532\,
            I => \N__42521\
        );

    \I__8271\ : Span4Mux_v
    port map (
            O => \N__42529\,
            I => \N__42518\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__42524\,
            I => \N__42515\
        );

    \I__8269\ : Odrv4
    port map (
            O => \N__42521\,
            I => \c0.n21686\
        );

    \I__8268\ : Odrv4
    port map (
            O => \N__42518\,
            I => \c0.n21686\
        );

    \I__8267\ : Odrv4
    port map (
            O => \N__42515\,
            I => \c0.n21686\
        );

    \I__8266\ : CascadeMux
    port map (
            O => \N__42508\,
            I => \N__42503\
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__42507\,
            I => \N__42499\
        );

    \I__8264\ : InMux
    port map (
            O => \N__42506\,
            I => \N__42495\
        );

    \I__8263\ : InMux
    port map (
            O => \N__42503\,
            I => \N__42490\
        );

    \I__8262\ : InMux
    port map (
            O => \N__42502\,
            I => \N__42487\
        );

    \I__8261\ : InMux
    port map (
            O => \N__42499\,
            I => \N__42484\
        );

    \I__8260\ : InMux
    port map (
            O => \N__42498\,
            I => \N__42481\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__42495\,
            I => \N__42478\
        );

    \I__8258\ : InMux
    port map (
            O => \N__42494\,
            I => \N__42473\
        );

    \I__8257\ : InMux
    port map (
            O => \N__42493\,
            I => \N__42473\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__42490\,
            I => \N__42470\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__42487\,
            I => \N__42463\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__42484\,
            I => \N__42463\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__42481\,
            I => \N__42463\
        );

    \I__8252\ : Span4Mux_h
    port map (
            O => \N__42478\,
            I => \N__42460\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__42473\,
            I => \N__42453\
        );

    \I__8250\ : Span4Mux_v
    port map (
            O => \N__42470\,
            I => \N__42453\
        );

    \I__8249\ : Span4Mux_v
    port map (
            O => \N__42463\,
            I => \N__42453\
        );

    \I__8248\ : Odrv4
    port map (
            O => \N__42460\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__8247\ : Odrv4
    port map (
            O => \N__42453\,
            I => \c0.FRAME_MATCHER_state_3\
        );

    \I__8246\ : CascadeMux
    port map (
            O => \N__42448\,
            I => \c0.n21686_cascade_\
        );

    \I__8245\ : SRMux
    port map (
            O => \N__42445\,
            I => \N__42442\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__42442\,
            I => \N__42439\
        );

    \I__8243\ : Span4Mux_h
    port map (
            O => \N__42439\,
            I => \N__42436\
        );

    \I__8242\ : Odrv4
    port map (
            O => \N__42436\,
            I => \c0.n21334\
        );

    \I__8241\ : CascadeMux
    port map (
            O => \N__42433\,
            I => \N__42430\
        );

    \I__8240\ : InMux
    port map (
            O => \N__42430\,
            I => \N__42426\
        );

    \I__8239\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42423\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__42426\,
            I => \N__42420\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__42423\,
            I => \N__42417\
        );

    \I__8236\ : Span4Mux_h
    port map (
            O => \N__42420\,
            I => \N__42412\
        );

    \I__8235\ : Span4Mux_h
    port map (
            O => \N__42417\,
            I => \N__42412\
        );

    \I__8234\ : Odrv4
    port map (
            O => \N__42412\,
            I => \c0.n44_adj_4336\
        );

    \I__8233\ : InMux
    port map (
            O => \N__42409\,
            I => \N__42406\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__42406\,
            I => \c0.n1_adj_4349\
        );

    \I__8231\ : CascadeMux
    port map (
            O => \N__42403\,
            I => \N__42400\
        );

    \I__8230\ : InMux
    port map (
            O => \N__42400\,
            I => \N__42397\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__42397\,
            I => \N__42392\
        );

    \I__8228\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42389\
        );

    \I__8227\ : InMux
    port map (
            O => \N__42395\,
            I => \N__42386\
        );

    \I__8226\ : Span4Mux_v
    port map (
            O => \N__42392\,
            I => \N__42382\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__42389\,
            I => \N__42379\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__42386\,
            I => \N__42376\
        );

    \I__8223\ : InMux
    port map (
            O => \N__42385\,
            I => \N__42372\
        );

    \I__8222\ : Sp12to4
    port map (
            O => \N__42382\,
            I => \N__42367\
        );

    \I__8221\ : Span12Mux_v
    port map (
            O => \N__42379\,
            I => \N__42367\
        );

    \I__8220\ : Span4Mux_v
    port map (
            O => \N__42376\,
            I => \N__42364\
        );

    \I__8219\ : InMux
    port map (
            O => \N__42375\,
            I => \N__42361\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__42372\,
            I => control_mode_4
        );

    \I__8217\ : Odrv12
    port map (
            O => \N__42367\,
            I => control_mode_4
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__42364\,
            I => control_mode_4
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__42361\,
            I => control_mode_4
        );

    \I__8214\ : CascadeMux
    port map (
            O => \N__42352\,
            I => \N__42348\
        );

    \I__8213\ : InMux
    port map (
            O => \N__42351\,
            I => \N__42345\
        );

    \I__8212\ : InMux
    port map (
            O => \N__42348\,
            I => \N__42342\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__42345\,
            I => \N__42339\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__42342\,
            I => \N__42333\
        );

    \I__8209\ : Span4Mux_h
    port map (
            O => \N__42339\,
            I => \N__42330\
        );

    \I__8208\ : InMux
    port map (
            O => \N__42338\,
            I => \N__42325\
        );

    \I__8207\ : InMux
    port map (
            O => \N__42337\,
            I => \N__42325\
        );

    \I__8206\ : InMux
    port map (
            O => \N__42336\,
            I => \N__42322\
        );

    \I__8205\ : Span4Mux_h
    port map (
            O => \N__42333\,
            I => \N__42315\
        );

    \I__8204\ : Span4Mux_v
    port map (
            O => \N__42330\,
            I => \N__42315\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__42325\,
            I => \N__42315\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__42322\,
            I => control_mode_7
        );

    \I__8201\ : Odrv4
    port map (
            O => \N__42315\,
            I => control_mode_7
        );

    \I__8200\ : CascadeMux
    port map (
            O => \N__42310\,
            I => \n23726_cascade_\
        );

    \I__8199\ : InMux
    port map (
            O => \N__42307\,
            I => \N__42303\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__42306\,
            I => \N__42300\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__42303\,
            I => \N__42297\
        );

    \I__8196\ : InMux
    port map (
            O => \N__42300\,
            I => \N__42294\
        );

    \I__8195\ : Span4Mux_v
    port map (
            O => \N__42297\,
            I => \N__42290\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__42294\,
            I => \N__42287\
        );

    \I__8193\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42283\
        );

    \I__8192\ : Sp12to4
    port map (
            O => \N__42290\,
            I => \N__42280\
        );

    \I__8191\ : Span4Mux_h
    port map (
            O => \N__42287\,
            I => \N__42277\
        );

    \I__8190\ : InMux
    port map (
            O => \N__42286\,
            I => \N__42274\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__42283\,
            I => control_mode_6
        );

    \I__8188\ : Odrv12
    port map (
            O => \N__42280\,
            I => control_mode_6
        );

    \I__8187\ : Odrv4
    port map (
            O => \N__42277\,
            I => control_mode_6
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__42274\,
            I => control_mode_6
        );

    \I__8185\ : InMux
    port map (
            O => \N__42265\,
            I => \N__42262\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__42262\,
            I => \N__42259\
        );

    \I__8183\ : Span4Mux_h
    port map (
            O => \N__42259\,
            I => \N__42256\
        );

    \I__8182\ : Odrv4
    port map (
            O => \N__42256\,
            I => n2249
        );

    \I__8181\ : CascadeMux
    port map (
            O => \N__42253\,
            I => \N__42245\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__42252\,
            I => \N__42242\
        );

    \I__8179\ : InMux
    port map (
            O => \N__42251\,
            I => \N__42224\
        );

    \I__8178\ : InMux
    port map (
            O => \N__42250\,
            I => \N__42224\
        );

    \I__8177\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42224\
        );

    \I__8176\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42210\
        );

    \I__8175\ : InMux
    port map (
            O => \N__42245\,
            I => \N__42210\
        );

    \I__8174\ : InMux
    port map (
            O => \N__42242\,
            I => \N__42210\
        );

    \I__8173\ : InMux
    port map (
            O => \N__42241\,
            I => \N__42210\
        );

    \I__8172\ : InMux
    port map (
            O => \N__42240\,
            I => \N__42210\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__42239\,
            I => \N__42205\
        );

    \I__8170\ : InMux
    port map (
            O => \N__42238\,
            I => \N__42199\
        );

    \I__8169\ : InMux
    port map (
            O => \N__42237\,
            I => \N__42190\
        );

    \I__8168\ : InMux
    port map (
            O => \N__42236\,
            I => \N__42190\
        );

    \I__8167\ : InMux
    port map (
            O => \N__42235\,
            I => \N__42190\
        );

    \I__8166\ : InMux
    port map (
            O => \N__42234\,
            I => \N__42190\
        );

    \I__8165\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42187\
        );

    \I__8164\ : InMux
    port map (
            O => \N__42232\,
            I => \N__42184\
        );

    \I__8163\ : CascadeMux
    port map (
            O => \N__42231\,
            I => \N__42181\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__42224\,
            I => \N__42177\
        );

    \I__8161\ : InMux
    port map (
            O => \N__42223\,
            I => \N__42172\
        );

    \I__8160\ : InMux
    port map (
            O => \N__42222\,
            I => \N__42172\
        );

    \I__8159\ : CascadeMux
    port map (
            O => \N__42221\,
            I => \N__42169\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__42210\,
            I => \N__42164\
        );

    \I__8157\ : InMux
    port map (
            O => \N__42209\,
            I => \N__42155\
        );

    \I__8156\ : InMux
    port map (
            O => \N__42208\,
            I => \N__42155\
        );

    \I__8155\ : InMux
    port map (
            O => \N__42205\,
            I => \N__42155\
        );

    \I__8154\ : InMux
    port map (
            O => \N__42204\,
            I => \N__42155\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__42203\,
            I => \N__42152\
        );

    \I__8152\ : InMux
    port map (
            O => \N__42202\,
            I => \N__42147\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__42199\,
            I => \N__42138\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__42190\,
            I => \N__42138\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__42187\,
            I => \N__42138\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__42184\,
            I => \N__42138\
        );

    \I__8147\ : InMux
    port map (
            O => \N__42181\,
            I => \N__42133\
        );

    \I__8146\ : InMux
    port map (
            O => \N__42180\,
            I => \N__42133\
        );

    \I__8145\ : Span4Mux_h
    port map (
            O => \N__42177\,
            I => \N__42128\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__42172\,
            I => \N__42128\
        );

    \I__8143\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42123\
        );

    \I__8142\ : InMux
    port map (
            O => \N__42168\,
            I => \N__42123\
        );

    \I__8141\ : InMux
    port map (
            O => \N__42167\,
            I => \N__42120\
        );

    \I__8140\ : Span4Mux_v
    port map (
            O => \N__42164\,
            I => \N__42115\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__42155\,
            I => \N__42115\
        );

    \I__8138\ : InMux
    port map (
            O => \N__42152\,
            I => \N__42108\
        );

    \I__8137\ : InMux
    port map (
            O => \N__42151\,
            I => \N__42108\
        );

    \I__8136\ : InMux
    port map (
            O => \N__42150\,
            I => \N__42108\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__42147\,
            I => \N__42103\
        );

    \I__8134\ : Span4Mux_v
    port map (
            O => \N__42138\,
            I => \N__42100\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__42133\,
            I => \N__42097\
        );

    \I__8132\ : Span4Mux_h
    port map (
            O => \N__42128\,
            I => \N__42090\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__42123\,
            I => \N__42090\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__42120\,
            I => \N__42090\
        );

    \I__8129\ : Span4Mux_v
    port map (
            O => \N__42115\,
            I => \N__42085\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__42108\,
            I => \N__42085\
        );

    \I__8127\ : InMux
    port map (
            O => \N__42107\,
            I => \N__42082\
        );

    \I__8126\ : InMux
    port map (
            O => \N__42106\,
            I => \N__42079\
        );

    \I__8125\ : Span4Mux_v
    port map (
            O => \N__42103\,
            I => \N__42076\
        );

    \I__8124\ : Span4Mux_h
    port map (
            O => \N__42100\,
            I => \N__42071\
        );

    \I__8123\ : Span4Mux_v
    port map (
            O => \N__42097\,
            I => \N__42071\
        );

    \I__8122\ : Span4Mux_v
    port map (
            O => \N__42090\,
            I => \N__42062\
        );

    \I__8121\ : Span4Mux_h
    port map (
            O => \N__42085\,
            I => \N__42062\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__42082\,
            I => \N__42062\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__42079\,
            I => \N__42062\
        );

    \I__8118\ : Span4Mux_v
    port map (
            O => \N__42076\,
            I => \N__42059\
        );

    \I__8117\ : Span4Mux_v
    port map (
            O => \N__42071\,
            I => \N__42056\
        );

    \I__8116\ : Span4Mux_h
    port map (
            O => \N__42062\,
            I => \N__42053\
        );

    \I__8115\ : Odrv4
    port map (
            O => \N__42059\,
            I => count_enable
        );

    \I__8114\ : Odrv4
    port map (
            O => \N__42056\,
            I => count_enable
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__42053\,
            I => count_enable
        );

    \I__8112\ : InMux
    port map (
            O => \N__42046\,
            I => \N__42042\
        );

    \I__8111\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42038\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__42042\,
            I => \N__42035\
        );

    \I__8109\ : CascadeMux
    port map (
            O => \N__42041\,
            I => \N__42031\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__42038\,
            I => \N__42027\
        );

    \I__8107\ : Span4Mux_h
    port map (
            O => \N__42035\,
            I => \N__42024\
        );

    \I__8106\ : InMux
    port map (
            O => \N__42034\,
            I => \N__42021\
        );

    \I__8105\ : InMux
    port map (
            O => \N__42031\,
            I => \N__42018\
        );

    \I__8104\ : InMux
    port map (
            O => \N__42030\,
            I => \N__42015\
        );

    \I__8103\ : Span4Mux_h
    port map (
            O => \N__42027\,
            I => \N__42010\
        );

    \I__8102\ : Span4Mux_v
    port map (
            O => \N__42024\,
            I => \N__42010\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__42021\,
            I => \N__42007\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__42018\,
            I => encoder0_position_22
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__42015\,
            I => encoder0_position_22
        );

    \I__8098\ : Odrv4
    port map (
            O => \N__42010\,
            I => encoder0_position_22
        );

    \I__8097\ : Odrv4
    port map (
            O => \N__42007\,
            I => encoder0_position_22
        );

    \I__8096\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41995\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__41995\,
            I => \N__41989\
        );

    \I__8094\ : InMux
    port map (
            O => \N__41994\,
            I => \N__41986\
        );

    \I__8093\ : InMux
    port map (
            O => \N__41993\,
            I => \N__41981\
        );

    \I__8092\ : InMux
    port map (
            O => \N__41992\,
            I => \N__41981\
        );

    \I__8091\ : Span4Mux_v
    port map (
            O => \N__41989\,
            I => \N__41976\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__41986\,
            I => \N__41976\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__41981\,
            I => \N__41971\
        );

    \I__8088\ : Span4Mux_h
    port map (
            O => \N__41976\,
            I => \N__41971\
        );

    \I__8087\ : Odrv4
    port map (
            O => \N__41971\,
            I => data_in_2_4
        );

    \I__8086\ : InMux
    port map (
            O => \N__41968\,
            I => \N__41964\
        );

    \I__8085\ : InMux
    port map (
            O => \N__41967\,
            I => \N__41961\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__41964\,
            I => \N__41957\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__41961\,
            I => \N__41954\
        );

    \I__8082\ : CascadeMux
    port map (
            O => \N__41960\,
            I => \N__41951\
        );

    \I__8081\ : Span4Mux_v
    port map (
            O => \N__41957\,
            I => \N__41947\
        );

    \I__8080\ : Span4Mux_v
    port map (
            O => \N__41954\,
            I => \N__41944\
        );

    \I__8079\ : InMux
    port map (
            O => \N__41951\,
            I => \N__41941\
        );

    \I__8078\ : InMux
    port map (
            O => \N__41950\,
            I => \N__41938\
        );

    \I__8077\ : Span4Mux_h
    port map (
            O => \N__41947\,
            I => \N__41935\
        );

    \I__8076\ : Sp12to4
    port map (
            O => \N__41944\,
            I => \N__41930\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__41941\,
            I => \N__41930\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__41938\,
            I => data_in_1_4
        );

    \I__8073\ : Odrv4
    port map (
            O => \N__41935\,
            I => data_in_1_4
        );

    \I__8072\ : Odrv12
    port map (
            O => \N__41930\,
            I => data_in_1_4
        );

    \I__8071\ : InMux
    port map (
            O => \N__41923\,
            I => \N__41920\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__41920\,
            I => \N__41917\
        );

    \I__8069\ : Span4Mux_h
    port map (
            O => \N__41917\,
            I => \N__41914\
        );

    \I__8068\ : Span4Mux_h
    port map (
            O => \N__41914\,
            I => \N__41910\
        );

    \I__8067\ : InMux
    port map (
            O => \N__41913\,
            I => \N__41907\
        );

    \I__8066\ : Span4Mux_v
    port map (
            O => \N__41910\,
            I => \N__41904\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__41907\,
            I => \c0.FRAME_MATCHER_rx_data_ready_prev\
        );

    \I__8064\ : Odrv4
    port map (
            O => \N__41904\,
            I => \c0.FRAME_MATCHER_rx_data_ready_prev\
        );

    \I__8063\ : CascadeMux
    port map (
            O => \N__41899\,
            I => \c0.n17790_cascade_\
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__41896\,
            I => \c0.n21775_cascade_\
        );

    \I__8061\ : InMux
    port map (
            O => \N__41893\,
            I => \N__41890\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__41890\,
            I => \N__41885\
        );

    \I__8059\ : InMux
    port map (
            O => \N__41889\,
            I => \N__41880\
        );

    \I__8058\ : InMux
    port map (
            O => \N__41888\,
            I => \N__41880\
        );

    \I__8057\ : Span4Mux_h
    port map (
            O => \N__41885\,
            I => \N__41877\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__41880\,
            I => data_in_3_4
        );

    \I__8055\ : Odrv4
    port map (
            O => \N__41877\,
            I => data_in_3_4
        );

    \I__8054\ : InMux
    port map (
            O => \N__41872\,
            I => \N__41866\
        );

    \I__8053\ : InMux
    port map (
            O => \N__41871\,
            I => \N__41863\
        );

    \I__8052\ : InMux
    port map (
            O => \N__41870\,
            I => \N__41859\
        );

    \I__8051\ : InMux
    port map (
            O => \N__41869\,
            I => \N__41856\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__41866\,
            I => \N__41853\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__41863\,
            I => \N__41850\
        );

    \I__8048\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41847\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__41859\,
            I => \N__41844\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__41856\,
            I => \N__41840\
        );

    \I__8045\ : Span4Mux_v
    port map (
            O => \N__41853\,
            I => \N__41833\
        );

    \I__8044\ : Span4Mux_v
    port map (
            O => \N__41850\,
            I => \N__41833\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__41847\,
            I => \N__41833\
        );

    \I__8042\ : Span4Mux_h
    port map (
            O => \N__41844\,
            I => \N__41830\
        );

    \I__8041\ : InMux
    port map (
            O => \N__41843\,
            I => \N__41827\
        );

    \I__8040\ : Span4Mux_v
    port map (
            O => \N__41840\,
            I => \N__41822\
        );

    \I__8039\ : Span4Mux_h
    port map (
            O => \N__41833\,
            I => \N__41822\
        );

    \I__8038\ : Odrv4
    port map (
            O => \N__41830\,
            I => control_mode_1
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__41827\,
            I => control_mode_1
        );

    \I__8036\ : Odrv4
    port map (
            O => \N__41822\,
            I => control_mode_1
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__41815\,
            I => \N__41812\
        );

    \I__8034\ : InMux
    port map (
            O => \N__41812\,
            I => \N__41807\
        );

    \I__8033\ : InMux
    port map (
            O => \N__41811\,
            I => \N__41804\
        );

    \I__8032\ : InMux
    port map (
            O => \N__41810\,
            I => \N__41801\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__41807\,
            I => \N__41796\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__41804\,
            I => \N__41791\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__41801\,
            I => \N__41791\
        );

    \I__8028\ : InMux
    port map (
            O => \N__41800\,
            I => \N__41788\
        );

    \I__8027\ : InMux
    port map (
            O => \N__41799\,
            I => \N__41785\
        );

    \I__8026\ : Span4Mux_v
    port map (
            O => \N__41796\,
            I => \N__41781\
        );

    \I__8025\ : Span4Mux_v
    port map (
            O => \N__41791\,
            I => \N__41774\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__41788\,
            I => \N__41774\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__41785\,
            I => \N__41774\
        );

    \I__8022\ : InMux
    port map (
            O => \N__41784\,
            I => \N__41771\
        );

    \I__8021\ : Span4Mux_h
    port map (
            O => \N__41781\,
            I => \N__41768\
        );

    \I__8020\ : Span4Mux_h
    port map (
            O => \N__41774\,
            I => \N__41765\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__41771\,
            I => control_mode_3
        );

    \I__8018\ : Odrv4
    port map (
            O => \N__41768\,
            I => control_mode_3
        );

    \I__8017\ : Odrv4
    port map (
            O => \N__41765\,
            I => control_mode_3
        );

    \I__8016\ : CascadeMux
    port map (
            O => \N__41758\,
            I => \N__41755\
        );

    \I__8015\ : InMux
    port map (
            O => \N__41755\,
            I => \N__41751\
        );

    \I__8014\ : InMux
    port map (
            O => \N__41754\,
            I => \N__41747\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__41751\,
            I => \N__41741\
        );

    \I__8012\ : InMux
    port map (
            O => \N__41750\,
            I => \N__41738\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__41747\,
            I => \N__41735\
        );

    \I__8010\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41728\
        );

    \I__8009\ : InMux
    port map (
            O => \N__41745\,
            I => \N__41728\
        );

    \I__8008\ : InMux
    port map (
            O => \N__41744\,
            I => \N__41728\
        );

    \I__8007\ : Span4Mux_h
    port map (
            O => \N__41741\,
            I => \N__41723\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__41738\,
            I => \N__41723\
        );

    \I__8005\ : Span4Mux_h
    port map (
            O => \N__41735\,
            I => \N__41719\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__41728\,
            I => \N__41714\
        );

    \I__8003\ : Span4Mux_h
    port map (
            O => \N__41723\,
            I => \N__41714\
        );

    \I__8002\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41711\
        );

    \I__8001\ : Odrv4
    port map (
            O => \N__41719\,
            I => encoder0_position_18
        );

    \I__8000\ : Odrv4
    port map (
            O => \N__41714\,
            I => encoder0_position_18
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__41711\,
            I => encoder0_position_18
        );

    \I__7998\ : CascadeMux
    port map (
            O => \N__41704\,
            I => \N__41701\
        );

    \I__7997\ : InMux
    port map (
            O => \N__41701\,
            I => \N__41697\
        );

    \I__7996\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41693\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__41697\,
            I => \N__41690\
        );

    \I__7994\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41687\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__41693\,
            I => \N__41684\
        );

    \I__7992\ : Span4Mux_v
    port map (
            O => \N__41690\,
            I => \N__41679\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__41687\,
            I => \N__41674\
        );

    \I__7990\ : Span4Mux_v
    port map (
            O => \N__41684\,
            I => \N__41674\
        );

    \I__7989\ : CascadeMux
    port map (
            O => \N__41683\,
            I => \N__41670\
        );

    \I__7988\ : InMux
    port map (
            O => \N__41682\,
            I => \N__41667\
        );

    \I__7987\ : Span4Mux_h
    port map (
            O => \N__41679\,
            I => \N__41662\
        );

    \I__7986\ : Span4Mux_h
    port map (
            O => \N__41674\,
            I => \N__41662\
        );

    \I__7985\ : InMux
    port map (
            O => \N__41673\,
            I => \N__41657\
        );

    \I__7984\ : InMux
    port map (
            O => \N__41670\,
            I => \N__41657\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__41667\,
            I => encoder0_position_3
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__41662\,
            I => encoder0_position_3
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__41657\,
            I => encoder0_position_3
        );

    \I__7980\ : InMux
    port map (
            O => \N__41650\,
            I => \N__41642\
        );

    \I__7979\ : InMux
    port map (
            O => \N__41649\,
            I => \N__41635\
        );

    \I__7978\ : InMux
    port map (
            O => \N__41648\,
            I => \N__41635\
        );

    \I__7977\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41635\
        );

    \I__7976\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41632\
        );

    \I__7975\ : CascadeMux
    port map (
            O => \N__41645\,
            I => \N__41629\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__41642\,
            I => \N__41623\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__41635\,
            I => \N__41623\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__41632\,
            I => \N__41620\
        );

    \I__7971\ : InMux
    port map (
            O => \N__41629\,
            I => \N__41615\
        );

    \I__7970\ : InMux
    port map (
            O => \N__41628\,
            I => \N__41615\
        );

    \I__7969\ : Span4Mux_h
    port map (
            O => \N__41623\,
            I => \N__41612\
        );

    \I__7968\ : Odrv12
    port map (
            O => \N__41620\,
            I => encoder0_position_31
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__41615\,
            I => encoder0_position_31
        );

    \I__7966\ : Odrv4
    port map (
            O => \N__41612\,
            I => encoder0_position_31
        );

    \I__7965\ : CascadeMux
    port map (
            O => \N__41605\,
            I => \N__41602\
        );

    \I__7964\ : InMux
    port map (
            O => \N__41602\,
            I => \N__41598\
        );

    \I__7963\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41595\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__41598\,
            I => \N__41592\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__41595\,
            I => \N__41587\
        );

    \I__7960\ : Span4Mux_v
    port map (
            O => \N__41592\,
            I => \N__41587\
        );

    \I__7959\ : Span4Mux_h
    port map (
            O => \N__41587\,
            I => \N__41584\
        );

    \I__7958\ : Odrv4
    port map (
            O => \N__41584\,
            I => \c0.n21813\
        );

    \I__7957\ : CascadeMux
    port map (
            O => \N__41581\,
            I => \N__41578\
        );

    \I__7956\ : InMux
    port map (
            O => \N__41578\,
            I => \N__41574\
        );

    \I__7955\ : InMux
    port map (
            O => \N__41577\,
            I => \N__41571\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__41574\,
            I => \N__41568\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__41571\,
            I => data_in_frame_6_5
        );

    \I__7952\ : Odrv12
    port map (
            O => \N__41568\,
            I => data_in_frame_6_5
        );

    \I__7951\ : InMux
    port map (
            O => \N__41563\,
            I => \N__41560\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__41560\,
            I => \N__41557\
        );

    \I__7949\ : Span4Mux_h
    port map (
            O => \N__41557\,
            I => \N__41554\
        );

    \I__7948\ : Span4Mux_v
    port map (
            O => \N__41554\,
            I => \N__41551\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__41551\,
            I => \c0.tx.n23987\
        );

    \I__7946\ : InMux
    port map (
            O => \N__41548\,
            I => \N__41541\
        );

    \I__7945\ : InMux
    port map (
            O => \N__41547\,
            I => \N__41541\
        );

    \I__7944\ : InMux
    port map (
            O => \N__41546\,
            I => \N__41538\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__41541\,
            I => \N__41535\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__41538\,
            I => \N__41531\
        );

    \I__7941\ : Span4Mux_h
    port map (
            O => \N__41535\,
            I => \N__41528\
        );

    \I__7940\ : InMux
    port map (
            O => \N__41534\,
            I => \N__41525\
        );

    \I__7939\ : Span12Mux_h
    port map (
            O => \N__41531\,
            I => \N__41522\
        );

    \I__7938\ : Span4Mux_v
    port map (
            O => \N__41528\,
            I => \N__41519\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__41525\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__7936\ : Odrv12
    port map (
            O => \N__41522\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__7935\ : Odrv4
    port map (
            O => \N__41519\,
            I => \c0.tx.r_Clock_Count_6\
        );

    \I__7934\ : InMux
    port map (
            O => \N__41512\,
            I => \N__41509\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__41509\,
            I => \N__41506\
        );

    \I__7932\ : Span4Mux_v
    port map (
            O => \N__41506\,
            I => \N__41503\
        );

    \I__7931\ : Span4Mux_h
    port map (
            O => \N__41503\,
            I => \N__41500\
        );

    \I__7930\ : Odrv4
    port map (
            O => \N__41500\,
            I => n313
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__41497\,
            I => \N__41493\
        );

    \I__7928\ : CascadeMux
    port map (
            O => \N__41496\,
            I => \N__41487\
        );

    \I__7927\ : InMux
    port map (
            O => \N__41493\,
            I => \N__41479\
        );

    \I__7926\ : InMux
    port map (
            O => \N__41492\,
            I => \N__41479\
        );

    \I__7925\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41476\
        );

    \I__7924\ : InMux
    port map (
            O => \N__41490\,
            I => \N__41471\
        );

    \I__7923\ : InMux
    port map (
            O => \N__41487\,
            I => \N__41471\
        );

    \I__7922\ : InMux
    port map (
            O => \N__41486\,
            I => \N__41468\
        );

    \I__7921\ : InMux
    port map (
            O => \N__41485\,
            I => \N__41462\
        );

    \I__7920\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41462\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__41479\,
            I => \N__41459\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__41476\,
            I => \N__41451\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__41471\,
            I => \N__41446\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__41468\,
            I => \N__41446\
        );

    \I__7915\ : CascadeMux
    port map (
            O => \N__41467\,
            I => \N__41440\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__41462\,
            I => \N__41437\
        );

    \I__7913\ : Span4Mux_h
    port map (
            O => \N__41459\,
            I => \N__41434\
        );

    \I__7912\ : InMux
    port map (
            O => \N__41458\,
            I => \N__41429\
        );

    \I__7911\ : InMux
    port map (
            O => \N__41457\,
            I => \N__41429\
        );

    \I__7910\ : InMux
    port map (
            O => \N__41456\,
            I => \N__41422\
        );

    \I__7909\ : InMux
    port map (
            O => \N__41455\,
            I => \N__41422\
        );

    \I__7908\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41422\
        );

    \I__7907\ : Span4Mux_h
    port map (
            O => \N__41451\,
            I => \N__41419\
        );

    \I__7906\ : Span4Mux_v
    port map (
            O => \N__41446\,
            I => \N__41416\
        );

    \I__7905\ : InMux
    port map (
            O => \N__41445\,
            I => \N__41413\
        );

    \I__7904\ : InMux
    port map (
            O => \N__41444\,
            I => \N__41406\
        );

    \I__7903\ : InMux
    port map (
            O => \N__41443\,
            I => \N__41406\
        );

    \I__7902\ : InMux
    port map (
            O => \N__41440\,
            I => \N__41406\
        );

    \I__7901\ : Span4Mux_v
    port map (
            O => \N__41437\,
            I => \N__41399\
        );

    \I__7900\ : Span4Mux_v
    port map (
            O => \N__41434\,
            I => \N__41399\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__41429\,
            I => \N__41399\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__41422\,
            I => \r_SM_Main_2_adj_4549\
        );

    \I__7897\ : Odrv4
    port map (
            O => \N__41419\,
            I => \r_SM_Main_2_adj_4549\
        );

    \I__7896\ : Odrv4
    port map (
            O => \N__41416\,
            I => \r_SM_Main_2_adj_4549\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__41413\,
            I => \r_SM_Main_2_adj_4549\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__41406\,
            I => \r_SM_Main_2_adj_4549\
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__41399\,
            I => \r_SM_Main_2_adj_4549\
        );

    \I__7892\ : InMux
    port map (
            O => \N__41386\,
            I => \N__41383\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__41383\,
            I => \N__41379\
        );

    \I__7890\ : InMux
    port map (
            O => \N__41382\,
            I => \N__41370\
        );

    \I__7889\ : Span4Mux_h
    port map (
            O => \N__41379\,
            I => \N__41367\
        );

    \I__7888\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41362\
        );

    \I__7887\ : InMux
    port map (
            O => \N__41377\,
            I => \N__41362\
        );

    \I__7886\ : InMux
    port map (
            O => \N__41376\,
            I => \N__41353\
        );

    \I__7885\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41353\
        );

    \I__7884\ : InMux
    port map (
            O => \N__41374\,
            I => \N__41353\
        );

    \I__7883\ : InMux
    port map (
            O => \N__41373\,
            I => \N__41353\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__41370\,
            I => n8
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__41367\,
            I => n8
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__41362\,
            I => n8
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__41353\,
            I => n8
        );

    \I__7878\ : InMux
    port map (
            O => \N__41344\,
            I => \N__41339\
        );

    \I__7877\ : InMux
    port map (
            O => \N__41343\,
            I => \N__41334\
        );

    \I__7876\ : InMux
    port map (
            O => \N__41342\,
            I => \N__41334\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__41339\,
            I => \N__41331\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__41334\,
            I => \N__41328\
        );

    \I__7873\ : Span4Mux_v
    port map (
            O => \N__41331\,
            I => \N__41324\
        );

    \I__7872\ : Span4Mux_h
    port map (
            O => \N__41328\,
            I => \N__41321\
        );

    \I__7871\ : InMux
    port map (
            O => \N__41327\,
            I => \N__41318\
        );

    \I__7870\ : Span4Mux_h
    port map (
            O => \N__41324\,
            I => \N__41315\
        );

    \I__7869\ : Span4Mux_v
    port map (
            O => \N__41321\,
            I => \N__41312\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__41318\,
            I => \r_Clock_Count_8\
        );

    \I__7867\ : Odrv4
    port map (
            O => \N__41315\,
            I => \r_Clock_Count_8\
        );

    \I__7866\ : Odrv4
    port map (
            O => \N__41312\,
            I => \r_Clock_Count_8\
        );

    \I__7865\ : InMux
    port map (
            O => \N__41305\,
            I => \N__41302\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__41302\,
            I => \N__41299\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__41299\,
            I => \N__41296\
        );

    \I__7862\ : Odrv4
    port map (
            O => \N__41296\,
            I => n2253
        );

    \I__7861\ : InMux
    port map (
            O => \N__41293\,
            I => \N__41290\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__41290\,
            I => \N__41287\
        );

    \I__7859\ : Span12Mux_h
    port map (
            O => \N__41287\,
            I => \N__41284\
        );

    \I__7858\ : Odrv12
    port map (
            O => \N__41284\,
            I => \c0.n21816\
        );

    \I__7857\ : CascadeMux
    port map (
            O => \N__41281\,
            I => \c0.n21740_cascade_\
        );

    \I__7856\ : InMux
    port map (
            O => \N__41278\,
            I => \N__41274\
        );

    \I__7855\ : CascadeMux
    port map (
            O => \N__41277\,
            I => \N__41271\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__41274\,
            I => \N__41268\
        );

    \I__7853\ : InMux
    port map (
            O => \N__41271\,
            I => \N__41265\
        );

    \I__7852\ : Span4Mux_v
    port map (
            O => \N__41268\,
            I => \N__41262\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__41265\,
            I => \c0.data_in_frame_20_6\
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__41262\,
            I => \c0.data_in_frame_20_6\
        );

    \I__7849\ : CascadeMux
    port map (
            O => \N__41257\,
            I => \n21744_cascade_\
        );

    \I__7848\ : InMux
    port map (
            O => \N__41254\,
            I => \N__41250\
        );

    \I__7847\ : InMux
    port map (
            O => \N__41253\,
            I => \N__41247\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__41250\,
            I => \N__41244\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__41247\,
            I => data_in_frame_6_3
        );

    \I__7844\ : Odrv12
    port map (
            O => \N__41244\,
            I => data_in_frame_6_3
        );

    \I__7843\ : InMux
    port map (
            O => \N__41239\,
            I => \N__41236\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__41236\,
            I => \N__41233\
        );

    \I__7841\ : Span4Mux_h
    port map (
            O => \N__41233\,
            I => \N__41230\
        );

    \I__7840\ : Odrv4
    port map (
            O => \N__41230\,
            I => \c0.n25_adj_4408\
        );

    \I__7839\ : CascadeMux
    port map (
            O => \N__41227\,
            I => \N__41224\
        );

    \I__7838\ : InMux
    port map (
            O => \N__41224\,
            I => \N__41221\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__41221\,
            I => \N__41218\
        );

    \I__7836\ : Odrv4
    port map (
            O => \N__41218\,
            I => \c0.n23648\
        );

    \I__7835\ : InMux
    port map (
            O => \N__41215\,
            I => \N__41212\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__41212\,
            I => \c0.n16_adj_4401\
        );

    \I__7833\ : InMux
    port map (
            O => \N__41209\,
            I => \N__41205\
        );

    \I__7832\ : InMux
    port map (
            O => \N__41208\,
            I => \N__41202\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__41205\,
            I => \c0.n21893\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__41202\,
            I => \c0.n21893\
        );

    \I__7829\ : InMux
    port map (
            O => \N__41197\,
            I => \N__41194\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__41194\,
            I => \N__41191\
        );

    \I__7827\ : Odrv12
    port map (
            O => \N__41191\,
            I => \c0.n44_adj_4409\
        );

    \I__7826\ : CascadeMux
    port map (
            O => \N__41188\,
            I => \c0.n6_adj_4393_cascade_\
        );

    \I__7825\ : CascadeMux
    port map (
            O => \N__41185\,
            I => \c0.n13086_cascade_\
        );

    \I__7824\ : CascadeMux
    port map (
            O => \N__41182\,
            I => \c0.n21986_cascade_\
        );

    \I__7823\ : InMux
    port map (
            O => \N__41179\,
            I => \N__41173\
        );

    \I__7822\ : InMux
    port map (
            O => \N__41178\,
            I => \N__41173\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__41173\,
            I => data_in_frame_6_0
        );

    \I__7820\ : CascadeMux
    port map (
            O => \N__41170\,
            I => \c0.n38_adj_4407_cascade_\
        );

    \I__7819\ : InMux
    port map (
            O => \N__41167\,
            I => \N__41164\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__41164\,
            I => \c0.n23836\
        );

    \I__7817\ : CascadeMux
    port map (
            O => \N__41161\,
            I => \c0.n43_adj_4410_cascade_\
        );

    \I__7816\ : CascadeMux
    port map (
            O => \N__41158\,
            I => \c0.n22443_cascade_\
        );

    \I__7815\ : CascadeMux
    port map (
            O => \N__41155\,
            I => \N__41152\
        );

    \I__7814\ : InMux
    port map (
            O => \N__41152\,
            I => \N__41148\
        );

    \I__7813\ : InMux
    port map (
            O => \N__41151\,
            I => \N__41143\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__41148\,
            I => \N__41140\
        );

    \I__7811\ : InMux
    port map (
            O => \N__41147\,
            I => \N__41135\
        );

    \I__7810\ : InMux
    port map (
            O => \N__41146\,
            I => \N__41135\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__41143\,
            I => \N__41132\
        );

    \I__7808\ : Span4Mux_h
    port map (
            O => \N__41140\,
            I => \N__41129\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__41135\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__7806\ : Odrv4
    port map (
            O => \N__41132\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__7805\ : Odrv4
    port map (
            O => \N__41129\,
            I => \c0.FRAME_MATCHER_state_30\
        );

    \I__7804\ : SRMux
    port map (
            O => \N__41122\,
            I => \N__41119\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__41119\,
            I => \N__41116\
        );

    \I__7802\ : Span4Mux_h
    port map (
            O => \N__41116\,
            I => \N__41113\
        );

    \I__7801\ : Span4Mux_h
    port map (
            O => \N__41113\,
            I => \N__41110\
        );

    \I__7800\ : Odrv4
    port map (
            O => \N__41110\,
            I => \c0.n8_adj_4396\
        );

    \I__7799\ : CascadeMux
    port map (
            O => \N__41107\,
            I => \c0.n21737_cascade_\
        );

    \I__7798\ : CascadeMux
    port map (
            O => \N__41104\,
            I => \N__41101\
        );

    \I__7797\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41096\
        );

    \I__7796\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41093\
        );

    \I__7795\ : InMux
    port map (
            O => \N__41099\,
            I => \N__41090\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__41096\,
            I => \N__41087\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__41093\,
            I => \N__41084\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__41090\,
            I => \N__41076\
        );

    \I__7791\ : Sp12to4
    port map (
            O => \N__41087\,
            I => \N__41076\
        );

    \I__7790\ : Sp12to4
    port map (
            O => \N__41084\,
            I => \N__41076\
        );

    \I__7789\ : InMux
    port map (
            O => \N__41083\,
            I => \N__41073\
        );

    \I__7788\ : Span12Mux_v
    port map (
            O => \N__41076\,
            I => \N__41070\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__41073\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__7786\ : Odrv12
    port map (
            O => \N__41070\,
            I => \c0.FRAME_MATCHER_state_6\
        );

    \I__7785\ : SRMux
    port map (
            O => \N__41065\,
            I => \N__41062\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__41062\,
            I => \N__41059\
        );

    \I__7783\ : Span12Mux_v
    port map (
            O => \N__41059\,
            I => \N__41056\
        );

    \I__7782\ : Odrv12
    port map (
            O => \N__41056\,
            I => \c0.n21340\
        );

    \I__7781\ : InMux
    port map (
            O => \N__41053\,
            I => \N__41049\
        );

    \I__7780\ : CascadeMux
    port map (
            O => \N__41052\,
            I => \N__41045\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__41049\,
            I => \N__41042\
        );

    \I__7778\ : InMux
    port map (
            O => \N__41048\,
            I => \N__41038\
        );

    \I__7777\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41035\
        );

    \I__7776\ : Span4Mux_v
    port map (
            O => \N__41042\,
            I => \N__41032\
        );

    \I__7775\ : InMux
    port map (
            O => \N__41041\,
            I => \N__41029\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__41038\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__41035\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__7772\ : Odrv4
    port map (
            O => \N__41032\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__41029\,
            I => \c0.FRAME_MATCHER_state_19\
        );

    \I__7770\ : SRMux
    port map (
            O => \N__41020\,
            I => \N__41017\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__41017\,
            I => \N__41014\
        );

    \I__7768\ : Odrv12
    port map (
            O => \N__41014\,
            I => \c0.n8_adj_4398\
        );

    \I__7767\ : CascadeMux
    port map (
            O => \N__41011\,
            I => \N__41008\
        );

    \I__7766\ : InMux
    port map (
            O => \N__41008\,
            I => \N__41004\
        );

    \I__7765\ : InMux
    port map (
            O => \N__41007\,
            I => \N__41000\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__41004\,
            I => \N__40997\
        );

    \I__7763\ : InMux
    port map (
            O => \N__41003\,
            I => \N__40993\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__41000\,
            I => \N__40990\
        );

    \I__7761\ : Span4Mux_v
    port map (
            O => \N__40997\,
            I => \N__40987\
        );

    \I__7760\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40984\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__40993\,
            I => \N__40981\
        );

    \I__7758\ : Span4Mux_h
    port map (
            O => \N__40990\,
            I => \N__40978\
        );

    \I__7757\ : Span4Mux_h
    port map (
            O => \N__40987\,
            I => \N__40975\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__40984\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__7755\ : Odrv12
    port map (
            O => \N__40981\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__7754\ : Odrv4
    port map (
            O => \N__40978\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__7753\ : Odrv4
    port map (
            O => \N__40975\,
            I => \c0.FRAME_MATCHER_state_5\
        );

    \I__7752\ : SRMux
    port map (
            O => \N__40966\,
            I => \N__40963\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__40963\,
            I => \N__40960\
        );

    \I__7750\ : Span4Mux_h
    port map (
            O => \N__40960\,
            I => \N__40957\
        );

    \I__7749\ : Odrv4
    port map (
            O => \N__40957\,
            I => \c0.n21338\
        );

    \I__7748\ : CEMux
    port map (
            O => \N__40954\,
            I => \N__40947\
        );

    \I__7747\ : CEMux
    port map (
            O => \N__40953\,
            I => \N__40941\
        );

    \I__7746\ : CEMux
    port map (
            O => \N__40952\,
            I => \N__40938\
        );

    \I__7745\ : CEMux
    port map (
            O => \N__40951\,
            I => \N__40935\
        );

    \I__7744\ : CEMux
    port map (
            O => \N__40950\,
            I => \N__40931\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__40947\,
            I => \N__40928\
        );

    \I__7742\ : CEMux
    port map (
            O => \N__40946\,
            I => \N__40924\
        );

    \I__7741\ : CEMux
    port map (
            O => \N__40945\,
            I => \N__40921\
        );

    \I__7740\ : CEMux
    port map (
            O => \N__40944\,
            I => \N__40918\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__40941\,
            I => \N__40915\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__40938\,
            I => \N__40912\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__40935\,
            I => \N__40909\
        );

    \I__7736\ : SRMux
    port map (
            O => \N__40934\,
            I => \N__40906\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__40931\,
            I => \N__40903\
        );

    \I__7734\ : Span4Mux_v
    port map (
            O => \N__40928\,
            I => \N__40900\
        );

    \I__7733\ : SRMux
    port map (
            O => \N__40927\,
            I => \N__40897\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__40924\,
            I => \N__40894\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__40921\,
            I => \N__40891\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__40918\,
            I => \N__40886\
        );

    \I__7729\ : Span4Mux_v
    port map (
            O => \N__40915\,
            I => \N__40886\
        );

    \I__7728\ : Span4Mux_h
    port map (
            O => \N__40912\,
            I => \N__40883\
        );

    \I__7727\ : Span4Mux_v
    port map (
            O => \N__40909\,
            I => \N__40880\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__40906\,
            I => \N__40877\
        );

    \I__7725\ : Span4Mux_h
    port map (
            O => \N__40903\,
            I => \N__40874\
        );

    \I__7724\ : Span4Mux_v
    port map (
            O => \N__40900\,
            I => \N__40871\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__40897\,
            I => \N__40868\
        );

    \I__7722\ : Span4Mux_h
    port map (
            O => \N__40894\,
            I => \N__40865\
        );

    \I__7721\ : Span4Mux_v
    port map (
            O => \N__40891\,
            I => \N__40858\
        );

    \I__7720\ : Span4Mux_h
    port map (
            O => \N__40886\,
            I => \N__40858\
        );

    \I__7719\ : Span4Mux_v
    port map (
            O => \N__40883\,
            I => \N__40858\
        );

    \I__7718\ : Span4Mux_v
    port map (
            O => \N__40880\,
            I => \N__40855\
        );

    \I__7717\ : Span4Mux_h
    port map (
            O => \N__40877\,
            I => \N__40852\
        );

    \I__7716\ : Span4Mux_v
    port map (
            O => \N__40874\,
            I => \N__40849\
        );

    \I__7715\ : Span4Mux_h
    port map (
            O => \N__40871\,
            I => \N__40846\
        );

    \I__7714\ : Span4Mux_h
    port map (
            O => \N__40868\,
            I => \N__40843\
        );

    \I__7713\ : Sp12to4
    port map (
            O => \N__40865\,
            I => \N__40840\
        );

    \I__7712\ : Span4Mux_v
    port map (
            O => \N__40858\,
            I => \N__40837\
        );

    \I__7711\ : Span4Mux_h
    port map (
            O => \N__40855\,
            I => \N__40834\
        );

    \I__7710\ : Span4Mux_h
    port map (
            O => \N__40852\,
            I => \N__40829\
        );

    \I__7709\ : Span4Mux_v
    port map (
            O => \N__40849\,
            I => \N__40829\
        );

    \I__7708\ : Span4Mux_v
    port map (
            O => \N__40846\,
            I => \N__40826\
        );

    \I__7707\ : Sp12to4
    port map (
            O => \N__40843\,
            I => \N__40821\
        );

    \I__7706\ : Span12Mux_v
    port map (
            O => \N__40840\,
            I => \N__40821\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__40837\,
            I => \N__40818\
        );

    \I__7704\ : Odrv4
    port map (
            O => \N__40834\,
            I => \c0.n8107\
        );

    \I__7703\ : Odrv4
    port map (
            O => \N__40829\,
            I => \c0.n8107\
        );

    \I__7702\ : Odrv4
    port map (
            O => \N__40826\,
            I => \c0.n8107\
        );

    \I__7701\ : Odrv12
    port map (
            O => \N__40821\,
            I => \c0.n8107\
        );

    \I__7700\ : Odrv4
    port map (
            O => \N__40818\,
            I => \c0.n8107\
        );

    \I__7699\ : InMux
    port map (
            O => \N__40807\,
            I => \N__40804\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__40804\,
            I => \N__40801\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__40801\,
            I => \c0.n49\
        );

    \I__7696\ : CascadeMux
    port map (
            O => \N__40798\,
            I => \N__40795\
        );

    \I__7695\ : InMux
    port map (
            O => \N__40795\,
            I => \N__40792\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__40792\,
            I => \N__40789\
        );

    \I__7693\ : Span4Mux_v
    port map (
            O => \N__40789\,
            I => \N__40786\
        );

    \I__7692\ : Odrv4
    port map (
            O => \N__40786\,
            I => \c0.n50\
        );

    \I__7691\ : InMux
    port map (
            O => \N__40783\,
            I => \N__40780\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__40780\,
            I => \c0.n54\
        );

    \I__7689\ : SRMux
    port map (
            O => \N__40777\,
            I => \N__40770\
        );

    \I__7688\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40770\
        );

    \I__7687\ : InMux
    port map (
            O => \N__40775\,
            I => \N__40767\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__40770\,
            I => \N__40764\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__40767\,
            I => \N__40761\
        );

    \I__7684\ : Span12Mux_v
    port map (
            O => \N__40764\,
            I => \N__40758\
        );

    \I__7683\ : Span4Mux_v
    port map (
            O => \N__40761\,
            I => \N__40755\
        );

    \I__7682\ : Odrv12
    port map (
            O => \N__40758\,
            I => \c0.n22665\
        );

    \I__7681\ : Odrv4
    port map (
            O => \N__40755\,
            I => \c0.n22665\
        );

    \I__7680\ : CascadeMux
    port map (
            O => \N__40750\,
            I => \N__40746\
        );

    \I__7679\ : InMux
    port map (
            O => \N__40749\,
            I => \N__40741\
        );

    \I__7678\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40738\
        );

    \I__7677\ : InMux
    port map (
            O => \N__40745\,
            I => \N__40735\
        );

    \I__7676\ : CascadeMux
    port map (
            O => \N__40744\,
            I => \N__40731\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__40741\,
            I => \N__40728\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__40738\,
            I => \N__40725\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__40735\,
            I => \N__40722\
        );

    \I__7672\ : InMux
    port map (
            O => \N__40734\,
            I => \N__40717\
        );

    \I__7671\ : InMux
    port map (
            O => \N__40731\,
            I => \N__40717\
        );

    \I__7670\ : Span4Mux_v
    port map (
            O => \N__40728\,
            I => \N__40714\
        );

    \I__7669\ : Odrv4
    port map (
            O => \N__40725\,
            I => \c0.n3239\
        );

    \I__7668\ : Odrv4
    port map (
            O => \N__40722\,
            I => \c0.n3239\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__40717\,
            I => \c0.n3239\
        );

    \I__7666\ : Odrv4
    port map (
            O => \N__40714\,
            I => \c0.n3239\
        );

    \I__7665\ : CascadeMux
    port map (
            O => \N__40705\,
            I => \c0.n63_adj_4293_cascade_\
        );

    \I__7664\ : InMux
    port map (
            O => \N__40702\,
            I => \N__40698\
        );

    \I__7663\ : InMux
    port map (
            O => \N__40701\,
            I => \N__40695\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__40698\,
            I => \N__40690\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__40695\,
            I => \N__40690\
        );

    \I__7660\ : Odrv4
    port map (
            O => \N__40690\,
            I => \c0.n13020\
        );

    \I__7659\ : InMux
    port map (
            O => \N__40687\,
            I => \N__40684\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__40684\,
            I => \N__40681\
        );

    \I__7657\ : Span4Mux_h
    port map (
            O => \N__40681\,
            I => \N__40678\
        );

    \I__7656\ : Odrv4
    port map (
            O => \N__40678\,
            I => \c0.n4_adj_4345\
        );

    \I__7655\ : CascadeMux
    port map (
            O => \N__40675\,
            I => \c0.n84_cascade_\
        );

    \I__7654\ : InMux
    port map (
            O => \N__40672\,
            I => \N__40667\
        );

    \I__7653\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40662\
        );

    \I__7652\ : InMux
    port map (
            O => \N__40670\,
            I => \N__40662\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__40667\,
            I => \c0.n12990\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__40662\,
            I => \c0.n12990\
        );

    \I__7649\ : InMux
    port map (
            O => \N__40657\,
            I => \N__40654\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__40654\,
            I => \N__40649\
        );

    \I__7647\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40644\
        );

    \I__7646\ : InMux
    port map (
            O => \N__40652\,
            I => \N__40644\
        );

    \I__7645\ : Span12Mux_v
    port map (
            O => \N__40649\,
            I => \N__40641\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__40644\,
            I => \N__40638\
        );

    \I__7643\ : Odrv12
    port map (
            O => \N__40641\,
            I => \c0.n7_adj_4344\
        );

    \I__7642\ : Odrv4
    port map (
            O => \N__40638\,
            I => \c0.n7_adj_4344\
        );

    \I__7641\ : InMux
    port map (
            O => \N__40633\,
            I => \N__40630\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__40630\,
            I => \N__40625\
        );

    \I__7639\ : InMux
    port map (
            O => \N__40629\,
            I => \N__40618\
        );

    \I__7638\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40618\
        );

    \I__7637\ : Span4Mux_v
    port map (
            O => \N__40625\,
            I => \N__40615\
        );

    \I__7636\ : InMux
    port map (
            O => \N__40624\,
            I => \N__40610\
        );

    \I__7635\ : InMux
    port map (
            O => \N__40623\,
            I => \N__40610\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__40618\,
            I => \N__40607\
        );

    \I__7633\ : Odrv4
    port map (
            O => \N__40615\,
            I => \c0.n12967\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__40610\,
            I => \c0.n12967\
        );

    \I__7631\ : Odrv4
    port map (
            O => \N__40607\,
            I => \c0.n12967\
        );

    \I__7630\ : InMux
    port map (
            O => \N__40600\,
            I => \N__40592\
        );

    \I__7629\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40589\
        );

    \I__7628\ : CascadeMux
    port map (
            O => \N__40598\,
            I => \N__40586\
        );

    \I__7627\ : CascadeMux
    port map (
            O => \N__40597\,
            I => \N__40582\
        );

    \I__7626\ : InMux
    port map (
            O => \N__40596\,
            I => \N__40577\
        );

    \I__7625\ : InMux
    port map (
            O => \N__40595\,
            I => \N__40577\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__40592\,
            I => \N__40572\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__40589\,
            I => \N__40569\
        );

    \I__7622\ : InMux
    port map (
            O => \N__40586\,
            I => \N__40562\
        );

    \I__7621\ : InMux
    port map (
            O => \N__40585\,
            I => \N__40562\
        );

    \I__7620\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40562\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__40577\,
            I => \N__40559\
        );

    \I__7618\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40556\
        );

    \I__7617\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40553\
        );

    \I__7616\ : Odrv12
    port map (
            O => \N__40572\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7615\ : Odrv4
    port map (
            O => \N__40569\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__40562\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7613\ : Odrv4
    port map (
            O => \N__40559\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__40556\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__40553\,
            I => \c0.FRAME_MATCHER_state_0\
        );

    \I__7610\ : CascadeMux
    port map (
            O => \N__40540\,
            I => \N__40536\
        );

    \I__7609\ : InMux
    port map (
            O => \N__40539\,
            I => \N__40528\
        );

    \I__7608\ : InMux
    port map (
            O => \N__40536\,
            I => \N__40528\
        );

    \I__7607\ : InMux
    port map (
            O => \N__40535\,
            I => \N__40528\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__40528\,
            I => \N__40524\
        );

    \I__7605\ : InMux
    port map (
            O => \N__40527\,
            I => \N__40521\
        );

    \I__7604\ : Span4Mux_h
    port map (
            O => \N__40524\,
            I => \N__40516\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__40521\,
            I => \N__40516\
        );

    \I__7602\ : Odrv4
    port map (
            O => \N__40516\,
            I => \c0.n12996\
        );

    \I__7601\ : InMux
    port map (
            O => \N__40513\,
            I => \N__40509\
        );

    \I__7600\ : CascadeMux
    port map (
            O => \N__40512\,
            I => \N__40506\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__40509\,
            I => \N__40502\
        );

    \I__7598\ : InMux
    port map (
            O => \N__40506\,
            I => \N__40497\
        );

    \I__7597\ : InMux
    port map (
            O => \N__40505\,
            I => \N__40497\
        );

    \I__7596\ : Odrv4
    port map (
            O => \N__40502\,
            I => \c0.n4_adj_4419\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__40497\,
            I => \c0.n4_adj_4419\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__40492\,
            I => \c0.data_out_frame_0__7__N_2568_cascade_\
        );

    \I__7593\ : CascadeMux
    port map (
            O => \N__40489\,
            I => \c0.n1220_cascade_\
        );

    \I__7592\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40483\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__40483\,
            I => \N__40480\
        );

    \I__7590\ : Span12Mux_v
    port map (
            O => \N__40480\,
            I => \N__40477\
        );

    \I__7589\ : Odrv12
    port map (
            O => \N__40477\,
            I => \c0.n4_adj_4373\
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__40474\,
            I => \c0.n5024_cascade_\
        );

    \I__7587\ : InMux
    port map (
            O => \N__40471\,
            I => \N__40468\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__40468\,
            I => \N__40465\
        );

    \I__7585\ : Span4Mux_h
    port map (
            O => \N__40465\,
            I => \N__40462\
        );

    \I__7584\ : Odrv4
    port map (
            O => \N__40462\,
            I => \c0.n21773\
        );

    \I__7583\ : CascadeMux
    port map (
            O => \N__40459\,
            I => \c0.n21773_cascade_\
        );

    \I__7582\ : InMux
    port map (
            O => \N__40456\,
            I => \N__40448\
        );

    \I__7581\ : InMux
    port map (
            O => \N__40455\,
            I => \N__40448\
        );

    \I__7580\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40440\
        );

    \I__7579\ : InMux
    port map (
            O => \N__40453\,
            I => \N__40440\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__40448\,
            I => \N__40437\
        );

    \I__7577\ : InMux
    port map (
            O => \N__40447\,
            I => \N__40430\
        );

    \I__7576\ : InMux
    port map (
            O => \N__40446\,
            I => \N__40430\
        );

    \I__7575\ : InMux
    port map (
            O => \N__40445\,
            I => \N__40430\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__40440\,
            I => \c0.data_out_frame_29_7_N_1483_1\
        );

    \I__7573\ : Odrv4
    port map (
            O => \N__40437\,
            I => \c0.data_out_frame_29_7_N_1483_1\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__40430\,
            I => \c0.data_out_frame_29_7_N_1483_1\
        );

    \I__7571\ : CascadeMux
    port map (
            O => \N__40423\,
            I => \c0.n4_adj_4328_cascade_\
        );

    \I__7570\ : InMux
    port map (
            O => \N__40420\,
            I => \N__40415\
        );

    \I__7569\ : InMux
    port map (
            O => \N__40419\,
            I => \N__40412\
        );

    \I__7568\ : InMux
    port map (
            O => \N__40418\,
            I => \N__40409\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__40415\,
            I => \c0.data_out_frame_0__7__N_2568\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__40412\,
            I => \c0.data_out_frame_0__7__N_2568\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__40409\,
            I => \c0.data_out_frame_0__7__N_2568\
        );

    \I__7564\ : InMux
    port map (
            O => \N__40402\,
            I => \N__40396\
        );

    \I__7563\ : InMux
    port map (
            O => \N__40401\,
            I => \N__40396\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__40396\,
            I => \c0.FRAME_MATCHER_state_1\
        );

    \I__7561\ : InMux
    port map (
            O => \N__40393\,
            I => \N__40390\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__40390\,
            I => \N__40387\
        );

    \I__7559\ : Span4Mux_h
    port map (
            O => \N__40387\,
            I => \N__40384\
        );

    \I__7558\ : Odrv4
    port map (
            O => \N__40384\,
            I => \c0.n4_adj_4391\
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__40381\,
            I => \N__40378\
        );

    \I__7556\ : InMux
    port map (
            O => \N__40378\,
            I => \N__40375\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__40375\,
            I => \N__40372\
        );

    \I__7554\ : Odrv12
    port map (
            O => \N__40372\,
            I => \c0.n38_adj_4390\
        );

    \I__7553\ : InMux
    port map (
            O => \N__40369\,
            I => \N__40363\
        );

    \I__7552\ : InMux
    port map (
            O => \N__40368\,
            I => \N__40360\
        );

    \I__7551\ : CascadeMux
    port map (
            O => \N__40367\,
            I => \N__40356\
        );

    \I__7550\ : CascadeMux
    port map (
            O => \N__40366\,
            I => \N__40352\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__40363\,
            I => \N__40349\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__40360\,
            I => \N__40346\
        );

    \I__7547\ : InMux
    port map (
            O => \N__40359\,
            I => \N__40343\
        );

    \I__7546\ : InMux
    port map (
            O => \N__40356\,
            I => \N__40340\
        );

    \I__7545\ : InMux
    port map (
            O => \N__40355\,
            I => \N__40337\
        );

    \I__7544\ : InMux
    port map (
            O => \N__40352\,
            I => \N__40334\
        );

    \I__7543\ : Span4Mux_v
    port map (
            O => \N__40349\,
            I => \N__40331\
        );

    \I__7542\ : Span4Mux_h
    port map (
            O => \N__40346\,
            I => \N__40328\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__40343\,
            I => \N__40325\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__40340\,
            I => encoder0_position_23
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__40337\,
            I => encoder0_position_23
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__40334\,
            I => encoder0_position_23
        );

    \I__7537\ : Odrv4
    port map (
            O => \N__40331\,
            I => encoder0_position_23
        );

    \I__7536\ : Odrv4
    port map (
            O => \N__40328\,
            I => encoder0_position_23
        );

    \I__7535\ : Odrv12
    port map (
            O => \N__40325\,
            I => encoder0_position_23
        );

    \I__7534\ : CascadeMux
    port map (
            O => \N__40312\,
            I => \N__40309\
        );

    \I__7533\ : InMux
    port map (
            O => \N__40309\,
            I => \N__40306\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__40306\,
            I => \N__40301\
        );

    \I__7531\ : InMux
    port map (
            O => \N__40305\,
            I => \N__40298\
        );

    \I__7530\ : InMux
    port map (
            O => \N__40304\,
            I => \N__40295\
        );

    \I__7529\ : Span4Mux_h
    port map (
            O => \N__40301\,
            I => \N__40291\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__40298\,
            I => \N__40288\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__40295\,
            I => \N__40285\
        );

    \I__7526\ : CascadeMux
    port map (
            O => \N__40294\,
            I => \N__40281\
        );

    \I__7525\ : Span4Mux_h
    port map (
            O => \N__40291\,
            I => \N__40276\
        );

    \I__7524\ : Span4Mux_h
    port map (
            O => \N__40288\,
            I => \N__40276\
        );

    \I__7523\ : Span4Mux_v
    port map (
            O => \N__40285\,
            I => \N__40273\
        );

    \I__7522\ : InMux
    port map (
            O => \N__40284\,
            I => \N__40268\
        );

    \I__7521\ : InMux
    port map (
            O => \N__40281\,
            I => \N__40268\
        );

    \I__7520\ : Odrv4
    port map (
            O => \N__40276\,
            I => encoder0_position_8
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__40273\,
            I => encoder0_position_8
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__40268\,
            I => encoder0_position_8
        );

    \I__7517\ : InMux
    port map (
            O => \N__40261\,
            I => \N__40258\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__40258\,
            I => \N__40254\
        );

    \I__7515\ : InMux
    port map (
            O => \N__40257\,
            I => \N__40251\
        );

    \I__7514\ : Span4Mux_v
    port map (
            O => \N__40254\,
            I => \N__40246\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__40251\,
            I => \N__40246\
        );

    \I__7512\ : Odrv4
    port map (
            O => \N__40246\,
            I => \c0.n22032\
        );

    \I__7511\ : InMux
    port map (
            O => \N__40243\,
            I => \N__40238\
        );

    \I__7510\ : InMux
    port map (
            O => \N__40242\,
            I => \N__40233\
        );

    \I__7509\ : InMux
    port map (
            O => \N__40241\,
            I => \N__40233\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__40238\,
            I => \N__40229\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__40233\,
            I => \N__40226\
        );

    \I__7506\ : InMux
    port map (
            O => \N__40232\,
            I => \N__40223\
        );

    \I__7505\ : Span4Mux_v
    port map (
            O => \N__40229\,
            I => \N__40218\
        );

    \I__7504\ : Span4Mux_h
    port map (
            O => \N__40226\,
            I => \N__40218\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__40223\,
            I => data_in_3_0
        );

    \I__7502\ : Odrv4
    port map (
            O => \N__40218\,
            I => data_in_3_0
        );

    \I__7501\ : InMux
    port map (
            O => \N__40213\,
            I => \N__40210\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__40210\,
            I => \N__40205\
        );

    \I__7499\ : InMux
    port map (
            O => \N__40209\,
            I => \N__40202\
        );

    \I__7498\ : InMux
    port map (
            O => \N__40208\,
            I => \N__40199\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__40205\,
            I => \N__40195\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__40202\,
            I => \N__40192\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__40199\,
            I => \N__40189\
        );

    \I__7494\ : InMux
    port map (
            O => \N__40198\,
            I => \N__40186\
        );

    \I__7493\ : Span4Mux_h
    port map (
            O => \N__40195\,
            I => \N__40179\
        );

    \I__7492\ : Span4Mux_v
    port map (
            O => \N__40192\,
            I => \N__40179\
        );

    \I__7491\ : Span4Mux_v
    port map (
            O => \N__40189\,
            I => \N__40179\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__40186\,
            I => control_mode_5
        );

    \I__7489\ : Odrv4
    port map (
            O => \N__40179\,
            I => control_mode_5
        );

    \I__7488\ : CascadeMux
    port map (
            O => \N__40174\,
            I => \c0.n23215_cascade_\
        );

    \I__7487\ : InMux
    port map (
            O => \N__40171\,
            I => \N__40166\
        );

    \I__7486\ : InMux
    port map (
            O => \N__40170\,
            I => \N__40163\
        );

    \I__7485\ : InMux
    port map (
            O => \N__40169\,
            I => \N__40160\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__40166\,
            I => \N__40154\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__40163\,
            I => \N__40151\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__40160\,
            I => \N__40146\
        );

    \I__7481\ : InMux
    port map (
            O => \N__40159\,
            I => \N__40143\
        );

    \I__7480\ : InMux
    port map (
            O => \N__40158\,
            I => \N__40138\
        );

    \I__7479\ : InMux
    port map (
            O => \N__40157\,
            I => \N__40138\
        );

    \I__7478\ : Span4Mux_v
    port map (
            O => \N__40154\,
            I => \N__40133\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__40151\,
            I => \N__40133\
        );

    \I__7476\ : InMux
    port map (
            O => \N__40150\,
            I => \N__40128\
        );

    \I__7475\ : InMux
    port map (
            O => \N__40149\,
            I => \N__40128\
        );

    \I__7474\ : Span4Mux_h
    port map (
            O => \N__40146\,
            I => \N__40125\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__40143\,
            I => \N__40120\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__40138\,
            I => \N__40120\
        );

    \I__7471\ : Span4Mux_h
    port map (
            O => \N__40133\,
            I => \N__40115\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__40128\,
            I => \N__40115\
        );

    \I__7469\ : Span4Mux_h
    port map (
            O => \N__40125\,
            I => \N__40110\
        );

    \I__7468\ : Span4Mux_v
    port map (
            O => \N__40120\,
            I => \N__40107\
        );

    \I__7467\ : Span4Mux_h
    port map (
            O => \N__40115\,
            I => \N__40104\
        );

    \I__7466\ : InMux
    port map (
            O => \N__40114\,
            I => \N__40099\
        );

    \I__7465\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40099\
        );

    \I__7464\ : Odrv4
    port map (
            O => \N__40110\,
            I => \data_out_frame_29_7_N_1483_2\
        );

    \I__7463\ : Odrv4
    port map (
            O => \N__40107\,
            I => \data_out_frame_29_7_N_1483_2\
        );

    \I__7462\ : Odrv4
    port map (
            O => \N__40104\,
            I => \data_out_frame_29_7_N_1483_2\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__40099\,
            I => \data_out_frame_29_7_N_1483_2\
        );

    \I__7460\ : InMux
    port map (
            O => \N__40090\,
            I => \N__40087\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__40087\,
            I => \c0.n6_adj_4338\
        );

    \I__7458\ : CascadeMux
    port map (
            O => \N__40084\,
            I => \c0.n17602_cascade_\
        );

    \I__7457\ : InMux
    port map (
            O => \N__40081\,
            I => \N__40078\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__40078\,
            I => \c0.n8_adj_4417\
        );

    \I__7455\ : InMux
    port map (
            O => \N__40075\,
            I => \N__40072\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__40072\,
            I => \N__40069\
        );

    \I__7453\ : Span4Mux_h
    port map (
            O => \N__40069\,
            I => \N__40066\
        );

    \I__7452\ : Odrv4
    port map (
            O => \N__40066\,
            I => n2245
        );

    \I__7451\ : InMux
    port map (
            O => \N__40063\,
            I => \N__40060\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__40060\,
            I => \N__40053\
        );

    \I__7449\ : InMux
    port map (
            O => \N__40059\,
            I => \N__40050\
        );

    \I__7448\ : InMux
    port map (
            O => \N__40058\,
            I => \N__40047\
        );

    \I__7447\ : InMux
    port map (
            O => \N__40057\,
            I => \N__40044\
        );

    \I__7446\ : InMux
    port map (
            O => \N__40056\,
            I => \N__40041\
        );

    \I__7445\ : Span4Mux_v
    port map (
            O => \N__40053\,
            I => \N__40036\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__40050\,
            I => \N__40033\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__40047\,
            I => \N__40028\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__40044\,
            I => \N__40028\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__40041\,
            I => \N__40025\
        );

    \I__7440\ : InMux
    port map (
            O => \N__40040\,
            I => \N__40022\
        );

    \I__7439\ : InMux
    port map (
            O => \N__40039\,
            I => \N__40019\
        );

    \I__7438\ : Span4Mux_h
    port map (
            O => \N__40036\,
            I => \N__40014\
        );

    \I__7437\ : Span4Mux_v
    port map (
            O => \N__40033\,
            I => \N__40014\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__40028\,
            I => \N__40011\
        );

    \I__7435\ : Span12Mux_h
    port map (
            O => \N__40025\,
            I => \N__40008\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__40022\,
            I => \N__40005\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__40019\,
            I => encoder0_position_26
        );

    \I__7432\ : Odrv4
    port map (
            O => \N__40014\,
            I => encoder0_position_26
        );

    \I__7431\ : Odrv4
    port map (
            O => \N__40011\,
            I => encoder0_position_26
        );

    \I__7430\ : Odrv12
    port map (
            O => \N__40008\,
            I => encoder0_position_26
        );

    \I__7429\ : Odrv4
    port map (
            O => \N__40005\,
            I => encoder0_position_26
        );

    \I__7428\ : InMux
    port map (
            O => \N__39994\,
            I => \N__39991\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__39991\,
            I => \N__39988\
        );

    \I__7426\ : Span4Mux_v
    port map (
            O => \N__39988\,
            I => \N__39985\
        );

    \I__7425\ : Sp12to4
    port map (
            O => \N__39985\,
            I => \N__39982\
        );

    \I__7424\ : Odrv12
    port map (
            O => \N__39982\,
            I => n2263
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__39979\,
            I => \N__39976\
        );

    \I__7422\ : InMux
    port map (
            O => \N__39976\,
            I => \N__39971\
        );

    \I__7421\ : InMux
    port map (
            O => \N__39975\,
            I => \N__39968\
        );

    \I__7420\ : InMux
    port map (
            O => \N__39974\,
            I => \N__39963\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__39971\,
            I => \N__39960\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__39968\,
            I => \N__39957\
        );

    \I__7417\ : InMux
    port map (
            O => \N__39967\,
            I => \N__39952\
        );

    \I__7416\ : InMux
    port map (
            O => \N__39966\,
            I => \N__39952\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__39963\,
            I => encoder0_position_10
        );

    \I__7414\ : Odrv12
    port map (
            O => \N__39960\,
            I => encoder0_position_10
        );

    \I__7413\ : Odrv4
    port map (
            O => \N__39957\,
            I => encoder0_position_10
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__39952\,
            I => encoder0_position_10
        );

    \I__7411\ : CascadeMux
    port map (
            O => \N__39943\,
            I => \N__39940\
        );

    \I__7410\ : InMux
    port map (
            O => \N__39940\,
            I => \N__39937\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__39937\,
            I => \N__39934\
        );

    \I__7408\ : Span4Mux_h
    port map (
            O => \N__39934\,
            I => \N__39930\
        );

    \I__7407\ : InMux
    port map (
            O => \N__39933\,
            I => \N__39927\
        );

    \I__7406\ : Span4Mux_h
    port map (
            O => \N__39930\,
            I => \N__39924\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__39927\,
            I => data_out_frame_8_2
        );

    \I__7404\ : Odrv4
    port map (
            O => \N__39924\,
            I => data_out_frame_8_2
        );

    \I__7403\ : InMux
    port map (
            O => \N__39919\,
            I => \N__39916\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__39916\,
            I => \N__39913\
        );

    \I__7401\ : Span4Mux_h
    port map (
            O => \N__39913\,
            I => \N__39910\
        );

    \I__7400\ : Odrv4
    port map (
            O => \N__39910\,
            I => n2246
        );

    \I__7399\ : CascadeMux
    port map (
            O => \N__39907\,
            I => \N__39904\
        );

    \I__7398\ : InMux
    port map (
            O => \N__39904\,
            I => \N__39899\
        );

    \I__7397\ : InMux
    port map (
            O => \N__39903\,
            I => \N__39895\
        );

    \I__7396\ : CascadeMux
    port map (
            O => \N__39902\,
            I => \N__39890\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__39899\,
            I => \N__39886\
        );

    \I__7394\ : InMux
    port map (
            O => \N__39898\,
            I => \N__39883\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__39895\,
            I => \N__39880\
        );

    \I__7392\ : InMux
    port map (
            O => \N__39894\,
            I => \N__39875\
        );

    \I__7391\ : InMux
    port map (
            O => \N__39893\,
            I => \N__39875\
        );

    \I__7390\ : InMux
    port map (
            O => \N__39890\,
            I => \N__39872\
        );

    \I__7389\ : InMux
    port map (
            O => \N__39889\,
            I => \N__39869\
        );

    \I__7388\ : Span4Mux_h
    port map (
            O => \N__39886\,
            I => \N__39866\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__39883\,
            I => \N__39863\
        );

    \I__7386\ : Span4Mux_v
    port map (
            O => \N__39880\,
            I => \N__39858\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__39875\,
            I => \N__39858\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__39872\,
            I => encoder0_position_25
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__39869\,
            I => encoder0_position_25
        );

    \I__7382\ : Odrv4
    port map (
            O => \N__39866\,
            I => encoder0_position_25
        );

    \I__7381\ : Odrv12
    port map (
            O => \N__39863\,
            I => encoder0_position_25
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__39858\,
            I => encoder0_position_25
        );

    \I__7379\ : InMux
    port map (
            O => \N__39847\,
            I => \N__39841\
        );

    \I__7378\ : InMux
    port map (
            O => \N__39846\,
            I => \N__39841\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__39841\,
            I => data_out_frame_7_6
        );

    \I__7376\ : InMux
    port map (
            O => \N__39838\,
            I => \N__39829\
        );

    \I__7375\ : InMux
    port map (
            O => \N__39837\,
            I => \N__39826\
        );

    \I__7374\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39823\
        );

    \I__7373\ : InMux
    port map (
            O => \N__39835\,
            I => \N__39819\
        );

    \I__7372\ : InMux
    port map (
            O => \N__39834\,
            I => \N__39811\
        );

    \I__7371\ : InMux
    port map (
            O => \N__39833\,
            I => \N__39808\
        );

    \I__7370\ : InMux
    port map (
            O => \N__39832\,
            I => \N__39801\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__39829\,
            I => \N__39796\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__39826\,
            I => \N__39791\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__39823\,
            I => \N__39791\
        );

    \I__7366\ : InMux
    port map (
            O => \N__39822\,
            I => \N__39788\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__39819\,
            I => \N__39785\
        );

    \I__7364\ : InMux
    port map (
            O => \N__39818\,
            I => \N__39782\
        );

    \I__7363\ : InMux
    port map (
            O => \N__39817\,
            I => \N__39768\
        );

    \I__7362\ : InMux
    port map (
            O => \N__39816\,
            I => \N__39763\
        );

    \I__7361\ : InMux
    port map (
            O => \N__39815\,
            I => \N__39763\
        );

    \I__7360\ : InMux
    port map (
            O => \N__39814\,
            I => \N__39760\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__39811\,
            I => \N__39751\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__39808\,
            I => \N__39751\
        );

    \I__7357\ : InMux
    port map (
            O => \N__39807\,
            I => \N__39744\
        );

    \I__7356\ : InMux
    port map (
            O => \N__39806\,
            I => \N__39744\
        );

    \I__7355\ : InMux
    port map (
            O => \N__39805\,
            I => \N__39741\
        );

    \I__7354\ : InMux
    port map (
            O => \N__39804\,
            I => \N__39738\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__39801\,
            I => \N__39735\
        );

    \I__7352\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39727\
        );

    \I__7351\ : InMux
    port map (
            O => \N__39799\,
            I => \N__39727\
        );

    \I__7350\ : Span4Mux_v
    port map (
            O => \N__39796\,
            I => \N__39721\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__39791\,
            I => \N__39721\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__39788\,
            I => \N__39715\
        );

    \I__7347\ : Span4Mux_h
    port map (
            O => \N__39785\,
            I => \N__39715\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__39782\,
            I => \N__39712\
        );

    \I__7345\ : InMux
    port map (
            O => \N__39781\,
            I => \N__39709\
        );

    \I__7344\ : InMux
    port map (
            O => \N__39780\,
            I => \N__39702\
        );

    \I__7343\ : InMux
    port map (
            O => \N__39779\,
            I => \N__39702\
        );

    \I__7342\ : InMux
    port map (
            O => \N__39778\,
            I => \N__39702\
        );

    \I__7341\ : InMux
    port map (
            O => \N__39777\,
            I => \N__39697\
        );

    \I__7340\ : InMux
    port map (
            O => \N__39776\,
            I => \N__39690\
        );

    \I__7339\ : InMux
    port map (
            O => \N__39775\,
            I => \N__39690\
        );

    \I__7338\ : InMux
    port map (
            O => \N__39774\,
            I => \N__39690\
        );

    \I__7337\ : InMux
    port map (
            O => \N__39773\,
            I => \N__39687\
        );

    \I__7336\ : InMux
    port map (
            O => \N__39772\,
            I => \N__39682\
        );

    \I__7335\ : InMux
    port map (
            O => \N__39771\,
            I => \N__39682\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__39768\,
            I => \N__39679\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__39763\,
            I => \N__39676\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__39760\,
            I => \N__39673\
        );

    \I__7331\ : InMux
    port map (
            O => \N__39759\,
            I => \N__39668\
        );

    \I__7330\ : InMux
    port map (
            O => \N__39758\,
            I => \N__39668\
        );

    \I__7329\ : InMux
    port map (
            O => \N__39757\,
            I => \N__39663\
        );

    \I__7328\ : InMux
    port map (
            O => \N__39756\,
            I => \N__39663\
        );

    \I__7327\ : Span4Mux_v
    port map (
            O => \N__39751\,
            I => \N__39660\
        );

    \I__7326\ : InMux
    port map (
            O => \N__39750\,
            I => \N__39655\
        );

    \I__7325\ : InMux
    port map (
            O => \N__39749\,
            I => \N__39655\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__39744\,
            I => \N__39650\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__39741\,
            I => \N__39650\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__39738\,
            I => \N__39647\
        );

    \I__7321\ : Span4Mux_h
    port map (
            O => \N__39735\,
            I => \N__39644\
        );

    \I__7320\ : InMux
    port map (
            O => \N__39734\,
            I => \N__39639\
        );

    \I__7319\ : InMux
    port map (
            O => \N__39733\,
            I => \N__39639\
        );

    \I__7318\ : InMux
    port map (
            O => \N__39732\,
            I => \N__39636\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__39727\,
            I => \N__39633\
        );

    \I__7316\ : InMux
    port map (
            O => \N__39726\,
            I => \N__39630\
        );

    \I__7315\ : Sp12to4
    port map (
            O => \N__39721\,
            I => \N__39627\
        );

    \I__7314\ : CascadeMux
    port map (
            O => \N__39720\,
            I => \N__39623\
        );

    \I__7313\ : Span4Mux_v
    port map (
            O => \N__39715\,
            I => \N__39616\
        );

    \I__7312\ : Span4Mux_h
    port map (
            O => \N__39712\,
            I => \N__39616\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__39709\,
            I => \N__39616\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__39702\,
            I => \N__39613\
        );

    \I__7309\ : InMux
    port map (
            O => \N__39701\,
            I => \N__39608\
        );

    \I__7308\ : InMux
    port map (
            O => \N__39700\,
            I => \N__39608\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__39697\,
            I => \N__39603\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__39690\,
            I => \N__39603\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__39687\,
            I => \N__39598\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__39682\,
            I => \N__39598\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__39679\,
            I => \N__39591\
        );

    \I__7302\ : Span4Mux_v
    port map (
            O => \N__39676\,
            I => \N__39591\
        );

    \I__7301\ : Span4Mux_v
    port map (
            O => \N__39673\,
            I => \N__39591\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__39668\,
            I => \N__39586\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__39663\,
            I => \N__39586\
        );

    \I__7298\ : Span4Mux_h
    port map (
            O => \N__39660\,
            I => \N__39583\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__39655\,
            I => \N__39574\
        );

    \I__7296\ : Span4Mux_v
    port map (
            O => \N__39650\,
            I => \N__39574\
        );

    \I__7295\ : Span4Mux_v
    port map (
            O => \N__39647\,
            I => \N__39574\
        );

    \I__7294\ : Span4Mux_h
    port map (
            O => \N__39644\,
            I => \N__39574\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__39639\,
            I => \N__39569\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__39636\,
            I => \N__39569\
        );

    \I__7291\ : Span4Mux_v
    port map (
            O => \N__39633\,
            I => \N__39564\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__39630\,
            I => \N__39564\
        );

    \I__7289\ : Span12Mux_h
    port map (
            O => \N__39627\,
            I => \N__39561\
        );

    \I__7288\ : InMux
    port map (
            O => \N__39626\,
            I => \N__39558\
        );

    \I__7287\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39555\
        );

    \I__7286\ : Span4Mux_h
    port map (
            O => \N__39616\,
            I => \N__39552\
        );

    \I__7285\ : Span4Mux_v
    port map (
            O => \N__39613\,
            I => \N__39541\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__39608\,
            I => \N__39541\
        );

    \I__7283\ : Span4Mux_v
    port map (
            O => \N__39603\,
            I => \N__39541\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__39598\,
            I => \N__39541\
        );

    \I__7281\ : Span4Mux_h
    port map (
            O => \N__39591\,
            I => \N__39541\
        );

    \I__7280\ : Span4Mux_h
    port map (
            O => \N__39586\,
            I => \N__39534\
        );

    \I__7279\ : Span4Mux_v
    port map (
            O => \N__39583\,
            I => \N__39534\
        );

    \I__7278\ : Span4Mux_h
    port map (
            O => \N__39574\,
            I => \N__39534\
        );

    \I__7277\ : Span12Mux_v
    port map (
            O => \N__39569\,
            I => \N__39525\
        );

    \I__7276\ : Sp12to4
    port map (
            O => \N__39564\,
            I => \N__39525\
        );

    \I__7275\ : Span12Mux_v
    port map (
            O => \N__39561\,
            I => \N__39525\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__39558\,
            I => \N__39525\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__39555\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7272\ : Odrv4
    port map (
            O => \N__39552\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7271\ : Odrv4
    port map (
            O => \N__39541\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7270\ : Odrv4
    port map (
            O => \N__39534\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7269\ : Odrv12
    port map (
            O => \N__39525\,
            I => \c0.byte_transmit_counter_0\
        );

    \I__7268\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39511\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__39511\,
            I => \N__39508\
        );

    \I__7266\ : Span4Mux_v
    port map (
            O => \N__39508\,
            I => \N__39505\
        );

    \I__7265\ : Span4Mux_h
    port map (
            O => \N__39505\,
            I => \N__39502\
        );

    \I__7264\ : Odrv4
    port map (
            O => \N__39502\,
            I => \c0.n5_adj_4350\
        );

    \I__7263\ : InMux
    port map (
            O => \N__39499\,
            I => \N__39496\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__39496\,
            I => \N__39492\
        );

    \I__7261\ : InMux
    port map (
            O => \N__39495\,
            I => \N__39489\
        );

    \I__7260\ : Span4Mux_v
    port map (
            O => \N__39492\,
            I => \N__39481\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__39489\,
            I => \N__39481\
        );

    \I__7258\ : InMux
    port map (
            O => \N__39488\,
            I => \N__39478\
        );

    \I__7257\ : InMux
    port map (
            O => \N__39487\,
            I => \N__39472\
        );

    \I__7256\ : InMux
    port map (
            O => \N__39486\,
            I => \N__39469\
        );

    \I__7255\ : Span4Mux_h
    port map (
            O => \N__39481\,
            I => \N__39466\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__39478\,
            I => \N__39463\
        );

    \I__7253\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39458\
        );

    \I__7252\ : InMux
    port map (
            O => \N__39476\,
            I => \N__39458\
        );

    \I__7251\ : InMux
    port map (
            O => \N__39475\,
            I => \N__39455\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__39472\,
            I => \N__39452\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__39469\,
            I => \N__39447\
        );

    \I__7248\ : Span4Mux_v
    port map (
            O => \N__39466\,
            I => \N__39447\
        );

    \I__7247\ : Span12Mux_h
    port map (
            O => \N__39463\,
            I => \N__39440\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__39458\,
            I => \N__39440\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__39455\,
            I => \N__39440\
        );

    \I__7244\ : Odrv12
    port map (
            O => \N__39452\,
            I => control_mode_2
        );

    \I__7243\ : Odrv4
    port map (
            O => \N__39447\,
            I => control_mode_2
        );

    \I__7242\ : Odrv12
    port map (
            O => \N__39440\,
            I => control_mode_2
        );

    \I__7241\ : CascadeMux
    port map (
            O => \N__39433\,
            I => \c0.n6_adj_4315_cascade_\
        );

    \I__7240\ : InMux
    port map (
            O => \N__39430\,
            I => \N__39427\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__39427\,
            I => \N__39423\
        );

    \I__7238\ : InMux
    port map (
            O => \N__39426\,
            I => \N__39420\
        );

    \I__7237\ : Span4Mux_h
    port map (
            O => \N__39423\,
            I => \N__39417\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__39420\,
            I => \N__39414\
        );

    \I__7235\ : Span4Mux_v
    port map (
            O => \N__39417\,
            I => \N__39411\
        );

    \I__7234\ : Span4Mux_v
    port map (
            O => \N__39414\,
            I => \N__39408\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__39411\,
            I => \c0.n20171\
        );

    \I__7232\ : Odrv4
    port map (
            O => \N__39408\,
            I => \c0.n20171\
        );

    \I__7231\ : InMux
    port map (
            O => \N__39403\,
            I => \N__39400\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__39400\,
            I => \c0.data_out_frame_29__7__N_847\
        );

    \I__7229\ : CascadeMux
    port map (
            O => \N__39397\,
            I => \c0.data_out_frame_29__7__N_847_cascade_\
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__39394\,
            I => \N__39387\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__39393\,
            I => \N__39384\
        );

    \I__7226\ : CascadeMux
    port map (
            O => \N__39392\,
            I => \N__39381\
        );

    \I__7225\ : CascadeMux
    port map (
            O => \N__39391\,
            I => \N__39378\
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__39390\,
            I => \N__39375\
        );

    \I__7223\ : InMux
    port map (
            O => \N__39387\,
            I => \N__39372\
        );

    \I__7222\ : InMux
    port map (
            O => \N__39384\,
            I => \N__39367\
        );

    \I__7221\ : InMux
    port map (
            O => \N__39381\,
            I => \N__39367\
        );

    \I__7220\ : InMux
    port map (
            O => \N__39378\,
            I => \N__39364\
        );

    \I__7219\ : InMux
    port map (
            O => \N__39375\,
            I => \N__39361\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__39372\,
            I => \N__39355\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__39367\,
            I => \N__39355\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__39364\,
            I => \N__39350\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__39361\,
            I => \N__39350\
        );

    \I__7214\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39347\
        );

    \I__7213\ : Odrv4
    port map (
            O => \N__39355\,
            I => encoder0_position_11
        );

    \I__7212\ : Odrv12
    port map (
            O => \N__39350\,
            I => encoder0_position_11
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__39347\,
            I => encoder0_position_11
        );

    \I__7210\ : InMux
    port map (
            O => \N__39340\,
            I => \N__39337\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__39337\,
            I => \c0.n10_adj_4332\
        );

    \I__7208\ : CascadeMux
    port map (
            O => \N__39334\,
            I => \N__39331\
        );

    \I__7207\ : InMux
    port map (
            O => \N__39331\,
            I => \N__39328\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__39328\,
            I => \N__39325\
        );

    \I__7205\ : Span4Mux_h
    port map (
            O => \N__39325\,
            I => \N__39321\
        );

    \I__7204\ : InMux
    port map (
            O => \N__39324\,
            I => \N__39314\
        );

    \I__7203\ : Span4Mux_h
    port map (
            O => \N__39321\,
            I => \N__39311\
        );

    \I__7202\ : InMux
    port map (
            O => \N__39320\,
            I => \N__39308\
        );

    \I__7201\ : InMux
    port map (
            O => \N__39319\,
            I => \N__39301\
        );

    \I__7200\ : InMux
    port map (
            O => \N__39318\,
            I => \N__39301\
        );

    \I__7199\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39301\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__39314\,
            I => encoder0_position_24
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__39311\,
            I => encoder0_position_24
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__39308\,
            I => encoder0_position_24
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__39301\,
            I => encoder0_position_24
        );

    \I__7194\ : InMux
    port map (
            O => \N__39292\,
            I => \N__39289\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__39289\,
            I => \N__39285\
        );

    \I__7192\ : InMux
    port map (
            O => \N__39288\,
            I => \N__39282\
        );

    \I__7191\ : Span12Mux_v
    port map (
            O => \N__39285\,
            I => \N__39279\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__39282\,
            I => \c0.n21931\
        );

    \I__7189\ : Odrv12
    port map (
            O => \N__39279\,
            I => \c0.n21931\
        );

    \I__7188\ : InMux
    port map (
            O => \N__39274\,
            I => \N__39270\
        );

    \I__7187\ : InMux
    port map (
            O => \N__39273\,
            I => \N__39265\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__39270\,
            I => \N__39261\
        );

    \I__7185\ : InMux
    port map (
            O => \N__39269\,
            I => \N__39258\
        );

    \I__7184\ : InMux
    port map (
            O => \N__39268\,
            I => \N__39255\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__39265\,
            I => \N__39252\
        );

    \I__7182\ : InMux
    port map (
            O => \N__39264\,
            I => \N__39249\
        );

    \I__7181\ : Span4Mux_h
    port map (
            O => \N__39261\,
            I => \N__39243\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__39258\,
            I => \N__39243\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__39255\,
            I => \N__39236\
        );

    \I__7178\ : Span4Mux_v
    port map (
            O => \N__39252\,
            I => \N__39236\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__39249\,
            I => \N__39236\
        );

    \I__7176\ : InMux
    port map (
            O => \N__39248\,
            I => \N__39233\
        );

    \I__7175\ : Span4Mux_v
    port map (
            O => \N__39243\,
            I => \N__39230\
        );

    \I__7174\ : Span4Mux_h
    port map (
            O => \N__39236\,
            I => \N__39225\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__39233\,
            I => \N__39225\
        );

    \I__7172\ : Odrv4
    port map (
            O => \N__39230\,
            I => \c0.r_SM_Main_2_N_3755_0\
        );

    \I__7171\ : Odrv4
    port map (
            O => \N__39225\,
            I => \c0.r_SM_Main_2_N_3755_0\
        );

    \I__7170\ : CEMux
    port map (
            O => \N__39220\,
            I => \N__39217\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__39217\,
            I => \N__39214\
        );

    \I__7168\ : Span4Mux_h
    port map (
            O => \N__39214\,
            I => \N__39211\
        );

    \I__7167\ : Span4Mux_h
    port map (
            O => \N__39211\,
            I => \N__39208\
        );

    \I__7166\ : Odrv4
    port map (
            O => \N__39208\,
            I => \c0.n14322\
        );

    \I__7165\ : CascadeMux
    port map (
            O => \N__39205\,
            I => \c0.n14322_cascade_\
        );

    \I__7164\ : SRMux
    port map (
            O => \N__39202\,
            I => \N__39199\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__39199\,
            I => \N__39196\
        );

    \I__7162\ : Span12Mux_s8_h
    port map (
            O => \N__39196\,
            I => \N__39193\
        );

    \I__7161\ : Odrv12
    port map (
            O => \N__39193\,
            I => \c0.n14871\
        );

    \I__7160\ : CascadeMux
    port map (
            O => \N__39190\,
            I => \N__39186\
        );

    \I__7159\ : InMux
    port map (
            O => \N__39189\,
            I => \N__39183\
        );

    \I__7158\ : InMux
    port map (
            O => \N__39186\,
            I => \N__39180\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__39183\,
            I => \N__39177\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__39180\,
            I => \N__39174\
        );

    \I__7155\ : Span4Mux_h
    port map (
            O => \N__39177\,
            I => \N__39171\
        );

    \I__7154\ : Odrv12
    port map (
            O => \N__39174\,
            I => \c0.tx_transmit_N_3651\
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__39171\,
            I => \c0.tx_transmit_N_3651\
        );

    \I__7152\ : InMux
    port map (
            O => \N__39166\,
            I => \N__39163\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__39163\,
            I => \c0.n23975\
        );

    \I__7150\ : InMux
    port map (
            O => \N__39160\,
            I => \N__39157\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__39157\,
            I => \N__39154\
        );

    \I__7148\ : Span4Mux_v
    port map (
            O => \N__39154\,
            I => \N__39151\
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__39151\,
            I => \c0.n18_adj_4403\
        );

    \I__7146\ : InMux
    port map (
            O => \N__39148\,
            I => \N__39145\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__39145\,
            I => \N__39142\
        );

    \I__7144\ : Odrv12
    port map (
            O => \N__39142\,
            I => \c0.n20875\
        );

    \I__7143\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39135\
        );

    \I__7142\ : InMux
    port map (
            O => \N__39138\,
            I => \N__39132\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__39135\,
            I => \c0.n17602\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__39132\,
            I => \c0.n17602\
        );

    \I__7139\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39124\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__39124\,
            I => \N__39121\
        );

    \I__7137\ : Span4Mux_v
    port map (
            O => \N__39121\,
            I => \N__39118\
        );

    \I__7136\ : Odrv4
    port map (
            O => \N__39118\,
            I => n2255
        );

    \I__7135\ : InMux
    port map (
            O => \N__39115\,
            I => \N__39111\
        );

    \I__7134\ : CascadeMux
    port map (
            O => \N__39114\,
            I => \N__39108\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__39111\,
            I => \N__39105\
        );

    \I__7132\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39102\
        );

    \I__7131\ : Span4Mux_v
    port map (
            O => \N__39105\,
            I => \N__39098\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__39102\,
            I => \N__39095\
        );

    \I__7129\ : InMux
    port map (
            O => \N__39101\,
            I => \N__39092\
        );

    \I__7128\ : Span4Mux_h
    port map (
            O => \N__39098\,
            I => \N__39086\
        );

    \I__7127\ : Span4Mux_h
    port map (
            O => \N__39095\,
            I => \N__39081\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__39092\,
            I => \N__39081\
        );

    \I__7125\ : InMux
    port map (
            O => \N__39091\,
            I => \N__39078\
        );

    \I__7124\ : InMux
    port map (
            O => \N__39090\,
            I => \N__39073\
        );

    \I__7123\ : InMux
    port map (
            O => \N__39089\,
            I => \N__39073\
        );

    \I__7122\ : Odrv4
    port map (
            O => \N__39086\,
            I => encoder0_position_16
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__39081\,
            I => encoder0_position_16
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__39078\,
            I => encoder0_position_16
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__39073\,
            I => encoder0_position_16
        );

    \I__7118\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39061\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__39061\,
            I => \N__39057\
        );

    \I__7116\ : InMux
    port map (
            O => \N__39060\,
            I => \N__39053\
        );

    \I__7115\ : Span4Mux_h
    port map (
            O => \N__39057\,
            I => \N__39050\
        );

    \I__7114\ : InMux
    port map (
            O => \N__39056\,
            I => \N__39047\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__39053\,
            I => \c0.n22408\
        );

    \I__7112\ : Odrv4
    port map (
            O => \N__39050\,
            I => \c0.n22408\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__39047\,
            I => \c0.n22408\
        );

    \I__7110\ : InMux
    port map (
            O => \N__39040\,
            I => \N__39037\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__39037\,
            I => \N__39032\
        );

    \I__7108\ : InMux
    port map (
            O => \N__39036\,
            I => \N__39029\
        );

    \I__7107\ : InMux
    port map (
            O => \N__39035\,
            I => \N__39026\
        );

    \I__7106\ : Span4Mux_h
    port map (
            O => \N__39032\,
            I => \N__39023\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__39029\,
            I => \N__39020\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__39026\,
            I => \N__39017\
        );

    \I__7103\ : Span4Mux_v
    port map (
            O => \N__39023\,
            I => \N__39009\
        );

    \I__7102\ : Span4Mux_v
    port map (
            O => \N__39020\,
            I => \N__39009\
        );

    \I__7101\ : Span4Mux_h
    port map (
            O => \N__39017\,
            I => \N__39006\
        );

    \I__7100\ : InMux
    port map (
            O => \N__39016\,
            I => \N__39001\
        );

    \I__7099\ : InMux
    port map (
            O => \N__39015\,
            I => \N__39001\
        );

    \I__7098\ : InMux
    port map (
            O => \N__39014\,
            I => \N__38998\
        );

    \I__7097\ : Odrv4
    port map (
            O => \N__39009\,
            I => encoder0_position_4
        );

    \I__7096\ : Odrv4
    port map (
            O => \N__39006\,
            I => encoder0_position_4
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__39001\,
            I => encoder0_position_4
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__38998\,
            I => encoder0_position_4
        );

    \I__7093\ : CascadeMux
    port map (
            O => \N__38989\,
            I => \c0.n22227_cascade_\
        );

    \I__7092\ : InMux
    port map (
            O => \N__38986\,
            I => \N__38982\
        );

    \I__7091\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38979\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__38982\,
            I => \N__38976\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__38979\,
            I => \c0.n22128\
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__38976\,
            I => \c0.n22128\
        );

    \I__7087\ : CascadeMux
    port map (
            O => \N__38971\,
            I => \N__38968\
        );

    \I__7086\ : InMux
    port map (
            O => \N__38968\,
            I => \N__38958\
        );

    \I__7085\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38958\
        );

    \I__7084\ : InMux
    port map (
            O => \N__38966\,
            I => \N__38958\
        );

    \I__7083\ : InMux
    port map (
            O => \N__38965\,
            I => \N__38955\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__38958\,
            I => \N__38950\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__38955\,
            I => \N__38950\
        );

    \I__7080\ : Span4Mux_h
    port map (
            O => \N__38950\,
            I => \N__38947\
        );

    \I__7079\ : Span4Mux_v
    port map (
            O => \N__38947\,
            I => \N__38944\
        );

    \I__7078\ : Odrv4
    port map (
            O => \N__38944\,
            I => \c0.n10444\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__38941\,
            I => \N__38938\
        );

    \I__7076\ : InMux
    port map (
            O => \N__38938\,
            I => \N__38935\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__38935\,
            I => \N__38931\
        );

    \I__7074\ : CascadeMux
    port map (
            O => \N__38934\,
            I => \N__38928\
        );

    \I__7073\ : Span4Mux_h
    port map (
            O => \N__38931\,
            I => \N__38925\
        );

    \I__7072\ : InMux
    port map (
            O => \N__38928\,
            I => \N__38922\
        );

    \I__7071\ : Span4Mux_v
    port map (
            O => \N__38925\,
            I => \N__38917\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__38922\,
            I => \N__38917\
        );

    \I__7069\ : Span4Mux_h
    port map (
            O => \N__38917\,
            I => \N__38911\
        );

    \I__7068\ : InMux
    port map (
            O => \N__38916\,
            I => \N__38906\
        );

    \I__7067\ : InMux
    port map (
            O => \N__38915\,
            I => \N__38906\
        );

    \I__7066\ : InMux
    port map (
            O => \N__38914\,
            I => \N__38902\
        );

    \I__7065\ : Span4Mux_h
    port map (
            O => \N__38911\,
            I => \N__38897\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__38906\,
            I => \N__38897\
        );

    \I__7063\ : InMux
    port map (
            O => \N__38905\,
            I => \N__38894\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__38902\,
            I => encoder1_position_20
        );

    \I__7061\ : Odrv4
    port map (
            O => \N__38897\,
            I => encoder1_position_20
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__38894\,
            I => encoder1_position_20
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__38887\,
            I => \N__38884\
        );

    \I__7058\ : InMux
    port map (
            O => \N__38884\,
            I => \N__38881\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__38881\,
            I => \N__38878\
        );

    \I__7056\ : Odrv12
    port map (
            O => \N__38878\,
            I => \c0.n6_adj_4312\
        );

    \I__7055\ : InMux
    port map (
            O => \N__38875\,
            I => \N__38871\
        );

    \I__7054\ : InMux
    port map (
            O => \N__38874\,
            I => \N__38866\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__38871\,
            I => \N__38863\
        );

    \I__7052\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38860\
        );

    \I__7051\ : InMux
    port map (
            O => \N__38869\,
            I => \N__38856\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__38866\,
            I => \N__38851\
        );

    \I__7049\ : Span4Mux_h
    port map (
            O => \N__38863\,
            I => \N__38851\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__38860\,
            I => \N__38848\
        );

    \I__7047\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38844\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__38856\,
            I => \N__38841\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__38851\,
            I => \N__38838\
        );

    \I__7044\ : Span12Mux_h
    port map (
            O => \N__38848\,
            I => \N__38835\
        );

    \I__7043\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38832\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__38844\,
            I => encoder0_position_12
        );

    \I__7041\ : Odrv4
    port map (
            O => \N__38841\,
            I => encoder0_position_12
        );

    \I__7040\ : Odrv4
    port map (
            O => \N__38838\,
            I => encoder0_position_12
        );

    \I__7039\ : Odrv12
    port map (
            O => \N__38835\,
            I => encoder0_position_12
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__38832\,
            I => encoder0_position_12
        );

    \I__7037\ : InMux
    port map (
            O => \N__38821\,
            I => \N__38818\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__38818\,
            I => \N__38815\
        );

    \I__7035\ : Odrv4
    port map (
            O => \N__38815\,
            I => \c0.n22477\
        );

    \I__7034\ : CascadeMux
    port map (
            O => \N__38812\,
            I => \c0.n22477_cascade_\
        );

    \I__7033\ : InMux
    port map (
            O => \N__38809\,
            I => \N__38806\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__38806\,
            I => \N__38803\
        );

    \I__7031\ : Odrv4
    port map (
            O => \N__38803\,
            I => \c0.n6_adj_4333\
        );

    \I__7030\ : InMux
    port map (
            O => \N__38800\,
            I => \N__38797\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__38797\,
            I => \N__38794\
        );

    \I__7028\ : Span4Mux_h
    port map (
            O => \N__38794\,
            I => \N__38791\
        );

    \I__7027\ : Span4Mux_h
    port map (
            O => \N__38791\,
            I => \N__38788\
        );

    \I__7026\ : Odrv4
    port map (
            O => \N__38788\,
            I => n2243
        );

    \I__7025\ : CascadeMux
    port map (
            O => \N__38785\,
            I => \N__38780\
        );

    \I__7024\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38777\
        );

    \I__7023\ : InMux
    port map (
            O => \N__38783\,
            I => \N__38774\
        );

    \I__7022\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38768\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__38777\,
            I => \N__38765\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__38774\,
            I => \N__38762\
        );

    \I__7019\ : InMux
    port map (
            O => \N__38773\,
            I => \N__38757\
        );

    \I__7018\ : InMux
    port map (
            O => \N__38772\,
            I => \N__38757\
        );

    \I__7017\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38753\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__38768\,
            I => \N__38750\
        );

    \I__7015\ : Span4Mux_h
    port map (
            O => \N__38765\,
            I => \N__38745\
        );

    \I__7014\ : Span4Mux_h
    port map (
            O => \N__38762\,
            I => \N__38745\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__38757\,
            I => \N__38742\
        );

    \I__7012\ : InMux
    port map (
            O => \N__38756\,
            I => \N__38739\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__38753\,
            I => encoder0_position_28
        );

    \I__7010\ : Odrv4
    port map (
            O => \N__38750\,
            I => encoder0_position_28
        );

    \I__7009\ : Odrv4
    port map (
            O => \N__38745\,
            I => encoder0_position_28
        );

    \I__7008\ : Odrv4
    port map (
            O => \N__38742\,
            I => encoder0_position_28
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__38739\,
            I => encoder0_position_28
        );

    \I__7006\ : CascadeMux
    port map (
            O => \N__38728\,
            I => \N__38725\
        );

    \I__7005\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38719\
        );

    \I__7004\ : InMux
    port map (
            O => \N__38724\,
            I => \N__38716\
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__38723\,
            I => \N__38711\
        );

    \I__7002\ : InMux
    port map (
            O => \N__38722\,
            I => \N__38708\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__38719\,
            I => \N__38705\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__38716\,
            I => \N__38702\
        );

    \I__6999\ : InMux
    port map (
            O => \N__38715\,
            I => \N__38697\
        );

    \I__6998\ : InMux
    port map (
            O => \N__38714\,
            I => \N__38697\
        );

    \I__6997\ : InMux
    port map (
            O => \N__38711\,
            I => \N__38694\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__38708\,
            I => \N__38687\
        );

    \I__6995\ : Span4Mux_h
    port map (
            O => \N__38705\,
            I => \N__38687\
        );

    \I__6994\ : Span4Mux_h
    port map (
            O => \N__38702\,
            I => \N__38687\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__38697\,
            I => \N__38684\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__38694\,
            I => encoder0_position_9
        );

    \I__6991\ : Odrv4
    port map (
            O => \N__38687\,
            I => encoder0_position_9
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__38684\,
            I => encoder0_position_9
        );

    \I__6989\ : InMux
    port map (
            O => \N__38677\,
            I => \N__38671\
        );

    \I__6988\ : InMux
    port map (
            O => \N__38676\,
            I => \N__38671\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__38671\,
            I => \c0.n22427\
        );

    \I__6986\ : CascadeMux
    port map (
            O => \N__38668\,
            I => \N__38663\
        );

    \I__6985\ : InMux
    port map (
            O => \N__38667\,
            I => \N__38659\
        );

    \I__6984\ : InMux
    port map (
            O => \N__38666\,
            I => \N__38656\
        );

    \I__6983\ : InMux
    port map (
            O => \N__38663\,
            I => \N__38653\
        );

    \I__6982\ : CascadeMux
    port map (
            O => \N__38662\,
            I => \N__38649\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__38659\,
            I => \N__38645\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__38656\,
            I => \N__38642\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__38653\,
            I => \N__38639\
        );

    \I__6978\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38636\
        );

    \I__6977\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38633\
        );

    \I__6976\ : InMux
    port map (
            O => \N__38648\,
            I => \N__38630\
        );

    \I__6975\ : Span4Mux_h
    port map (
            O => \N__38645\,
            I => \N__38627\
        );

    \I__6974\ : Span4Mux_h
    port map (
            O => \N__38642\,
            I => \N__38622\
        );

    \I__6973\ : Span4Mux_h
    port map (
            O => \N__38639\,
            I => \N__38622\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__38636\,
            I => encoder0_position_19
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__38633\,
            I => encoder0_position_19
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__38630\,
            I => encoder0_position_19
        );

    \I__6969\ : Odrv4
    port map (
            O => \N__38627\,
            I => encoder0_position_19
        );

    \I__6968\ : Odrv4
    port map (
            O => \N__38622\,
            I => encoder0_position_19
        );

    \I__6967\ : CascadeMux
    port map (
            O => \N__38611\,
            I => \N__38607\
        );

    \I__6966\ : InMux
    port map (
            O => \N__38610\,
            I => \N__38602\
        );

    \I__6965\ : InMux
    port map (
            O => \N__38607\,
            I => \N__38602\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__38602\,
            I => \c0.n21885\
        );

    \I__6963\ : InMux
    port map (
            O => \N__38599\,
            I => \N__38596\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__38596\,
            I => \c0.n22200\
        );

    \I__6961\ : CascadeMux
    port map (
            O => \N__38593\,
            I => \c0.n22200_cascade_\
        );

    \I__6960\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38587\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__38587\,
            I => \N__38583\
        );

    \I__6958\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38580\
        );

    \I__6957\ : Span4Mux_h
    port map (
            O => \N__38583\,
            I => \N__38576\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__38580\,
            I => \N__38573\
        );

    \I__6955\ : InMux
    port map (
            O => \N__38579\,
            I => \N__38570\
        );

    \I__6954\ : Odrv4
    port map (
            O => \N__38576\,
            I => \c0.n21970\
        );

    \I__6953\ : Odrv12
    port map (
            O => \N__38573\,
            I => \c0.n21970\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__38570\,
            I => \c0.n21970\
        );

    \I__6951\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38560\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__38560\,
            I => \N__38557\
        );

    \I__6949\ : Span4Mux_h
    port map (
            O => \N__38557\,
            I => \N__38553\
        );

    \I__6948\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38550\
        );

    \I__6947\ : Odrv4
    port map (
            O => \N__38553\,
            I => \c0.n13705\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__38550\,
            I => \c0.n13705\
        );

    \I__6945\ : InMux
    port map (
            O => \N__38545\,
            I => \N__38542\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__38542\,
            I => \N__38539\
        );

    \I__6943\ : Odrv12
    port map (
            O => \N__38539\,
            I => n2259
        );

    \I__6942\ : InMux
    port map (
            O => \N__38536\,
            I => \N__38533\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__38533\,
            I => \N__38530\
        );

    \I__6940\ : Span4Mux_v
    port map (
            O => \N__38530\,
            I => \N__38527\
        );

    \I__6939\ : Odrv4
    port map (
            O => \N__38527\,
            I => n2267
        );

    \I__6938\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38521\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__38521\,
            I => \N__38518\
        );

    \I__6936\ : Odrv4
    port map (
            O => \N__38518\,
            I => n2261
        );

    \I__6935\ : InMux
    port map (
            O => \N__38515\,
            I => \N__38512\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__38512\,
            I => \N__38509\
        );

    \I__6933\ : Odrv12
    port map (
            O => \N__38509\,
            I => \c0.n21908\
        );

    \I__6932\ : InMux
    port map (
            O => \N__38506\,
            I => \N__38493\
        );

    \I__6931\ : InMux
    port map (
            O => \N__38505\,
            I => \N__38488\
        );

    \I__6930\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38485\
        );

    \I__6929\ : InMux
    port map (
            O => \N__38503\,
            I => \N__38482\
        );

    \I__6928\ : InMux
    port map (
            O => \N__38502\,
            I => \N__38473\
        );

    \I__6927\ : InMux
    port map (
            O => \N__38501\,
            I => \N__38473\
        );

    \I__6926\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38473\
        );

    \I__6925\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38473\
        );

    \I__6924\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38470\
        );

    \I__6923\ : InMux
    port map (
            O => \N__38497\,
            I => \N__38467\
        );

    \I__6922\ : CascadeMux
    port map (
            O => \N__38496\,
            I => \N__38462\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__38493\,
            I => \N__38454\
        );

    \I__6920\ : InMux
    port map (
            O => \N__38492\,
            I => \N__38449\
        );

    \I__6919\ : InMux
    port map (
            O => \N__38491\,
            I => \N__38449\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__38488\,
            I => \N__38446\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__38485\,
            I => \N__38443\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__38482\,
            I => \N__38434\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__38473\,
            I => \N__38434\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__38470\,
            I => \N__38434\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__38467\,
            I => \N__38434\
        );

    \I__6912\ : InMux
    port map (
            O => \N__38466\,
            I => \N__38431\
        );

    \I__6911\ : InMux
    port map (
            O => \N__38465\,
            I => \N__38424\
        );

    \I__6910\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38424\
        );

    \I__6909\ : InMux
    port map (
            O => \N__38461\,
            I => \N__38424\
        );

    \I__6908\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38419\
        );

    \I__6907\ : InMux
    port map (
            O => \N__38459\,
            I => \N__38419\
        );

    \I__6906\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38416\
        );

    \I__6905\ : InMux
    port map (
            O => \N__38457\,
            I => \N__38413\
        );

    \I__6904\ : Span4Mux_h
    port map (
            O => \N__38454\,
            I => \N__38405\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__38449\,
            I => \N__38405\
        );

    \I__6902\ : Span4Mux_v
    port map (
            O => \N__38446\,
            I => \N__38402\
        );

    \I__6901\ : Span4Mux_v
    port map (
            O => \N__38443\,
            I => \N__38397\
        );

    \I__6900\ : Span4Mux_v
    port map (
            O => \N__38434\,
            I => \N__38397\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__38431\,
            I => \N__38388\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__38424\,
            I => \N__38388\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__38419\,
            I => \N__38388\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__38416\,
            I => \N__38383\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__38413\,
            I => \N__38383\
        );

    \I__6894\ : InMux
    port map (
            O => \N__38412\,
            I => \N__38378\
        );

    \I__6893\ : InMux
    port map (
            O => \N__38411\,
            I => \N__38378\
        );

    \I__6892\ : CascadeMux
    port map (
            O => \N__38410\,
            I => \N__38374\
        );

    \I__6891\ : Span4Mux_v
    port map (
            O => \N__38405\,
            I => \N__38367\
        );

    \I__6890\ : Span4Mux_h
    port map (
            O => \N__38402\,
            I => \N__38367\
        );

    \I__6889\ : Span4Mux_h
    port map (
            O => \N__38397\,
            I => \N__38367\
        );

    \I__6888\ : InMux
    port map (
            O => \N__38396\,
            I => \N__38364\
        );

    \I__6887\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38361\
        );

    \I__6886\ : Span12Mux_v
    port map (
            O => \N__38388\,
            I => \N__38353\
        );

    \I__6885\ : Span4Mux_v
    port map (
            O => \N__38383\,
            I => \N__38348\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__38378\,
            I => \N__38348\
        );

    \I__6883\ : InMux
    port map (
            O => \N__38377\,
            I => \N__38343\
        );

    \I__6882\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38343\
        );

    \I__6881\ : Sp12to4
    port map (
            O => \N__38367\,
            I => \N__38336\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__38364\,
            I => \N__38336\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__38361\,
            I => \N__38336\
        );

    \I__6878\ : InMux
    port map (
            O => \N__38360\,
            I => \N__38327\
        );

    \I__6877\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38327\
        );

    \I__6876\ : InMux
    port map (
            O => \N__38358\,
            I => \N__38327\
        );

    \I__6875\ : InMux
    port map (
            O => \N__38357\,
            I => \N__38327\
        );

    \I__6874\ : InMux
    port map (
            O => \N__38356\,
            I => \N__38324\
        );

    \I__6873\ : Odrv12
    port map (
            O => \N__38353\,
            I => count_enable_adj_4544
        );

    \I__6872\ : Odrv4
    port map (
            O => \N__38348\,
            I => count_enable_adj_4544
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__38343\,
            I => count_enable_adj_4544
        );

    \I__6870\ : Odrv12
    port map (
            O => \N__38336\,
            I => count_enable_adj_4544
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__38327\,
            I => count_enable_adj_4544
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__38324\,
            I => count_enable_adj_4544
        );

    \I__6867\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38308\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__38308\,
            I => \N__38305\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__38305\,
            I => \N__38302\
        );

    \I__6864\ : Span4Mux_h
    port map (
            O => \N__38302\,
            I => \N__38299\
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__38299\,
            I => n2185
        );

    \I__6862\ : InMux
    port map (
            O => \N__38296\,
            I => \N__38291\
        );

    \I__6861\ : InMux
    port map (
            O => \N__38295\,
            I => \N__38288\
        );

    \I__6860\ : InMux
    port map (
            O => \N__38294\,
            I => \N__38285\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__38291\,
            I => \N__38282\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__38288\,
            I => \N__38279\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__38285\,
            I => \N__38276\
        );

    \I__6856\ : Span4Mux_v
    port map (
            O => \N__38282\,
            I => \N__38273\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__38279\,
            I => \N__38270\
        );

    \I__6854\ : Span4Mux_h
    port map (
            O => \N__38276\,
            I => \N__38267\
        );

    \I__6853\ : Sp12to4
    port map (
            O => \N__38273\,
            I => \N__38264\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__38270\,
            I => \c0.n13839\
        );

    \I__6851\ : Odrv4
    port map (
            O => \N__38267\,
            I => \c0.n13839\
        );

    \I__6850\ : Odrv12
    port map (
            O => \N__38264\,
            I => \c0.n13839\
        );

    \I__6849\ : InMux
    port map (
            O => \N__38257\,
            I => \N__38254\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__38254\,
            I => \N__38251\
        );

    \I__6847\ : Odrv4
    port map (
            O => \N__38251\,
            I => \c0.n22015\
        );

    \I__6846\ : CascadeMux
    port map (
            O => \N__38248\,
            I => \N__38239\
        );

    \I__6845\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38236\
        );

    \I__6844\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38233\
        );

    \I__6843\ : CascadeMux
    port map (
            O => \N__38245\,
            I => \N__38230\
        );

    \I__6842\ : InMux
    port map (
            O => \N__38244\,
            I => \N__38227\
        );

    \I__6841\ : InMux
    port map (
            O => \N__38243\,
            I => \N__38222\
        );

    \I__6840\ : InMux
    port map (
            O => \N__38242\,
            I => \N__38222\
        );

    \I__6839\ : InMux
    port map (
            O => \N__38239\,
            I => \N__38218\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__38236\,
            I => \N__38215\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__38233\,
            I => \N__38212\
        );

    \I__6836\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38209\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__38227\,
            I => \N__38204\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__38222\,
            I => \N__38204\
        );

    \I__6833\ : InMux
    port map (
            O => \N__38221\,
            I => \N__38201\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__38218\,
            I => \N__38196\
        );

    \I__6831\ : Span4Mux_v
    port map (
            O => \N__38215\,
            I => \N__38196\
        );

    \I__6830\ : Span4Mux_h
    port map (
            O => \N__38212\,
            I => \N__38193\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__38209\,
            I => \N__38188\
        );

    \I__6828\ : Span4Mux_h
    port map (
            O => \N__38204\,
            I => \N__38188\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__38201\,
            I => encoder0_position_29
        );

    \I__6826\ : Odrv4
    port map (
            O => \N__38196\,
            I => encoder0_position_29
        );

    \I__6825\ : Odrv4
    port map (
            O => \N__38193\,
            I => encoder0_position_29
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__38188\,
            I => encoder0_position_29
        );

    \I__6823\ : InMux
    port map (
            O => \N__38179\,
            I => \N__38176\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__38176\,
            I => \N__38173\
        );

    \I__6821\ : Span4Mux_h
    port map (
            O => \N__38173\,
            I => \N__38170\
        );

    \I__6820\ : Odrv4
    port map (
            O => \N__38170\,
            I => \c0.data_out_frame_29__7__N_856\
        );

    \I__6819\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38164\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__38164\,
            I => \N__38160\
        );

    \I__6817\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38157\
        );

    \I__6816\ : Span4Mux_h
    port map (
            O => \N__38160\,
            I => \N__38154\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__38157\,
            I => \c0.n22382\
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__38154\,
            I => \c0.n22382\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__38149\,
            I => \N__38146\
        );

    \I__6812\ : InMux
    port map (
            O => \N__38146\,
            I => \N__38143\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__38143\,
            I => \N__38140\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__38140\,
            I => \c0.n6_adj_4311\
        );

    \I__6809\ : InMux
    port map (
            O => \N__38137\,
            I => \N__38134\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__38134\,
            I => \c0.n14_adj_4400\
        );

    \I__6807\ : CascadeMux
    port map (
            O => \N__38131\,
            I => \c0.n17600_cascade_\
        );

    \I__6806\ : InMux
    port map (
            O => \N__38128\,
            I => \N__38122\
        );

    \I__6805\ : InMux
    port map (
            O => \N__38127\,
            I => \N__38122\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__38122\,
            I => \c0.data_in_frame_10_4\
        );

    \I__6803\ : SRMux
    port map (
            O => \N__38119\,
            I => \N__38116\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__38116\,
            I => \N__38113\
        );

    \I__6801\ : Odrv12
    port map (
            O => \N__38113\,
            I => \c0.n21342\
        );

    \I__6800\ : InMux
    port map (
            O => \N__38110\,
            I => \N__38104\
        );

    \I__6799\ : InMux
    port map (
            O => \N__38109\,
            I => \N__38101\
        );

    \I__6798\ : InMux
    port map (
            O => \N__38108\,
            I => \N__38098\
        );

    \I__6797\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38095\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__38104\,
            I => \N__38088\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__38101\,
            I => \N__38088\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__38098\,
            I => \N__38088\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__38095\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__6792\ : Odrv12
    port map (
            O => \N__38088\,
            I => \c0.FRAME_MATCHER_state_11\
        );

    \I__6791\ : SRMux
    port map (
            O => \N__38083\,
            I => \N__38080\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__38080\,
            I => \N__38077\
        );

    \I__6789\ : Span4Mux_h
    port map (
            O => \N__38077\,
            I => \N__38074\
        );

    \I__6788\ : Odrv4
    port map (
            O => \N__38074\,
            I => \c0.n21350\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__38071\,
            I => \N__38067\
        );

    \I__6786\ : CascadeMux
    port map (
            O => \N__38070\,
            I => \N__38064\
        );

    \I__6785\ : InMux
    port map (
            O => \N__38067\,
            I => \N__38060\
        );

    \I__6784\ : InMux
    port map (
            O => \N__38064\,
            I => \N__38056\
        );

    \I__6783\ : InMux
    port map (
            O => \N__38063\,
            I => \N__38053\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__38060\,
            I => \N__38050\
        );

    \I__6781\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38047\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__38056\,
            I => \N__38043\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__38053\,
            I => \N__38040\
        );

    \I__6778\ : Span4Mux_v
    port map (
            O => \N__38050\,
            I => \N__38035\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__38047\,
            I => \N__38035\
        );

    \I__6776\ : InMux
    port map (
            O => \N__38046\,
            I => \N__38032\
        );

    \I__6775\ : Span4Mux_h
    port map (
            O => \N__38043\,
            I => \N__38025\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__38040\,
            I => \N__38025\
        );

    \I__6773\ : Span4Mux_v
    port map (
            O => \N__38035\,
            I => \N__38025\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__38032\,
            I => encoder1_position_13
        );

    \I__6771\ : Odrv4
    port map (
            O => \N__38025\,
            I => encoder1_position_13
        );

    \I__6770\ : InMux
    port map (
            O => \N__38020\,
            I => \N__38017\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__38017\,
            I => \N__38014\
        );

    \I__6768\ : Span4Mux_v
    port map (
            O => \N__38014\,
            I => \N__38011\
        );

    \I__6767\ : Span4Mux_h
    port map (
            O => \N__38011\,
            I => \N__38008\
        );

    \I__6766\ : Span4Mux_h
    port map (
            O => \N__38008\,
            I => \N__38004\
        );

    \I__6765\ : InMux
    port map (
            O => \N__38007\,
            I => \N__38001\
        );

    \I__6764\ : Span4Mux_v
    port map (
            O => \N__38004\,
            I => \N__37998\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__38001\,
            I => data_out_frame_12_5
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__37998\,
            I => data_out_frame_12_5
        );

    \I__6761\ : InMux
    port map (
            O => \N__37993\,
            I => \N__37990\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__37990\,
            I => \N__37987\
        );

    \I__6759\ : Odrv4
    port map (
            O => \N__37987\,
            I => \c0.n14_adj_4364\
        );

    \I__6758\ : InMux
    port map (
            O => \N__37984\,
            I => \N__37981\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__37981\,
            I => \c0.n13\
        );

    \I__6756\ : CascadeMux
    port map (
            O => \N__37978\,
            I => \c0.n13_adj_4366_cascade_\
        );

    \I__6755\ : InMux
    port map (
            O => \N__37975\,
            I => \N__37972\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__37972\,
            I => \c0.n14_adj_4365\
        );

    \I__6753\ : InMux
    port map (
            O => \N__37969\,
            I => \N__37966\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__37966\,
            I => \N__37963\
        );

    \I__6751\ : Span4Mux_v
    port map (
            O => \N__37963\,
            I => \N__37960\
        );

    \I__6750\ : Odrv4
    port map (
            O => \N__37960\,
            I => \c0.n20_adj_4482\
        );

    \I__6749\ : CascadeMux
    port map (
            O => \N__37957\,
            I => \c0.n21_adj_4480_cascade_\
        );

    \I__6748\ : InMux
    port map (
            O => \N__37954\,
            I => \N__37951\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__37951\,
            I => \N__37948\
        );

    \I__6746\ : Odrv4
    port map (
            O => \N__37948\,
            I => \c0.n19_adj_4481\
        );

    \I__6745\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37941\
        );

    \I__6744\ : CascadeMux
    port map (
            O => \N__37944\,
            I => \N__37937\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__37941\,
            I => \N__37934\
        );

    \I__6742\ : InMux
    port map (
            O => \N__37940\,
            I => \N__37931\
        );

    \I__6741\ : InMux
    port map (
            O => \N__37937\,
            I => \N__37928\
        );

    \I__6740\ : Span12Mux_h
    port map (
            O => \N__37934\,
            I => \N__37921\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__37931\,
            I => \N__37921\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__37928\,
            I => \N__37921\
        );

    \I__6737\ : Odrv12
    port map (
            O => \N__37921\,
            I => \c0.n14789\
        );

    \I__6736\ : CascadeMux
    port map (
            O => \N__37918\,
            I => \N__37915\
        );

    \I__6735\ : InMux
    port map (
            O => \N__37915\,
            I => \N__37910\
        );

    \I__6734\ : InMux
    port map (
            O => \N__37914\,
            I => \N__37907\
        );

    \I__6733\ : InMux
    port map (
            O => \N__37913\,
            I => \N__37904\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__37910\,
            I => \N__37896\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__37907\,
            I => \N__37896\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__37904\,
            I => \N__37896\
        );

    \I__6729\ : InMux
    port map (
            O => \N__37903\,
            I => \N__37893\
        );

    \I__6728\ : Span4Mux_v
    port map (
            O => \N__37896\,
            I => \N__37890\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__37893\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__37890\,
            I => \c0.FRAME_MATCHER_state_18\
        );

    \I__6725\ : CascadeMux
    port map (
            O => \N__37885\,
            I => \N__37882\
        );

    \I__6724\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37877\
        );

    \I__6723\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37873\
        );

    \I__6722\ : InMux
    port map (
            O => \N__37880\,
            I => \N__37870\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__37877\,
            I => \N__37867\
        );

    \I__6720\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37864\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__37873\,
            I => \N__37857\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__37870\,
            I => \N__37857\
        );

    \I__6717\ : Span4Mux_v
    port map (
            O => \N__37867\,
            I => \N__37857\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__37864\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__37857\,
            I => \c0.FRAME_MATCHER_state_16\
        );

    \I__6714\ : InMux
    port map (
            O => \N__37852\,
            I => \N__37849\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__37849\,
            I => \N__37843\
        );

    \I__6712\ : InMux
    port map (
            O => \N__37848\,
            I => \N__37840\
        );

    \I__6711\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37837\
        );

    \I__6710\ : InMux
    port map (
            O => \N__37846\,
            I => \N__37834\
        );

    \I__6709\ : Span4Mux_h
    port map (
            O => \N__37843\,
            I => \N__37831\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__37840\,
            I => \N__37828\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__37837\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__37834\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__6705\ : Odrv4
    port map (
            O => \N__37831\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__6704\ : Odrv4
    port map (
            O => \N__37828\,
            I => \c0.FRAME_MATCHER_state_17\
        );

    \I__6703\ : InMux
    port map (
            O => \N__37819\,
            I => \N__37815\
        );

    \I__6702\ : InMux
    port map (
            O => \N__37818\,
            I => \N__37812\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__37815\,
            I => \N__37807\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__37812\,
            I => \N__37807\
        );

    \I__6699\ : Odrv4
    port map (
            O => \N__37807\,
            I => \c0.n21682\
        );

    \I__6698\ : InMux
    port map (
            O => \N__37804\,
            I => \N__37800\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__37803\,
            I => \N__37796\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__37800\,
            I => \N__37793\
        );

    \I__6695\ : InMux
    port map (
            O => \N__37799\,
            I => \N__37790\
        );

    \I__6694\ : InMux
    port map (
            O => \N__37796\,
            I => \N__37786\
        );

    \I__6693\ : Span4Mux_h
    port map (
            O => \N__37793\,
            I => \N__37783\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__37790\,
            I => \N__37780\
        );

    \I__6691\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37777\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__37786\,
            I => \N__37774\
        );

    \I__6689\ : Span4Mux_h
    port map (
            O => \N__37783\,
            I => \N__37769\
        );

    \I__6688\ : Span4Mux_h
    port map (
            O => \N__37780\,
            I => \N__37769\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__37777\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__6686\ : Odrv12
    port map (
            O => \N__37774\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__6685\ : Odrv4
    port map (
            O => \N__37769\,
            I => \c0.FRAME_MATCHER_state_4\
        );

    \I__6684\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37759\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__37759\,
            I => \N__37756\
        );

    \I__6682\ : Odrv4
    port map (
            O => \N__37756\,
            I => \c0.n47\
        );

    \I__6681\ : InMux
    port map (
            O => \N__37753\,
            I => \N__37747\
        );

    \I__6680\ : InMux
    port map (
            O => \N__37752\,
            I => \N__37744\
        );

    \I__6679\ : InMux
    port map (
            O => \N__37751\,
            I => \N__37741\
        );

    \I__6678\ : InMux
    port map (
            O => \N__37750\,
            I => \N__37738\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__37747\,
            I => \N__37735\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__37744\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__37741\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__37738\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__6673\ : Odrv4
    port map (
            O => \N__37735\,
            I => \c0.FRAME_MATCHER_state_25\
        );

    \I__6672\ : SRMux
    port map (
            O => \N__37726\,
            I => \N__37723\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__37723\,
            I => \N__37720\
        );

    \I__6670\ : Odrv12
    port map (
            O => \N__37720\,
            I => \c0.n21374\
        );

    \I__6669\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37711\
        );

    \I__6668\ : InMux
    port map (
            O => \N__37716\,
            I => \N__37708\
        );

    \I__6667\ : InMux
    port map (
            O => \N__37715\,
            I => \N__37703\
        );

    \I__6666\ : InMux
    port map (
            O => \N__37714\,
            I => \N__37703\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__37711\,
            I => \N__37698\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__37708\,
            I => \N__37698\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__37703\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__37698\,
            I => \c0.FRAME_MATCHER_state_10\
        );

    \I__6661\ : SRMux
    port map (
            O => \N__37693\,
            I => \N__37690\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__37690\,
            I => \c0.n21348\
        );

    \I__6659\ : InMux
    port map (
            O => \N__37687\,
            I => \N__37681\
        );

    \I__6658\ : InMux
    port map (
            O => \N__37686\,
            I => \N__37676\
        );

    \I__6657\ : InMux
    port map (
            O => \N__37685\,
            I => \N__37676\
        );

    \I__6656\ : InMux
    port map (
            O => \N__37684\,
            I => \N__37673\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__37681\,
            I => \N__37668\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__37676\,
            I => \N__37668\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__37673\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__6652\ : Odrv4
    port map (
            O => \N__37668\,
            I => \c0.FRAME_MATCHER_state_7\
        );

    \I__6651\ : CascadeMux
    port map (
            O => \N__37663\,
            I => \c0.n48_cascade_\
        );

    \I__6650\ : InMux
    port map (
            O => \N__37660\,
            I => \N__37657\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__37657\,
            I => \c0.n45_adj_4413\
        );

    \I__6648\ : CascadeMux
    port map (
            O => \N__37654\,
            I => \N__37650\
        );

    \I__6647\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37645\
        );

    \I__6646\ : InMux
    port map (
            O => \N__37650\,
            I => \N__37645\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__37645\,
            I => \N__37642\
        );

    \I__6644\ : Span4Mux_v
    port map (
            O => \N__37642\,
            I => \N__37637\
        );

    \I__6643\ : InMux
    port map (
            O => \N__37641\,
            I => \N__37634\
        );

    \I__6642\ : InMux
    port map (
            O => \N__37640\,
            I => \N__37631\
        );

    \I__6641\ : Sp12to4
    port map (
            O => \N__37637\,
            I => \N__37628\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__37634\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__37631\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__6638\ : Odrv12
    port map (
            O => \N__37628\,
            I => \c0.FRAME_MATCHER_state_23\
        );

    \I__6637\ : InMux
    port map (
            O => \N__37621\,
            I => \N__37617\
        );

    \I__6636\ : InMux
    port map (
            O => \N__37620\,
            I => \N__37614\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__37617\,
            I => \c0.n14_adj_4316\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__37614\,
            I => \c0.n14_adj_4316\
        );

    \I__6633\ : InMux
    port map (
            O => \N__37609\,
            I => \N__37606\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__37606\,
            I => \N__37600\
        );

    \I__6631\ : InMux
    port map (
            O => \N__37605\,
            I => \N__37593\
        );

    \I__6630\ : InMux
    port map (
            O => \N__37604\,
            I => \N__37593\
        );

    \I__6629\ : InMux
    port map (
            O => \N__37603\,
            I => \N__37593\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__37600\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__37593\,
            I => \c0.FRAME_MATCHER_state_24\
        );

    \I__6626\ : SRMux
    port map (
            O => \N__37588\,
            I => \N__37585\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__37585\,
            I => \c0.n21372\
        );

    \I__6624\ : SRMux
    port map (
            O => \N__37582\,
            I => \N__37579\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__37579\,
            I => \N__37576\
        );

    \I__6622\ : Span4Mux_h
    port map (
            O => \N__37576\,
            I => \N__37573\
        );

    \I__6621\ : Odrv4
    port map (
            O => \N__37573\,
            I => \c0.n21346\
        );

    \I__6620\ : SRMux
    port map (
            O => \N__37570\,
            I => \N__37567\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__37567\,
            I => \N__37564\
        );

    \I__6618\ : Span4Mux_v
    port map (
            O => \N__37564\,
            I => \N__37561\
        );

    \I__6617\ : Span4Mux_h
    port map (
            O => \N__37561\,
            I => \N__37558\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__37558\,
            I => \c0.n21364\
        );

    \I__6615\ : CascadeMux
    port map (
            O => \N__37555\,
            I => \N__37552\
        );

    \I__6614\ : InMux
    port map (
            O => \N__37552\,
            I => \N__37546\
        );

    \I__6613\ : InMux
    port map (
            O => \N__37551\,
            I => \N__37546\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__37546\,
            I => \N__37542\
        );

    \I__6611\ : InMux
    port map (
            O => \N__37545\,
            I => \N__37538\
        );

    \I__6610\ : Span4Mux_v
    port map (
            O => \N__37542\,
            I => \N__37535\
        );

    \I__6609\ : InMux
    port map (
            O => \N__37541\,
            I => \N__37532\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__37538\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__6607\ : Odrv4
    port map (
            O => \N__37535\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__37532\,
            I => \c0.FRAME_MATCHER_state_9\
        );

    \I__6605\ : InMux
    port map (
            O => \N__37525\,
            I => \N__37522\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__37522\,
            I => \c0.n46\
        );

    \I__6603\ : CascadeMux
    port map (
            O => \N__37519\,
            I => \N__37516\
        );

    \I__6602\ : InMux
    port map (
            O => \N__37516\,
            I => \N__37510\
        );

    \I__6601\ : InMux
    port map (
            O => \N__37515\,
            I => \N__37503\
        );

    \I__6600\ : InMux
    port map (
            O => \N__37514\,
            I => \N__37503\
        );

    \I__6599\ : InMux
    port map (
            O => \N__37513\,
            I => \N__37503\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__37510\,
            I => \N__37496\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__37503\,
            I => \N__37496\
        );

    \I__6596\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37489\
        );

    \I__6595\ : InMux
    port map (
            O => \N__37501\,
            I => \N__37489\
        );

    \I__6594\ : Span4Mux_h
    port map (
            O => \N__37496\,
            I => \N__37486\
        );

    \I__6593\ : InMux
    port map (
            O => \N__37495\,
            I => \N__37481\
        );

    \I__6592\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37481\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__37489\,
            I => \c0.n117\
        );

    \I__6590\ : Odrv4
    port map (
            O => \N__37486\,
            I => \c0.n117\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__37481\,
            I => \c0.n117\
        );

    \I__6588\ : InMux
    port map (
            O => \N__37474\,
            I => \N__37459\
        );

    \I__6587\ : InMux
    port map (
            O => \N__37473\,
            I => \N__37459\
        );

    \I__6586\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37459\
        );

    \I__6585\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37459\
        );

    \I__6584\ : InMux
    port map (
            O => \N__37470\,
            I => \N__37454\
        );

    \I__6583\ : InMux
    port map (
            O => \N__37469\,
            I => \N__37454\
        );

    \I__6582\ : InMux
    port map (
            O => \N__37468\,
            I => \N__37451\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__37459\,
            I => \N__37446\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__37454\,
            I => \N__37446\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__37451\,
            I => \N__37443\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__37446\,
            I => \N__37440\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__37443\,
            I => \c0.n63_adj_4301\
        );

    \I__6576\ : Odrv4
    port map (
            O => \N__37440\,
            I => \c0.n63_adj_4301\
        );

    \I__6575\ : CascadeMux
    port map (
            O => \N__37435\,
            I => \c0.n16958_cascade_\
        );

    \I__6574\ : CascadeMux
    port map (
            O => \N__37432\,
            I => \N__37425\
        );

    \I__6573\ : InMux
    port map (
            O => \N__37431\,
            I => \N__37415\
        );

    \I__6572\ : InMux
    port map (
            O => \N__37430\,
            I => \N__37415\
        );

    \I__6571\ : InMux
    port map (
            O => \N__37429\,
            I => \N__37415\
        );

    \I__6570\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37415\
        );

    \I__6569\ : InMux
    port map (
            O => \N__37425\,
            I => \N__37410\
        );

    \I__6568\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37410\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__37415\,
            I => \N__37404\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__37410\,
            I => \N__37404\
        );

    \I__6565\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37401\
        );

    \I__6564\ : Span4Mux_h
    port map (
            O => \N__37404\,
            I => \N__37398\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__37401\,
            I => \c0.n63\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__37398\,
            I => \c0.n63\
        );

    \I__6561\ : CascadeMux
    port map (
            O => \N__37393\,
            I => \c0.n22695_cascade_\
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__37390\,
            I => \N__37385\
        );

    \I__6559\ : InMux
    port map (
            O => \N__37389\,
            I => \N__37382\
        );

    \I__6558\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37377\
        );

    \I__6557\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37377\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__37382\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__37377\,
            I => \c0.FRAME_MATCHER_state_2\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__37372\,
            I => \N__37369\
        );

    \I__6553\ : InMux
    port map (
            O => \N__37369\,
            I => \N__37366\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__37366\,
            I => \N__37363\
        );

    \I__6551\ : Odrv4
    port map (
            O => \N__37363\,
            I => \c0.n13_adj_4388\
        );

    \I__6550\ : InMux
    port map (
            O => \N__37360\,
            I => \N__37357\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__37357\,
            I => \N__37353\
        );

    \I__6548\ : InMux
    port map (
            O => \N__37356\,
            I => \N__37350\
        );

    \I__6547\ : Odrv4
    port map (
            O => \N__37353\,
            I => \c0.n9207\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__37350\,
            I => \c0.n9207\
        );

    \I__6545\ : InMux
    port map (
            O => \N__37345\,
            I => \N__37342\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__37342\,
            I => \c0.n14_adj_4337\
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__37339\,
            I => \c0.n7_adj_4352_cascade_\
        );

    \I__6542\ : InMux
    port map (
            O => \N__37336\,
            I => \N__37331\
        );

    \I__6541\ : CascadeMux
    port map (
            O => \N__37335\,
            I => \N__37328\
        );

    \I__6540\ : InMux
    port map (
            O => \N__37334\,
            I => \N__37325\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__37331\,
            I => \N__37322\
        );

    \I__6538\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37319\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__37325\,
            I => \N__37313\
        );

    \I__6536\ : Span4Mux_h
    port map (
            O => \N__37322\,
            I => \N__37313\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__37319\,
            I => \N__37310\
        );

    \I__6534\ : InMux
    port map (
            O => \N__37318\,
            I => \N__37307\
        );

    \I__6533\ : Sp12to4
    port map (
            O => \N__37313\,
            I => \N__37302\
        );

    \I__6532\ : Span12Mux_v
    port map (
            O => \N__37310\,
            I => \N__37302\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__37307\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__6530\ : Odrv12
    port map (
            O => \N__37302\,
            I => \c0.FRAME_MATCHER_state_26\
        );

    \I__6529\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37294\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__37294\,
            I => \N__37291\
        );

    \I__6527\ : Odrv4
    port map (
            O => \N__37291\,
            I => \c0.n21789\
        );

    \I__6526\ : CascadeMux
    port map (
            O => \N__37288\,
            I => \c0.n12996_cascade_\
        );

    \I__6525\ : CascadeMux
    port map (
            O => \N__37285\,
            I => \c0.n13020_cascade_\
        );

    \I__6524\ : CascadeMux
    port map (
            O => \N__37282\,
            I => \c0.data_out_frame_29_7_N_1483_1_cascade_\
        );

    \I__6523\ : InMux
    port map (
            O => \N__37279\,
            I => \N__37276\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__37276\,
            I => \c0.n6650\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__37273\,
            I => \c0.n6650_cascade_\
        );

    \I__6520\ : InMux
    port map (
            O => \N__37270\,
            I => \N__37267\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__37267\,
            I => \c0.n6_adj_4270\
        );

    \I__6518\ : CascadeMux
    port map (
            O => \N__37264\,
            I => \N__37260\
        );

    \I__6517\ : InMux
    port map (
            O => \N__37263\,
            I => \N__37257\
        );

    \I__6516\ : InMux
    port map (
            O => \N__37260\,
            I => \N__37254\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__37257\,
            I => \N__37251\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__37254\,
            I => \N__37247\
        );

    \I__6513\ : Span4Mux_h
    port map (
            O => \N__37251\,
            I => \N__37243\
        );

    \I__6512\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37240\
        );

    \I__6511\ : Span4Mux_h
    port map (
            O => \N__37247\,
            I => \N__37237\
        );

    \I__6510\ : InMux
    port map (
            O => \N__37246\,
            I => \N__37234\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__37243\,
            I => \N__37231\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__37240\,
            I => encoder1_position_17
        );

    \I__6507\ : Odrv4
    port map (
            O => \N__37237\,
            I => encoder1_position_17
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__37234\,
            I => encoder1_position_17
        );

    \I__6505\ : Odrv4
    port map (
            O => \N__37231\,
            I => encoder1_position_17
        );

    \I__6504\ : CascadeMux
    port map (
            O => \N__37222\,
            I => \N__37218\
        );

    \I__6503\ : InMux
    port map (
            O => \N__37221\,
            I => \N__37215\
        );

    \I__6502\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37212\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__37215\,
            I => data_out_frame_11_1
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__37212\,
            I => data_out_frame_11_1
        );

    \I__6499\ : CascadeMux
    port map (
            O => \N__37207\,
            I => \c0.n9_adj_4415_cascade_\
        );

    \I__6498\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37200\
        );

    \I__6497\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37197\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__37200\,
            I => \N__37194\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__37197\,
            I => \N__37190\
        );

    \I__6494\ : Span4Mux_v
    port map (
            O => \N__37194\,
            I => \N__37187\
        );

    \I__6493\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37184\
        );

    \I__6492\ : Span12Mux_h
    port map (
            O => \N__37190\,
            I => \N__37181\
        );

    \I__6491\ : Sp12to4
    port map (
            O => \N__37187\,
            I => \N__37176\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__37184\,
            I => \N__37176\
        );

    \I__6489\ : Odrv12
    port map (
            O => \N__37181\,
            I => n14252
        );

    \I__6488\ : Odrv12
    port map (
            O => \N__37176\,
            I => n14252
        );

    \I__6487\ : InMux
    port map (
            O => \N__37171\,
            I => \N__37167\
        );

    \I__6486\ : InMux
    port map (
            O => \N__37170\,
            I => \N__37164\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__37167\,
            I => \N__37161\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__37164\,
            I => \N__37158\
        );

    \I__6483\ : Span4Mux_h
    port map (
            O => \N__37161\,
            I => \N__37155\
        );

    \I__6482\ : Span4Mux_v
    port map (
            O => \N__37158\,
            I => \N__37152\
        );

    \I__6481\ : Odrv4
    port map (
            O => \N__37155\,
            I => \c0.n38_adj_4387\
        );

    \I__6480\ : Odrv4
    port map (
            O => \N__37152\,
            I => \c0.n38_adj_4387\
        );

    \I__6479\ : InMux
    port map (
            O => \N__37147\,
            I => \N__37143\
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__37146\,
            I => \N__37139\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__37143\,
            I => \N__37136\
        );

    \I__6476\ : InMux
    port map (
            O => \N__37142\,
            I => \N__37132\
        );

    \I__6475\ : InMux
    port map (
            O => \N__37139\,
            I => \N__37129\
        );

    \I__6474\ : Span4Mux_h
    port map (
            O => \N__37136\,
            I => \N__37126\
        );

    \I__6473\ : InMux
    port map (
            O => \N__37135\,
            I => \N__37123\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__37132\,
            I => \N__37118\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__37129\,
            I => \N__37118\
        );

    \I__6470\ : Odrv4
    port map (
            O => \N__37126\,
            I => \c0.tx_active\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__37123\,
            I => \c0.tx_active\
        );

    \I__6468\ : Odrv12
    port map (
            O => \N__37118\,
            I => \c0.tx_active\
        );

    \I__6467\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37108\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__37108\,
            I => \c0.n22651\
        );

    \I__6465\ : CascadeMux
    port map (
            O => \N__37105\,
            I => \n22661_cascade_\
        );

    \I__6464\ : InMux
    port map (
            O => \N__37102\,
            I => \N__37099\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__37099\,
            I => \N__37095\
        );

    \I__6462\ : InMux
    port map (
            O => \N__37098\,
            I => \N__37092\
        );

    \I__6461\ : Span4Mux_h
    port map (
            O => \N__37095\,
            I => \N__37089\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__37092\,
            I => data_out_frame_7_3
        );

    \I__6459\ : Odrv4
    port map (
            O => \N__37089\,
            I => data_out_frame_7_3
        );

    \I__6458\ : InMux
    port map (
            O => \N__37084\,
            I => \N__37080\
        );

    \I__6457\ : InMux
    port map (
            O => \N__37083\,
            I => \N__37077\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__37080\,
            I => data_out_frame_6_1
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__37077\,
            I => data_out_frame_6_1
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__37072\,
            I => \N__37068\
        );

    \I__6453\ : CascadeMux
    port map (
            O => \N__37071\,
            I => \N__37065\
        );

    \I__6452\ : InMux
    port map (
            O => \N__37068\,
            I => \N__37062\
        );

    \I__6451\ : InMux
    port map (
            O => \N__37065\,
            I => \N__37057\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__37062\,
            I => \N__37054\
        );

    \I__6449\ : InMux
    port map (
            O => \N__37061\,
            I => \N__37051\
        );

    \I__6448\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37048\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__37057\,
            I => \N__37043\
        );

    \I__6446\ : Span4Mux_v
    port map (
            O => \N__37054\,
            I => \N__37036\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__37051\,
            I => \N__37036\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__37048\,
            I => \N__37036\
        );

    \I__6443\ : InMux
    port map (
            O => \N__37047\,
            I => \N__37033\
        );

    \I__6442\ : InMux
    port map (
            O => \N__37046\,
            I => \N__37030\
        );

    \I__6441\ : Span4Mux_v
    port map (
            O => \N__37043\,
            I => \N__37025\
        );

    \I__6440\ : Span4Mux_h
    port map (
            O => \N__37036\,
            I => \N__37025\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__37033\,
            I => encoder0_position_0
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__37030\,
            I => encoder0_position_0
        );

    \I__6437\ : Odrv4
    port map (
            O => \N__37025\,
            I => encoder0_position_0
        );

    \I__6436\ : InMux
    port map (
            O => \N__37018\,
            I => \N__37015\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__37015\,
            I => \N__37011\
        );

    \I__6434\ : InMux
    port map (
            O => \N__37014\,
            I => \N__37008\
        );

    \I__6433\ : Span4Mux_v
    port map (
            O => \N__37011\,
            I => \N__37005\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__37008\,
            I => data_out_frame_9_0
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__37005\,
            I => data_out_frame_9_0
        );

    \I__6430\ : InMux
    port map (
            O => \N__37000\,
            I => \N__36997\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__36997\,
            I => n2242
        );

    \I__6428\ : InMux
    port map (
            O => \N__36994\,
            I => \N__36990\
        );

    \I__6427\ : InMux
    port map (
            O => \N__36993\,
            I => \N__36987\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__36990\,
            I => \N__36982\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__36987\,
            I => \N__36979\
        );

    \I__6424\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36974\
        );

    \I__6423\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36974\
        );

    \I__6422\ : Span12Mux_v
    port map (
            O => \N__36982\,
            I => \N__36971\
        );

    \I__6421\ : Span4Mux_v
    port map (
            O => \N__36979\,
            I => \N__36968\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__36974\,
            I => data_in_3_6
        );

    \I__6419\ : Odrv12
    port map (
            O => \N__36971\,
            I => data_in_3_6
        );

    \I__6418\ : Odrv4
    port map (
            O => \N__36968\,
            I => data_in_3_6
        );

    \I__6417\ : CascadeMux
    port map (
            O => \N__36961\,
            I => \N__36957\
        );

    \I__6416\ : InMux
    port map (
            O => \N__36960\,
            I => \N__36952\
        );

    \I__6415\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36952\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__36952\,
            I => \N__36949\
        );

    \I__6413\ : Span4Mux_h
    port map (
            O => \N__36949\,
            I => \N__36944\
        );

    \I__6412\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36941\
        );

    \I__6411\ : InMux
    port map (
            O => \N__36947\,
            I => \N__36938\
        );

    \I__6410\ : Span4Mux_v
    port map (
            O => \N__36944\,
            I => \N__36933\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__36941\,
            I => \N__36933\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__36938\,
            I => data_in_2_6
        );

    \I__6407\ : Odrv4
    port map (
            O => \N__36933\,
            I => data_in_2_6
        );

    \I__6406\ : InMux
    port map (
            O => \N__36928\,
            I => \N__36925\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__36925\,
            I => \N__36921\
        );

    \I__6404\ : InMux
    port map (
            O => \N__36924\,
            I => \N__36918\
        );

    \I__6403\ : Span12Mux_v
    port map (
            O => \N__36921\,
            I => \N__36915\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__36918\,
            I => data_out_frame_10_1
        );

    \I__6401\ : Odrv12
    port map (
            O => \N__36915\,
            I => data_out_frame_10_1
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__36910\,
            I => \N__36903\
        );

    \I__6399\ : InMux
    port map (
            O => \N__36909\,
            I => \N__36891\
        );

    \I__6398\ : InMux
    port map (
            O => \N__36908\,
            I => \N__36884\
        );

    \I__6397\ : InMux
    port map (
            O => \N__36907\,
            I => \N__36877\
        );

    \I__6396\ : InMux
    port map (
            O => \N__36906\,
            I => \N__36877\
        );

    \I__6395\ : InMux
    port map (
            O => \N__36903\,
            I => \N__36874\
        );

    \I__6394\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36867\
        );

    \I__6393\ : CascadeMux
    port map (
            O => \N__36901\,
            I => \N__36864\
        );

    \I__6392\ : CascadeMux
    port map (
            O => \N__36900\,
            I => \N__36859\
        );

    \I__6391\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36854\
        );

    \I__6390\ : InMux
    port map (
            O => \N__36898\,
            I => \N__36854\
        );

    \I__6389\ : InMux
    port map (
            O => \N__36897\,
            I => \N__36849\
        );

    \I__6388\ : InMux
    port map (
            O => \N__36896\,
            I => \N__36849\
        );

    \I__6387\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36844\
        );

    \I__6386\ : InMux
    port map (
            O => \N__36894\,
            I => \N__36841\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__36891\,
            I => \N__36838\
        );

    \I__6384\ : InMux
    port map (
            O => \N__36890\,
            I => \N__36835\
        );

    \I__6383\ : InMux
    port map (
            O => \N__36889\,
            I => \N__36830\
        );

    \I__6382\ : InMux
    port map (
            O => \N__36888\,
            I => \N__36825\
        );

    \I__6381\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36825\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__36884\,
            I => \N__36822\
        );

    \I__6379\ : InMux
    port map (
            O => \N__36883\,
            I => \N__36819\
        );

    \I__6378\ : InMux
    port map (
            O => \N__36882\,
            I => \N__36814\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__36877\,
            I => \N__36809\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__36874\,
            I => \N__36809\
        );

    \I__6375\ : InMux
    port map (
            O => \N__36873\,
            I => \N__36800\
        );

    \I__6374\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36800\
        );

    \I__6373\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36800\
        );

    \I__6372\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36800\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__36867\,
            I => \N__36797\
        );

    \I__6370\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36788\
        );

    \I__6369\ : InMux
    port map (
            O => \N__36863\,
            I => \N__36788\
        );

    \I__6368\ : InMux
    port map (
            O => \N__36862\,
            I => \N__36788\
        );

    \I__6367\ : InMux
    port map (
            O => \N__36859\,
            I => \N__36788\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__36854\,
            I => \N__36783\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__36849\,
            I => \N__36783\
        );

    \I__6364\ : InMux
    port map (
            O => \N__36848\,
            I => \N__36778\
        );

    \I__6363\ : InMux
    port map (
            O => \N__36847\,
            I => \N__36778\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__36844\,
            I => \N__36769\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__36841\,
            I => \N__36769\
        );

    \I__6360\ : Span4Mux_v
    port map (
            O => \N__36838\,
            I => \N__36769\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__36835\,
            I => \N__36769\
        );

    \I__6358\ : InMux
    port map (
            O => \N__36834\,
            I => \N__36766\
        );

    \I__6357\ : CascadeMux
    port map (
            O => \N__36833\,
            I => \N__36762\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__36830\,
            I => \N__36756\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__36825\,
            I => \N__36749\
        );

    \I__6354\ : Span4Mux_v
    port map (
            O => \N__36822\,
            I => \N__36749\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__36819\,
            I => \N__36749\
        );

    \I__6352\ : InMux
    port map (
            O => \N__36818\,
            I => \N__36746\
        );

    \I__6351\ : CascadeMux
    port map (
            O => \N__36817\,
            I => \N__36743\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__36814\,
            I => \N__36738\
        );

    \I__6349\ : Span4Mux_v
    port map (
            O => \N__36809\,
            I => \N__36733\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__36800\,
            I => \N__36733\
        );

    \I__6347\ : Span4Mux_v
    port map (
            O => \N__36797\,
            I => \N__36728\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__36788\,
            I => \N__36728\
        );

    \I__6345\ : Span4Mux_v
    port map (
            O => \N__36783\,
            I => \N__36721\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__36778\,
            I => \N__36721\
        );

    \I__6343\ : Span4Mux_h
    port map (
            O => \N__36769\,
            I => \N__36721\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__36766\,
            I => \N__36718\
        );

    \I__6341\ : InMux
    port map (
            O => \N__36765\,
            I => \N__36715\
        );

    \I__6340\ : InMux
    port map (
            O => \N__36762\,
            I => \N__36712\
        );

    \I__6339\ : InMux
    port map (
            O => \N__36761\,
            I => \N__36705\
        );

    \I__6338\ : InMux
    port map (
            O => \N__36760\,
            I => \N__36705\
        );

    \I__6337\ : InMux
    port map (
            O => \N__36759\,
            I => \N__36705\
        );

    \I__6336\ : Span4Mux_v
    port map (
            O => \N__36756\,
            I => \N__36698\
        );

    \I__6335\ : Span4Mux_v
    port map (
            O => \N__36749\,
            I => \N__36698\
        );

    \I__6334\ : LocalMux
    port map (
            O => \N__36746\,
            I => \N__36698\
        );

    \I__6333\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36695\
        );

    \I__6332\ : InMux
    port map (
            O => \N__36742\,
            I => \N__36692\
        );

    \I__6331\ : InMux
    port map (
            O => \N__36741\,
            I => \N__36689\
        );

    \I__6330\ : Span4Mux_v
    port map (
            O => \N__36738\,
            I => \N__36682\
        );

    \I__6329\ : Span4Mux_v
    port map (
            O => \N__36733\,
            I => \N__36682\
        );

    \I__6328\ : Span4Mux_v
    port map (
            O => \N__36728\,
            I => \N__36682\
        );

    \I__6327\ : Span4Mux_h
    port map (
            O => \N__36721\,
            I => \N__36679\
        );

    \I__6326\ : Span4Mux_h
    port map (
            O => \N__36718\,
            I => \N__36676\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__36715\,
            I => \N__36665\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__36712\,
            I => \N__36665\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__36705\,
            I => \N__36665\
        );

    \I__6322\ : Sp12to4
    port map (
            O => \N__36698\,
            I => \N__36665\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__36695\,
            I => \N__36665\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__36692\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__36689\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6318\ : Odrv4
    port map (
            O => \N__36682\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6317\ : Odrv4
    port map (
            O => \N__36679\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6316\ : Odrv4
    port map (
            O => \N__36676\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6315\ : Odrv12
    port map (
            O => \N__36665\,
            I => \c0.byte_transmit_counter_1\
        );

    \I__6314\ : InMux
    port map (
            O => \N__36652\,
            I => \N__36649\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__36649\,
            I => \c0.n24183\
        );

    \I__6312\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36638\
        );

    \I__6311\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36638\
        );

    \I__6310\ : InMux
    port map (
            O => \N__36644\,
            I => \N__36633\
        );

    \I__6309\ : InMux
    port map (
            O => \N__36643\,
            I => \N__36633\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__36638\,
            I => \N__36630\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__36633\,
            I => data_in_3_7
        );

    \I__6306\ : Odrv12
    port map (
            O => \N__36630\,
            I => data_in_3_7
        );

    \I__6305\ : InMux
    port map (
            O => \N__36625\,
            I => \N__36620\
        );

    \I__6304\ : InMux
    port map (
            O => \N__36624\,
            I => \N__36617\
        );

    \I__6303\ : InMux
    port map (
            O => \N__36623\,
            I => \N__36614\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__36620\,
            I => \N__36611\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__36617\,
            I => \N__36608\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__36614\,
            I => \N__36605\
        );

    \I__6299\ : Span4Mux_h
    port map (
            O => \N__36611\,
            I => \N__36600\
        );

    \I__6298\ : Span4Mux_v
    port map (
            O => \N__36608\,
            I => \N__36600\
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__36605\,
            I => data_in_2_7
        );

    \I__6296\ : Odrv4
    port map (
            O => \N__36600\,
            I => data_in_2_7
        );

    \I__6295\ : InMux
    port map (
            O => \N__36595\,
            I => \N__36591\
        );

    \I__6294\ : InMux
    port map (
            O => \N__36594\,
            I => \N__36588\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__36591\,
            I => \N__36583\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__36588\,
            I => \N__36580\
        );

    \I__6291\ : InMux
    port map (
            O => \N__36587\,
            I => \N__36577\
        );

    \I__6290\ : InMux
    port map (
            O => \N__36586\,
            I => \N__36574\
        );

    \I__6289\ : Span4Mux_h
    port map (
            O => \N__36583\,
            I => \N__36571\
        );

    \I__6288\ : Span4Mux_v
    port map (
            O => \N__36580\,
            I => \N__36566\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__36577\,
            I => \N__36566\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__36574\,
            I => data_in_3_2
        );

    \I__6285\ : Odrv4
    port map (
            O => \N__36571\,
            I => data_in_3_2
        );

    \I__6284\ : Odrv4
    port map (
            O => \N__36566\,
            I => data_in_3_2
        );

    \I__6283\ : InMux
    port map (
            O => \N__36559\,
            I => \N__36553\
        );

    \I__6282\ : InMux
    port map (
            O => \N__36558\,
            I => \N__36550\
        );

    \I__6281\ : CascadeMux
    port map (
            O => \N__36557\,
            I => \N__36546\
        );

    \I__6280\ : CascadeMux
    port map (
            O => \N__36556\,
            I => \N__36543\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__36553\,
            I => \N__36540\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__36550\,
            I => \N__36537\
        );

    \I__6277\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36532\
        );

    \I__6276\ : InMux
    port map (
            O => \N__36546\,
            I => \N__36532\
        );

    \I__6275\ : InMux
    port map (
            O => \N__36543\,
            I => \N__36527\
        );

    \I__6274\ : Span4Mux_v
    port map (
            O => \N__36540\,
            I => \N__36522\
        );

    \I__6273\ : Span4Mux_h
    port map (
            O => \N__36537\,
            I => \N__36522\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__36532\,
            I => \N__36519\
        );

    \I__6271\ : InMux
    port map (
            O => \N__36531\,
            I => \N__36514\
        );

    \I__6270\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36514\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__36527\,
            I => encoder0_position_17
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__36522\,
            I => encoder0_position_17
        );

    \I__6267\ : Odrv4
    port map (
            O => \N__36519\,
            I => encoder0_position_17
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__36514\,
            I => encoder0_position_17
        );

    \I__6265\ : CascadeMux
    port map (
            O => \N__36505\,
            I => \N__36500\
        );

    \I__6264\ : InMux
    port map (
            O => \N__36504\,
            I => \N__36496\
        );

    \I__6263\ : CascadeMux
    port map (
            O => \N__36503\,
            I => \N__36492\
        );

    \I__6262\ : InMux
    port map (
            O => \N__36500\,
            I => \N__36489\
        );

    \I__6261\ : InMux
    port map (
            O => \N__36499\,
            I => \N__36486\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__36496\,
            I => \N__36483\
        );

    \I__6259\ : InMux
    port map (
            O => \N__36495\,
            I => \N__36480\
        );

    \I__6258\ : InMux
    port map (
            O => \N__36492\,
            I => \N__36477\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__36489\,
            I => \N__36472\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__36486\,
            I => \N__36472\
        );

    \I__6255\ : Span4Mux_h
    port map (
            O => \N__36483\,
            I => \N__36469\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__36480\,
            I => encoder1_position_28
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__36477\,
            I => encoder1_position_28
        );

    \I__6252\ : Odrv12
    port map (
            O => \N__36472\,
            I => encoder1_position_28
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__36469\,
            I => encoder1_position_28
        );

    \I__6250\ : CascadeMux
    port map (
            O => \N__36460\,
            I => \N__36455\
        );

    \I__6249\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36451\
        );

    \I__6248\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36446\
        );

    \I__6247\ : InMux
    port map (
            O => \N__36455\,
            I => \N__36446\
        );

    \I__6246\ : InMux
    port map (
            O => \N__36454\,
            I => \N__36443\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__36451\,
            I => \N__36440\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__36446\,
            I => \N__36433\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__36443\,
            I => \N__36433\
        );

    \I__6242\ : Span4Mux_h
    port map (
            O => \N__36440\,
            I => \N__36433\
        );

    \I__6241\ : Span4Mux_h
    port map (
            O => \N__36433\,
            I => \N__36430\
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__36430\,
            I => \c0.n13338\
        );

    \I__6239\ : InMux
    port map (
            O => \N__36427\,
            I => \N__36422\
        );

    \I__6238\ : InMux
    port map (
            O => \N__36426\,
            I => \N__36419\
        );

    \I__6237\ : CascadeMux
    port map (
            O => \N__36425\,
            I => \N__36416\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__36422\,
            I => \N__36413\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__36419\,
            I => \N__36410\
        );

    \I__6234\ : InMux
    port map (
            O => \N__36416\,
            I => \N__36407\
        );

    \I__6233\ : Span4Mux_h
    port map (
            O => \N__36413\,
            I => \N__36403\
        );

    \I__6232\ : Span4Mux_h
    port map (
            O => \N__36410\,
            I => \N__36398\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__36407\,
            I => \N__36398\
        );

    \I__6230\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36395\
        );

    \I__6229\ : Span4Mux_v
    port map (
            O => \N__36403\,
            I => \N__36392\
        );

    \I__6228\ : Span4Mux_v
    port map (
            O => \N__36398\,
            I => \N__36389\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__36395\,
            I => data_in_2_5
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__36392\,
            I => data_in_2_5
        );

    \I__6225\ : Odrv4
    port map (
            O => \N__36389\,
            I => data_in_2_5
        );

    \I__6224\ : InMux
    port map (
            O => \N__36382\,
            I => \N__36378\
        );

    \I__6223\ : InMux
    port map (
            O => \N__36381\,
            I => \N__36374\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__36378\,
            I => \N__36371\
        );

    \I__6221\ : InMux
    port map (
            O => \N__36377\,
            I => \N__36368\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__36374\,
            I => \N__36364\
        );

    \I__6219\ : Span4Mux_h
    port map (
            O => \N__36371\,
            I => \N__36359\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__36368\,
            I => \N__36359\
        );

    \I__6217\ : InMux
    port map (
            O => \N__36367\,
            I => \N__36356\
        );

    \I__6216\ : Span4Mux_v
    port map (
            O => \N__36364\,
            I => \N__36353\
        );

    \I__6215\ : Span4Mux_v
    port map (
            O => \N__36359\,
            I => \N__36350\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__36356\,
            I => data_in_1_3
        );

    \I__6213\ : Odrv4
    port map (
            O => \N__36353\,
            I => data_in_1_3
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__36350\,
            I => data_in_1_3
        );

    \I__6211\ : InMux
    port map (
            O => \N__36343\,
            I => \N__36340\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__36340\,
            I => \N__36337\
        );

    \I__6209\ : Span4Mux_h
    port map (
            O => \N__36337\,
            I => \N__36334\
        );

    \I__6208\ : Odrv4
    port map (
            O => \N__36334\,
            I => \c0.n16_adj_4478\
        );

    \I__6207\ : InMux
    port map (
            O => \N__36331\,
            I => \N__36328\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__36328\,
            I => \N__36325\
        );

    \I__6205\ : Span4Mux_h
    port map (
            O => \N__36325\,
            I => \N__36320\
        );

    \I__6204\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36315\
        );

    \I__6203\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36315\
        );

    \I__6202\ : Odrv4
    port map (
            O => \N__36320\,
            I => data_in_1_1
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__36315\,
            I => data_in_1_1
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__36310\,
            I => \N__36307\
        );

    \I__6199\ : InMux
    port map (
            O => \N__36307\,
            I => \N__36304\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__36304\,
            I => \N__36301\
        );

    \I__6197\ : Span4Mux_h
    port map (
            O => \N__36301\,
            I => \N__36296\
        );

    \I__6196\ : InMux
    port map (
            O => \N__36300\,
            I => \N__36291\
        );

    \I__6195\ : InMux
    port map (
            O => \N__36299\,
            I => \N__36291\
        );

    \I__6194\ : Odrv4
    port map (
            O => \N__36296\,
            I => data_in_0_1
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__36291\,
            I => data_in_0_1
        );

    \I__6192\ : InMux
    port map (
            O => \N__36286\,
            I => \N__36282\
        );

    \I__6191\ : InMux
    port map (
            O => \N__36285\,
            I => \N__36279\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__36282\,
            I => \N__36276\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__36279\,
            I => data_out_frame_6_5
        );

    \I__6188\ : Odrv12
    port map (
            O => \N__36276\,
            I => data_out_frame_6_5
        );

    \I__6187\ : InMux
    port map (
            O => \N__36271\,
            I => \N__36268\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__36268\,
            I => n2256
        );

    \I__6185\ : CascadeMux
    port map (
            O => \N__36265\,
            I => \N__36262\
        );

    \I__6184\ : InMux
    port map (
            O => \N__36262\,
            I => \N__36259\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__36259\,
            I => \N__36253\
        );

    \I__6182\ : InMux
    port map (
            O => \N__36258\,
            I => \N__36249\
        );

    \I__6181\ : CascadeMux
    port map (
            O => \N__36257\,
            I => \N__36246\
        );

    \I__6180\ : InMux
    port map (
            O => \N__36256\,
            I => \N__36243\
        );

    \I__6179\ : Span4Mux_h
    port map (
            O => \N__36253\,
            I => \N__36240\
        );

    \I__6178\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36237\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__36249\,
            I => \N__36234\
        );

    \I__6176\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36231\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__36243\,
            I => encoder0_position_15
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__36240\,
            I => encoder0_position_15
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__36237\,
            I => encoder0_position_15
        );

    \I__6172\ : Odrv12
    port map (
            O => \N__36234\,
            I => encoder0_position_15
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__36231\,
            I => encoder0_position_15
        );

    \I__6170\ : InMux
    port map (
            O => \N__36220\,
            I => \N__36217\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__36217\,
            I => \N__36213\
        );

    \I__6168\ : CascadeMux
    port map (
            O => \N__36216\,
            I => \N__36210\
        );

    \I__6167\ : Span4Mux_v
    port map (
            O => \N__36213\,
            I => \N__36207\
        );

    \I__6166\ : InMux
    port map (
            O => \N__36210\,
            I => \N__36204\
        );

    \I__6165\ : Span4Mux_h
    port map (
            O => \N__36207\,
            I => \N__36201\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__36204\,
            I => \N__36198\
        );

    \I__6163\ : Span4Mux_h
    port map (
            O => \N__36201\,
            I => \N__36193\
        );

    \I__6162\ : Span4Mux_h
    port map (
            O => \N__36198\,
            I => \N__36190\
        );

    \I__6161\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36185\
        );

    \I__6160\ : InMux
    port map (
            O => \N__36196\,
            I => \N__36185\
        );

    \I__6159\ : Odrv4
    port map (
            O => \N__36193\,
            I => data_in_2_0
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__36190\,
            I => data_in_2_0
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__36185\,
            I => data_in_2_0
        );

    \I__6156\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36175\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__36175\,
            I => n2247
        );

    \I__6154\ : InMux
    port map (
            O => \N__36172\,
            I => \N__36169\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__36169\,
            I => n2265
        );

    \I__6152\ : InMux
    port map (
            O => \N__36166\,
            I => \N__36160\
        );

    \I__6151\ : InMux
    port map (
            O => \N__36165\,
            I => \N__36160\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__36160\,
            I => \N__36156\
        );

    \I__6149\ : InMux
    port map (
            O => \N__36159\,
            I => \N__36151\
        );

    \I__6148\ : Span4Mux_h
    port map (
            O => \N__36156\,
            I => \N__36148\
        );

    \I__6147\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36143\
        );

    \I__6146\ : InMux
    port map (
            O => \N__36154\,
            I => \N__36143\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__36151\,
            I => encoder0_position_6
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__36148\,
            I => encoder0_position_6
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__36143\,
            I => encoder0_position_6
        );

    \I__6142\ : CascadeMux
    port map (
            O => \N__36136\,
            I => \N__36133\
        );

    \I__6141\ : InMux
    port map (
            O => \N__36133\,
            I => \N__36130\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__36130\,
            I => \N__36127\
        );

    \I__6139\ : Span4Mux_v
    port map (
            O => \N__36127\,
            I => \N__36124\
        );

    \I__6138\ : Span4Mux_h
    port map (
            O => \N__36124\,
            I => \N__36118\
        );

    \I__6137\ : InMux
    port map (
            O => \N__36123\,
            I => \N__36115\
        );

    \I__6136\ : InMux
    port map (
            O => \N__36122\,
            I => \N__36112\
        );

    \I__6135\ : InMux
    port map (
            O => \N__36121\,
            I => \N__36108\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__36118\,
            I => \N__36105\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36100\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__36112\,
            I => \N__36100\
        );

    \I__6131\ : InMux
    port map (
            O => \N__36111\,
            I => \N__36097\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__36108\,
            I => encoder0_position_20
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__36105\,
            I => encoder0_position_20
        );

    \I__6128\ : Odrv4
    port map (
            O => \N__36100\,
            I => encoder0_position_20
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__36097\,
            I => encoder0_position_20
        );

    \I__6126\ : InMux
    port map (
            O => \N__36088\,
            I => \N__36085\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__36085\,
            I => n2266
        );

    \I__6124\ : CascadeMux
    port map (
            O => \N__36082\,
            I => \N__36079\
        );

    \I__6123\ : InMux
    port map (
            O => \N__36079\,
            I => \N__36075\
        );

    \I__6122\ : CascadeMux
    port map (
            O => \N__36078\,
            I => \N__36072\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__36075\,
            I => \N__36069\
        );

    \I__6120\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36066\
        );

    \I__6119\ : Span4Mux_h
    port map (
            O => \N__36069\,
            I => \N__36063\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__36066\,
            I => \N__36059\
        );

    \I__6117\ : Span4Mux_h
    port map (
            O => \N__36063\,
            I => \N__36053\
        );

    \I__6116\ : InMux
    port map (
            O => \N__36062\,
            I => \N__36050\
        );

    \I__6115\ : Span4Mux_h
    port map (
            O => \N__36059\,
            I => \N__36047\
        );

    \I__6114\ : InMux
    port map (
            O => \N__36058\,
            I => \N__36044\
        );

    \I__6113\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36039\
        );

    \I__6112\ : InMux
    port map (
            O => \N__36056\,
            I => \N__36039\
        );

    \I__6111\ : Odrv4
    port map (
            O => \N__36053\,
            I => encoder0_position_5
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__36050\,
            I => encoder0_position_5
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__36047\,
            I => encoder0_position_5
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__36044\,
            I => encoder0_position_5
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__36039\,
            I => encoder0_position_5
        );

    \I__6106\ : InMux
    port map (
            O => \N__36028\,
            I => \N__36024\
        );

    \I__6105\ : InMux
    port map (
            O => \N__36027\,
            I => \N__36021\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__36024\,
            I => \N__36018\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__36021\,
            I => \N__36015\
        );

    \I__6102\ : Odrv12
    port map (
            O => \N__36018\,
            I => \c0.n21808\
        );

    \I__6101\ : Odrv4
    port map (
            O => \N__36015\,
            I => \c0.n21808\
        );

    \I__6100\ : InMux
    port map (
            O => \N__36010\,
            I => \N__36007\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__36007\,
            I => n2250
        );

    \I__6098\ : CascadeMux
    port map (
            O => \N__36004\,
            I => \N__36001\
        );

    \I__6097\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35998\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__35998\,
            I => \N__35994\
        );

    \I__6095\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35990\
        );

    \I__6094\ : Span4Mux_h
    port map (
            O => \N__35994\,
            I => \N__35986\
        );

    \I__6093\ : CascadeMux
    port map (
            O => \N__35993\,
            I => \N__35983\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__35990\,
            I => \N__35980\
        );

    \I__6091\ : InMux
    port map (
            O => \N__35989\,
            I => \N__35976\
        );

    \I__6090\ : Span4Mux_h
    port map (
            O => \N__35986\,
            I => \N__35973\
        );

    \I__6089\ : InMux
    port map (
            O => \N__35983\,
            I => \N__35970\
        );

    \I__6088\ : Span4Mux_h
    port map (
            O => \N__35980\,
            I => \N__35967\
        );

    \I__6087\ : InMux
    port map (
            O => \N__35979\,
            I => \N__35964\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__35976\,
            I => encoder0_position_21
        );

    \I__6085\ : Odrv4
    port map (
            O => \N__35973\,
            I => encoder0_position_21
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__35970\,
            I => encoder0_position_21
        );

    \I__6083\ : Odrv4
    port map (
            O => \N__35967\,
            I => encoder0_position_21
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__35964\,
            I => encoder0_position_21
        );

    \I__6081\ : InMux
    port map (
            O => \N__35953\,
            I => \N__35950\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__35950\,
            I => n2262
        );

    \I__6079\ : InMux
    port map (
            O => \N__35947\,
            I => \N__35944\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__35944\,
            I => \N__35941\
        );

    \I__6077\ : Odrv12
    port map (
            O => \N__35941\,
            I => n2260
        );

    \I__6076\ : InMux
    port map (
            O => \N__35938\,
            I => \N__35935\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__35935\,
            I => n2254
        );

    \I__6074\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35929\
        );

    \I__6073\ : LocalMux
    port map (
            O => \N__35929\,
            I => \N__35925\
        );

    \I__6072\ : InMux
    port map (
            O => \N__35928\,
            I => \N__35922\
        );

    \I__6071\ : Span4Mux_h
    port map (
            O => \N__35925\,
            I => \N__35919\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__35922\,
            I => \N__35916\
        );

    \I__6069\ : Odrv4
    port map (
            O => \N__35919\,
            I => \c0.n10394\
        );

    \I__6068\ : Odrv12
    port map (
            O => \N__35916\,
            I => \c0.n10394\
        );

    \I__6067\ : InMux
    port map (
            O => \N__35911\,
            I => \N__35908\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__35908\,
            I => \N__35905\
        );

    \I__6065\ : Span4Mux_h
    port map (
            O => \N__35905\,
            I => \N__35902\
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__35902\,
            I => \c0.n20328\
        );

    \I__6063\ : CascadeMux
    port map (
            O => \N__35899\,
            I => \N__35896\
        );

    \I__6062\ : InMux
    port map (
            O => \N__35896\,
            I => \N__35892\
        );

    \I__6061\ : InMux
    port map (
            O => \N__35895\,
            I => \N__35887\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__35892\,
            I => \N__35884\
        );

    \I__6059\ : InMux
    port map (
            O => \N__35891\,
            I => \N__35881\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__35890\,
            I => \N__35878\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__35887\,
            I => \N__35874\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__35884\,
            I => \N__35869\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__35881\,
            I => \N__35866\
        );

    \I__6054\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35861\
        );

    \I__6053\ : InMux
    port map (
            O => \N__35877\,
            I => \N__35861\
        );

    \I__6052\ : Span4Mux_h
    port map (
            O => \N__35874\,
            I => \N__35858\
        );

    \I__6051\ : InMux
    port map (
            O => \N__35873\,
            I => \N__35853\
        );

    \I__6050\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35853\
        );

    \I__6049\ : Odrv4
    port map (
            O => \N__35869\,
            I => encoder0_position_14
        );

    \I__6048\ : Odrv4
    port map (
            O => \N__35866\,
            I => encoder0_position_14
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__35861\,
            I => encoder0_position_14
        );

    \I__6046\ : Odrv4
    port map (
            O => \N__35858\,
            I => encoder0_position_14
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__35853\,
            I => encoder0_position_14
        );

    \I__6044\ : CascadeMux
    port map (
            O => \N__35842\,
            I => \c0.n20328_cascade_\
        );

    \I__6043\ : InMux
    port map (
            O => \N__35839\,
            I => \N__35836\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__35836\,
            I => \N__35833\
        );

    \I__6041\ : Span4Mux_h
    port map (
            O => \N__35833\,
            I => \N__35830\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__35830\,
            I => \c0.n22367\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__35827\,
            I => \c0.n22367_cascade_\
        );

    \I__6038\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35821\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__35821\,
            I => \c0.n23569\
        );

    \I__6036\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35815\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__35815\,
            I => n2271
        );

    \I__6034\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35807\
        );

    \I__6033\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35804\
        );

    \I__6032\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35801\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__35807\,
            I => \c0.n10_adj_4331\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__35804\,
            I => \c0.n10_adj_4331\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__35801\,
            I => \c0.n10_adj_4331\
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__35794\,
            I => \N__35791\
        );

    \I__6027\ : InMux
    port map (
            O => \N__35791\,
            I => \N__35788\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__35788\,
            I => \N__35784\
        );

    \I__6025\ : InMux
    port map (
            O => \N__35787\,
            I => \N__35781\
        );

    \I__6024\ : Odrv12
    port map (
            O => \N__35784\,
            I => \c0.n22230\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__35781\,
            I => \c0.n22230\
        );

    \I__6022\ : CascadeMux
    port map (
            O => \N__35776\,
            I => \N__35773\
        );

    \I__6021\ : InMux
    port map (
            O => \N__35773\,
            I => \N__35769\
        );

    \I__6020\ : InMux
    port map (
            O => \N__35772\,
            I => \N__35766\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__35769\,
            I => \N__35759\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__35766\,
            I => \N__35756\
        );

    \I__6017\ : InMux
    port map (
            O => \N__35765\,
            I => \N__35753\
        );

    \I__6016\ : InMux
    port map (
            O => \N__35764\,
            I => \N__35750\
        );

    \I__6015\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35747\
        );

    \I__6014\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35744\
        );

    \I__6013\ : Span4Mux_v
    port map (
            O => \N__35759\,
            I => \N__35739\
        );

    \I__6012\ : Span4Mux_h
    port map (
            O => \N__35756\,
            I => \N__35739\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__35753\,
            I => encoder0_position_1
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__35750\,
            I => encoder0_position_1
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__35747\,
            I => encoder0_position_1
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__35744\,
            I => encoder0_position_1
        );

    \I__6007\ : Odrv4
    port map (
            O => \N__35739\,
            I => encoder0_position_1
        );

    \I__6006\ : CascadeMux
    port map (
            O => \N__35728\,
            I => \c0.n22461_cascade_\
        );

    \I__6005\ : InMux
    port map (
            O => \N__35725\,
            I => \N__35720\
        );

    \I__6004\ : CascadeMux
    port map (
            O => \N__35724\,
            I => \N__35717\
        );

    \I__6003\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35714\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__35720\,
            I => \N__35710\
        );

    \I__6001\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35707\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__35714\,
            I => \N__35704\
        );

    \I__5999\ : InMux
    port map (
            O => \N__35713\,
            I => \N__35698\
        );

    \I__5998\ : Span12Mux_h
    port map (
            O => \N__35710\,
            I => \N__35695\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__35707\,
            I => \N__35690\
        );

    \I__5996\ : Span4Mux_h
    port map (
            O => \N__35704\,
            I => \N__35690\
        );

    \I__5995\ : InMux
    port map (
            O => \N__35703\,
            I => \N__35687\
        );

    \I__5994\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35684\
        );

    \I__5993\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35681\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__35698\,
            I => encoder0_position_13
        );

    \I__5991\ : Odrv12
    port map (
            O => \N__35695\,
            I => encoder0_position_13
        );

    \I__5990\ : Odrv4
    port map (
            O => \N__35690\,
            I => encoder0_position_13
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__35687\,
            I => encoder0_position_13
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__35684\,
            I => encoder0_position_13
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__35681\,
            I => encoder0_position_13
        );

    \I__5986\ : InMux
    port map (
            O => \N__35668\,
            I => \N__35665\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__35665\,
            I => \N__35662\
        );

    \I__5984\ : Odrv4
    port map (
            O => \N__35662\,
            I => \c0.n20_adj_4318\
        );

    \I__5983\ : CascadeMux
    port map (
            O => \N__35659\,
            I => \N__35656\
        );

    \I__5982\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35652\
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__35655\,
            I => \N__35649\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__35652\,
            I => \N__35646\
        );

    \I__5979\ : InMux
    port map (
            O => \N__35649\,
            I => \N__35641\
        );

    \I__5978\ : Span4Mux_h
    port map (
            O => \N__35646\,
            I => \N__35638\
        );

    \I__5977\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35635\
        );

    \I__5976\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35632\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__35641\,
            I => \N__35629\
        );

    \I__5974\ : Sp12to4
    port map (
            O => \N__35638\,
            I => \N__35624\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__35635\,
            I => \N__35624\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__35632\,
            I => \N__35619\
        );

    \I__5971\ : Span4Mux_h
    port map (
            O => \N__35629\,
            I => \N__35619\
        );

    \I__5970\ : Odrv12
    port map (
            O => \N__35624\,
            I => encoder1_position_26
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__35619\,
            I => encoder1_position_26
        );

    \I__5968\ : InMux
    port map (
            O => \N__35614\,
            I => \N__35611\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__35611\,
            I => \N__35606\
        );

    \I__5966\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35600\
        );

    \I__5965\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35600\
        );

    \I__5964\ : Span4Mux_v
    port map (
            O => \N__35606\,
            I => \N__35597\
        );

    \I__5963\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35594\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__35600\,
            I => \N__35591\
        );

    \I__5961\ : Span4Mux_h
    port map (
            O => \N__35597\,
            I => \N__35587\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__35594\,
            I => \N__35582\
        );

    \I__5959\ : Span4Mux_h
    port map (
            O => \N__35591\,
            I => \N__35582\
        );

    \I__5958\ : InMux
    port map (
            O => \N__35590\,
            I => \N__35579\
        );

    \I__5957\ : Odrv4
    port map (
            O => \N__35587\,
            I => \c0.n20236\
        );

    \I__5956\ : Odrv4
    port map (
            O => \N__35582\,
            I => \c0.n20236\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__35579\,
            I => \c0.n20236\
        );

    \I__5954\ : InMux
    port map (
            O => \N__35572\,
            I => \N__35569\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__35569\,
            I => \N__35565\
        );

    \I__5952\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35562\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__35565\,
            I => \N__35559\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__35562\,
            I => \N__35556\
        );

    \I__5949\ : Span4Mux_v
    port map (
            O => \N__35559\,
            I => \N__35553\
        );

    \I__5948\ : Span4Mux_v
    port map (
            O => \N__35556\,
            I => \N__35550\
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__35553\,
            I => \c0.n22449\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__35550\,
            I => \c0.n22449\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__35545\,
            I => \N__35542\
        );

    \I__5944\ : InMux
    port map (
            O => \N__35542\,
            I => \N__35539\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__35539\,
            I => \c0.n22474\
        );

    \I__5942\ : InMux
    port map (
            O => \N__35536\,
            I => \N__35533\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__35533\,
            I => \c0.n22483\
        );

    \I__5940\ : CascadeMux
    port map (
            O => \N__35530\,
            I => \N__35526\
        );

    \I__5939\ : InMux
    port map (
            O => \N__35529\,
            I => \N__35523\
        );

    \I__5938\ : InMux
    port map (
            O => \N__35526\,
            I => \N__35520\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__35523\,
            I => \N__35514\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__35520\,
            I => \N__35511\
        );

    \I__5935\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35508\
        );

    \I__5934\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35505\
        );

    \I__5933\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35502\
        );

    \I__5932\ : Span4Mux_h
    port map (
            O => \N__35514\,
            I => \N__35499\
        );

    \I__5931\ : Span4Mux_h
    port map (
            O => \N__35511\,
            I => \N__35496\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__35508\,
            I => \N__35493\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__35505\,
            I => \N__35486\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__35502\,
            I => \N__35486\
        );

    \I__5927\ : Span4Mux_v
    port map (
            O => \N__35499\,
            I => \N__35486\
        );

    \I__5926\ : Odrv4
    port map (
            O => \N__35496\,
            I => encoder1_position_30
        );

    \I__5925\ : Odrv12
    port map (
            O => \N__35493\,
            I => encoder1_position_30
        );

    \I__5924\ : Odrv4
    port map (
            O => \N__35486\,
            I => encoder1_position_30
        );

    \I__5923\ : CascadeMux
    port map (
            O => \N__35479\,
            I => \c0.n16_adj_4321_cascade_\
        );

    \I__5922\ : CascadeMux
    port map (
            O => \N__35476\,
            I => \c0.n18_adj_4322_cascade_\
        );

    \I__5921\ : InMux
    port map (
            O => \N__35473\,
            I => \N__35470\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__35470\,
            I => \N__35467\
        );

    \I__5919\ : Span4Mux_h
    port map (
            O => \N__35467\,
            I => \N__35464\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__35464\,
            I => \c0.n17_adj_4323\
        );

    \I__5917\ : InMux
    port map (
            O => \N__35461\,
            I => \N__35458\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__35458\,
            I => \N__35455\
        );

    \I__5915\ : Span4Mux_v
    port map (
            O => \N__35455\,
            I => \N__35452\
        );

    \I__5914\ : Odrv4
    port map (
            O => \N__35452\,
            I => \c0.n14_adj_4324\
        );

    \I__5913\ : InMux
    port map (
            O => \N__35449\,
            I => \N__35446\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__35446\,
            I => \N__35442\
        );

    \I__5911\ : InMux
    port map (
            O => \N__35445\,
            I => \N__35439\
        );

    \I__5910\ : Span12Mux_v
    port map (
            O => \N__35442\,
            I => \N__35434\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__35439\,
            I => \N__35434\
        );

    \I__5908\ : Odrv12
    port map (
            O => \N__35434\,
            I => \c0.n22376\
        );

    \I__5907\ : InMux
    port map (
            O => \N__35431\,
            I => \N__35428\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__35428\,
            I => \c0.n13619\
        );

    \I__5905\ : CascadeMux
    port map (
            O => \N__35425\,
            I => \c0.n13619_cascade_\
        );

    \I__5904\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35419\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__35419\,
            I => \N__35415\
        );

    \I__5902\ : InMux
    port map (
            O => \N__35418\,
            I => \N__35412\
        );

    \I__5901\ : Span4Mux_h
    port map (
            O => \N__35415\,
            I => \N__35409\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__35412\,
            I => \c0.n22412\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__35409\,
            I => \c0.n22412\
        );

    \I__5898\ : CascadeMux
    port map (
            O => \N__35404\,
            I => \c0.n13524_cascade_\
        );

    \I__5897\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35398\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__35398\,
            I => \c0.n10_adj_4317\
        );

    \I__5895\ : CascadeMux
    port map (
            O => \N__35395\,
            I => \N__35392\
        );

    \I__5894\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35387\
        );

    \I__5893\ : InMux
    port map (
            O => \N__35391\,
            I => \N__35382\
        );

    \I__5892\ : InMux
    port map (
            O => \N__35390\,
            I => \N__35378\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__35387\,
            I => \N__35375\
        );

    \I__5890\ : InMux
    port map (
            O => \N__35386\,
            I => \N__35370\
        );

    \I__5889\ : InMux
    port map (
            O => \N__35385\,
            I => \N__35370\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__35382\,
            I => \N__35366\
        );

    \I__5887\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35363\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__35378\,
            I => \N__35360\
        );

    \I__5885\ : Span4Mux_h
    port map (
            O => \N__35375\,
            I => \N__35355\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__35370\,
            I => \N__35355\
        );

    \I__5883\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35352\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__35366\,
            I => encoder1_position_8
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__35363\,
            I => encoder1_position_8
        );

    \I__5880\ : Odrv4
    port map (
            O => \N__35360\,
            I => encoder1_position_8
        );

    \I__5879\ : Odrv4
    port map (
            O => \N__35355\,
            I => encoder1_position_8
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__35352\,
            I => encoder1_position_8
        );

    \I__5877\ : InMux
    port map (
            O => \N__35341\,
            I => \N__35338\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__35338\,
            I => \N__35335\
        );

    \I__5875\ : Span4Mux_h
    port map (
            O => \N__35335\,
            I => \N__35331\
        );

    \I__5874\ : InMux
    port map (
            O => \N__35334\,
            I => \N__35328\
        );

    \I__5873\ : Span4Mux_h
    port map (
            O => \N__35331\,
            I => \N__35325\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__35328\,
            I => data_out_frame_12_0
        );

    \I__5871\ : Odrv4
    port map (
            O => \N__35325\,
            I => data_out_frame_12_0
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__35320\,
            I => \N__35317\
        );

    \I__5869\ : InMux
    port map (
            O => \N__35317\,
            I => \N__35311\
        );

    \I__5868\ : InMux
    port map (
            O => \N__35316\,
            I => \N__35311\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__35311\,
            I => \N__35305\
        );

    \I__5866\ : InMux
    port map (
            O => \N__35310\,
            I => \N__35300\
        );

    \I__5865\ : InMux
    port map (
            O => \N__35309\,
            I => \N__35300\
        );

    \I__5864\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35297\
        );

    \I__5863\ : Span4Mux_v
    port map (
            O => \N__35305\,
            I => \N__35294\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__35300\,
            I => \N__35289\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__35297\,
            I => \N__35289\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__35294\,
            I => \c0.n13079\
        );

    \I__5859\ : Odrv12
    port map (
            O => \N__35289\,
            I => \c0.n13079\
        );

    \I__5858\ : InMux
    port map (
            O => \N__35284\,
            I => \N__35280\
        );

    \I__5857\ : CascadeMux
    port map (
            O => \N__35283\,
            I => \N__35277\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__35280\,
            I => \N__35274\
        );

    \I__5855\ : InMux
    port map (
            O => \N__35277\,
            I => \N__35271\
        );

    \I__5854\ : Span4Mux_v
    port map (
            O => \N__35274\,
            I => \N__35268\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__35271\,
            I => \N__35265\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__35268\,
            I => \c0.n22174\
        );

    \I__5851\ : Odrv12
    port map (
            O => \N__35265\,
            I => \c0.n22174\
        );

    \I__5850\ : CascadeMux
    port map (
            O => \N__35260\,
            I => \N__35257\
        );

    \I__5849\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35254\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__35254\,
            I => \N__35249\
        );

    \I__5847\ : InMux
    port map (
            O => \N__35253\,
            I => \N__35246\
        );

    \I__5846\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35242\
        );

    \I__5845\ : Span4Mux_h
    port map (
            O => \N__35249\,
            I => \N__35239\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__35246\,
            I => \N__35236\
        );

    \I__5843\ : InMux
    port map (
            O => \N__35245\,
            I => \N__35233\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__35242\,
            I => \N__35226\
        );

    \I__5841\ : Sp12to4
    port map (
            O => \N__35239\,
            I => \N__35226\
        );

    \I__5840\ : Span12Mux_h
    port map (
            O => \N__35236\,
            I => \N__35226\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__35233\,
            I => data_in_3_5
        );

    \I__5838\ : Odrv12
    port map (
            O => \N__35226\,
            I => data_in_3_5
        );

    \I__5837\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35217\
        );

    \I__5836\ : InMux
    port map (
            O => \N__35220\,
            I => \N__35214\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__35217\,
            I => \N__35210\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__35214\,
            I => \N__35205\
        );

    \I__5833\ : InMux
    port map (
            O => \N__35213\,
            I => \N__35202\
        );

    \I__5832\ : Span12Mux_h
    port map (
            O => \N__35210\,
            I => \N__35197\
        );

    \I__5831\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35194\
        );

    \I__5830\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35191\
        );

    \I__5829\ : Span4Mux_h
    port map (
            O => \N__35205\,
            I => \N__35186\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__35202\,
            I => \N__35186\
        );

    \I__5827\ : InMux
    port map (
            O => \N__35201\,
            I => \N__35181\
        );

    \I__5826\ : InMux
    port map (
            O => \N__35200\,
            I => \N__35181\
        );

    \I__5825\ : Odrv12
    port map (
            O => \N__35197\,
            I => encoder1_position_10
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__35194\,
            I => encoder1_position_10
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__35191\,
            I => encoder1_position_10
        );

    \I__5822\ : Odrv4
    port map (
            O => \N__35186\,
            I => encoder1_position_10
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__35181\,
            I => encoder1_position_10
        );

    \I__5820\ : InMux
    port map (
            O => \N__35170\,
            I => \N__35166\
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__35169\,
            I => \N__35163\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__35166\,
            I => \N__35160\
        );

    \I__5817\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35157\
        );

    \I__5816\ : Span4Mux_v
    port map (
            O => \N__35160\,
            I => \N__35154\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__35157\,
            I => data_out_frame_12_2
        );

    \I__5814\ : Odrv4
    port map (
            O => \N__35154\,
            I => data_out_frame_12_2
        );

    \I__5813\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35146\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__35146\,
            I => \N__35143\
        );

    \I__5811\ : Odrv12
    port map (
            O => \N__35143\,
            I => \c0.n21918\
        );

    \I__5810\ : CascadeMux
    port map (
            O => \N__35140\,
            I => \N__35136\
        );

    \I__5809\ : InMux
    port map (
            O => \N__35139\,
            I => \N__35131\
        );

    \I__5808\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35128\
        );

    \I__5807\ : InMux
    port map (
            O => \N__35135\,
            I => \N__35123\
        );

    \I__5806\ : InMux
    port map (
            O => \N__35134\,
            I => \N__35123\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__35131\,
            I => \N__35117\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__35128\,
            I => \N__35111\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__35123\,
            I => \N__35111\
        );

    \I__5802\ : InMux
    port map (
            O => \N__35122\,
            I => \N__35108\
        );

    \I__5801\ : InMux
    port map (
            O => \N__35121\,
            I => \N__35103\
        );

    \I__5800\ : InMux
    port map (
            O => \N__35120\,
            I => \N__35103\
        );

    \I__5799\ : Span4Mux_v
    port map (
            O => \N__35117\,
            I => \N__35100\
        );

    \I__5798\ : InMux
    port map (
            O => \N__35116\,
            I => \N__35097\
        );

    \I__5797\ : Span4Mux_h
    port map (
            O => \N__35111\,
            I => \N__35094\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__35108\,
            I => \N__35091\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__35103\,
            I => encoder1_position_4
        );

    \I__5794\ : Odrv4
    port map (
            O => \N__35100\,
            I => encoder1_position_4
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__35097\,
            I => encoder1_position_4
        );

    \I__5792\ : Odrv4
    port map (
            O => \N__35094\,
            I => encoder1_position_4
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__35091\,
            I => encoder1_position_4
        );

    \I__5790\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35076\
        );

    \I__5789\ : InMux
    port map (
            O => \N__35079\,
            I => \N__35073\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__35076\,
            I => \N__35070\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__35073\,
            I => data_out_frame_13_4
        );

    \I__5786\ : Odrv4
    port map (
            O => \N__35070\,
            I => data_out_frame_13_4
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__35065\,
            I => \N__35061\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__35064\,
            I => \N__35058\
        );

    \I__5783\ : InMux
    port map (
            O => \N__35061\,
            I => \N__35054\
        );

    \I__5782\ : InMux
    port map (
            O => \N__35058\,
            I => \N__35051\
        );

    \I__5781\ : InMux
    port map (
            O => \N__35057\,
            I => \N__35048\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__35054\,
            I => \N__35043\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__35051\,
            I => \N__35043\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__35048\,
            I => \N__35039\
        );

    \I__5777\ : Span4Mux_h
    port map (
            O => \N__35043\,
            I => \N__35036\
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__35042\,
            I => \N__35032\
        );

    \I__5775\ : Span4Mux_h
    port map (
            O => \N__35039\,
            I => \N__35027\
        );

    \I__5774\ : Span4Mux_h
    port map (
            O => \N__35036\,
            I => \N__35024\
        );

    \I__5773\ : InMux
    port map (
            O => \N__35035\,
            I => \N__35021\
        );

    \I__5772\ : InMux
    port map (
            O => \N__35032\,
            I => \N__35016\
        );

    \I__5771\ : InMux
    port map (
            O => \N__35031\,
            I => \N__35016\
        );

    \I__5770\ : InMux
    port map (
            O => \N__35030\,
            I => \N__35013\
        );

    \I__5769\ : Odrv4
    port map (
            O => \N__35027\,
            I => encoder1_position_2
        );

    \I__5768\ : Odrv4
    port map (
            O => \N__35024\,
            I => encoder1_position_2
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__35021\,
            I => encoder1_position_2
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__35016\,
            I => encoder1_position_2
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__35013\,
            I => encoder1_position_2
        );

    \I__5764\ : InMux
    port map (
            O => \N__35002\,
            I => \N__34999\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__34999\,
            I => \N__34995\
        );

    \I__5762\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34992\
        );

    \I__5761\ : Span4Mux_h
    port map (
            O => \N__34995\,
            I => \N__34989\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__34992\,
            I => data_out_frame_13_2
        );

    \I__5759\ : Odrv4
    port map (
            O => \N__34989\,
            I => data_out_frame_13_2
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__34984\,
            I => \N__34981\
        );

    \I__5757\ : InMux
    port map (
            O => \N__34981\,
            I => \N__34975\
        );

    \I__5756\ : InMux
    port map (
            O => \N__34980\,
            I => \N__34972\
        );

    \I__5755\ : InMux
    port map (
            O => \N__34979\,
            I => \N__34967\
        );

    \I__5754\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34967\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__34975\,
            I => \N__34963\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__34972\,
            I => \N__34958\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__34967\,
            I => \N__34958\
        );

    \I__5750\ : CascadeMux
    port map (
            O => \N__34966\,
            I => \N__34954\
        );

    \I__5749\ : Span4Mux_v
    port map (
            O => \N__34963\,
            I => \N__34949\
        );

    \I__5748\ : Span4Mux_h
    port map (
            O => \N__34958\,
            I => \N__34949\
        );

    \I__5747\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34946\
        );

    \I__5746\ : InMux
    port map (
            O => \N__34954\,
            I => \N__34943\
        );

    \I__5745\ : Span4Mux_h
    port map (
            O => \N__34949\,
            I => \N__34940\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__34946\,
            I => encoder1_position_6
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__34943\,
            I => encoder1_position_6
        );

    \I__5742\ : Odrv4
    port map (
            O => \N__34940\,
            I => encoder1_position_6
        );

    \I__5741\ : CascadeMux
    port map (
            O => \N__34933\,
            I => \N__34930\
        );

    \I__5740\ : InMux
    port map (
            O => \N__34930\,
            I => \N__34922\
        );

    \I__5739\ : CascadeMux
    port map (
            O => \N__34929\,
            I => \N__34919\
        );

    \I__5738\ : InMux
    port map (
            O => \N__34928\,
            I => \N__34916\
        );

    \I__5737\ : InMux
    port map (
            O => \N__34927\,
            I => \N__34913\
        );

    \I__5736\ : InMux
    port map (
            O => \N__34926\,
            I => \N__34908\
        );

    \I__5735\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34908\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__34922\,
            I => \N__34904\
        );

    \I__5733\ : InMux
    port map (
            O => \N__34919\,
            I => \N__34901\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__34916\,
            I => \N__34898\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__34913\,
            I => \N__34893\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__34908\,
            I => \N__34893\
        );

    \I__5729\ : InMux
    port map (
            O => \N__34907\,
            I => \N__34890\
        );

    \I__5728\ : Span4Mux_h
    port map (
            O => \N__34904\,
            I => \N__34887\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__34901\,
            I => \N__34884\
        );

    \I__5726\ : Span4Mux_v
    port map (
            O => \N__34898\,
            I => \N__34879\
        );

    \I__5725\ : Span4Mux_h
    port map (
            O => \N__34893\,
            I => \N__34879\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__34890\,
            I => encoder1_position_7
        );

    \I__5723\ : Odrv4
    port map (
            O => \N__34887\,
            I => encoder1_position_7
        );

    \I__5722\ : Odrv12
    port map (
            O => \N__34884\,
            I => encoder1_position_7
        );

    \I__5721\ : Odrv4
    port map (
            O => \N__34879\,
            I => encoder1_position_7
        );

    \I__5720\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34867\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__34867\,
            I => \N__34864\
        );

    \I__5718\ : Odrv4
    port map (
            O => \N__34864\,
            I => \c0.n21896\
        );

    \I__5717\ : InMux
    port map (
            O => \N__34861\,
            I => \N__34858\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__34858\,
            I => \N__34854\
        );

    \I__5715\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34851\
        );

    \I__5714\ : Span4Mux_v
    port map (
            O => \N__34854\,
            I => \N__34845\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__34851\,
            I => \N__34845\
        );

    \I__5712\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34842\
        );

    \I__5711\ : Span4Mux_h
    port map (
            O => \N__34845\,
            I => \N__34839\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__34842\,
            I => \c0.n21998\
        );

    \I__5709\ : Odrv4
    port map (
            O => \N__34839\,
            I => \c0.n21998\
        );

    \I__5708\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34831\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__34831\,
            I => \c0.n21852\
        );

    \I__5706\ : InMux
    port map (
            O => \N__34828\,
            I => \N__34824\
        );

    \I__5705\ : CascadeMux
    port map (
            O => \N__34827\,
            I => \N__34821\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__34824\,
            I => \N__34818\
        );

    \I__5703\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34814\
        );

    \I__5702\ : Span4Mux_h
    port map (
            O => \N__34818\,
            I => \N__34811\
        );

    \I__5701\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34808\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__34814\,
            I => \c0.n20249\
        );

    \I__5699\ : Odrv4
    port map (
            O => \N__34811\,
            I => \c0.n20249\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__34808\,
            I => \c0.n20249\
        );

    \I__5697\ : InMux
    port map (
            O => \N__34801\,
            I => \N__34798\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__34798\,
            I => \N__34795\
        );

    \I__5695\ : Span4Mux_v
    port map (
            O => \N__34795\,
            I => \N__34789\
        );

    \I__5694\ : InMux
    port map (
            O => \N__34794\,
            I => \N__34784\
        );

    \I__5693\ : InMux
    port map (
            O => \N__34793\,
            I => \N__34784\
        );

    \I__5692\ : InMux
    port map (
            O => \N__34792\,
            I => \N__34781\
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__34789\,
            I => \c0.n21210\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__34784\,
            I => \c0.n21210\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__34781\,
            I => \c0.n21210\
        );

    \I__5688\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34771\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__34771\,
            I => \c0.n17_adj_4499\
        );

    \I__5686\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34765\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34762\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__34762\,
            I => \c0.data_out_frame_29_7\
        );

    \I__5683\ : InMux
    port map (
            O => \N__34759\,
            I => \N__34756\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__34756\,
            I => \c0.data_out_frame_28_7\
        );

    \I__5681\ : InMux
    port map (
            O => \N__34753\,
            I => \N__34750\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__34750\,
            I => \N__34747\
        );

    \I__5679\ : Span4Mux_h
    port map (
            O => \N__34747\,
            I => \N__34744\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__34744\,
            I => \N__34741\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__34741\,
            I => \N__34738\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__34738\,
            I => \c0.n26_adj_4359\
        );

    \I__5675\ : InMux
    port map (
            O => \N__34735\,
            I => \N__34732\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__34732\,
            I => \N__34728\
        );

    \I__5673\ : InMux
    port map (
            O => \N__34731\,
            I => \N__34725\
        );

    \I__5672\ : Span4Mux_h
    port map (
            O => \N__34728\,
            I => \N__34722\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__34725\,
            I => data_out_frame_13_1
        );

    \I__5670\ : Odrv4
    port map (
            O => \N__34722\,
            I => data_out_frame_13_1
        );

    \I__5669\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34714\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__34714\,
            I => \N__34711\
        );

    \I__5667\ : Span4Mux_h
    port map (
            O => \N__34711\,
            I => \N__34707\
        );

    \I__5666\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34704\
        );

    \I__5665\ : Span4Mux_h
    port map (
            O => \N__34707\,
            I => \N__34701\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__34704\,
            I => data_out_frame_12_1
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__34701\,
            I => data_out_frame_12_1
        );

    \I__5662\ : CascadeMux
    port map (
            O => \N__34696\,
            I => \N__34693\
        );

    \I__5661\ : InMux
    port map (
            O => \N__34693\,
            I => \N__34690\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__34690\,
            I => \N__34687\
        );

    \I__5659\ : Span4Mux_v
    port map (
            O => \N__34687\,
            I => \N__34684\
        );

    \I__5658\ : Span4Mux_h
    port map (
            O => \N__34684\,
            I => \N__34681\
        );

    \I__5657\ : Span4Mux_v
    port map (
            O => \N__34681\,
            I => \N__34678\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__34678\,
            I => \c0.n11_adj_4520\
        );

    \I__5655\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34672\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__34672\,
            I => \N__34669\
        );

    \I__5653\ : Span4Mux_v
    port map (
            O => \N__34669\,
            I => \N__34665\
        );

    \I__5652\ : InMux
    port map (
            O => \N__34668\,
            I => \N__34662\
        );

    \I__5651\ : Span4Mux_h
    port map (
            O => \N__34665\,
            I => \N__34659\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__34662\,
            I => data_out_frame_8_3
        );

    \I__5649\ : Odrv4
    port map (
            O => \N__34659\,
            I => data_out_frame_8_3
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__34654\,
            I => \N__34651\
        );

    \I__5647\ : InMux
    port map (
            O => \N__34651\,
            I => \N__34648\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__34648\,
            I => \N__34645\
        );

    \I__5645\ : Span4Mux_v
    port map (
            O => \N__34645\,
            I => \N__34642\
        );

    \I__5644\ : Span4Mux_h
    port map (
            O => \N__34642\,
            I => \N__34639\
        );

    \I__5643\ : Odrv4
    port map (
            O => \N__34639\,
            I => \c0.n11_adj_4303\
        );

    \I__5642\ : InMux
    port map (
            O => \N__34636\,
            I => \N__34632\
        );

    \I__5641\ : InMux
    port map (
            O => \N__34635\,
            I => \N__34628\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__34632\,
            I => \N__34624\
        );

    \I__5639\ : InMux
    port map (
            O => \N__34631\,
            I => \N__34618\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__34628\,
            I => \N__34615\
        );

    \I__5637\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34612\
        );

    \I__5636\ : Span4Mux_h
    port map (
            O => \N__34624\,
            I => \N__34609\
        );

    \I__5635\ : InMux
    port map (
            O => \N__34623\,
            I => \N__34602\
        );

    \I__5634\ : InMux
    port map (
            O => \N__34622\,
            I => \N__34602\
        );

    \I__5633\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34602\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__34618\,
            I => \N__34595\
        );

    \I__5631\ : Span4Mux_v
    port map (
            O => \N__34615\,
            I => \N__34595\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__34612\,
            I => \N__34595\
        );

    \I__5629\ : Odrv4
    port map (
            O => \N__34609\,
            I => encoder1_position_12
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__34602\,
            I => encoder1_position_12
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__34595\,
            I => encoder1_position_12
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__34588\,
            I => \N__34585\
        );

    \I__5625\ : InMux
    port map (
            O => \N__34585\,
            I => \N__34579\
        );

    \I__5624\ : InMux
    port map (
            O => \N__34584\,
            I => \N__34579\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__34579\,
            I => data_out_frame_12_4
        );

    \I__5622\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34573\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__34573\,
            I => \N__34570\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__34570\,
            I => \c0.n44_adj_4412\
        );

    \I__5619\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34559\
        );

    \I__5618\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34559\
        );

    \I__5617\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34556\
        );

    \I__5616\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34553\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__34559\,
            I => \N__34550\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__34556\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__34553\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__34550\,
            I => \c0.FRAME_MATCHER_state_14\
        );

    \I__5611\ : CascadeMux
    port map (
            O => \N__34543\,
            I => \N__34537\
        );

    \I__5610\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34534\
        );

    \I__5609\ : InMux
    port map (
            O => \N__34541\,
            I => \N__34531\
        );

    \I__5608\ : InMux
    port map (
            O => \N__34540\,
            I => \N__34526\
        );

    \I__5607\ : InMux
    port map (
            O => \N__34537\,
            I => \N__34526\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__34534\,
            I => \N__34523\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__34531\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__34526\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__5603\ : Odrv12
    port map (
            O => \N__34523\,
            I => \c0.FRAME_MATCHER_state_21\
        );

    \I__5602\ : SRMux
    port map (
            O => \N__34516\,
            I => \N__34513\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__34513\,
            I => \N__34510\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__34510\,
            I => \N__34507\
        );

    \I__5599\ : Odrv4
    port map (
            O => \N__34507\,
            I => \c0.n21368\
        );

    \I__5598\ : InMux
    port map (
            O => \N__34504\,
            I => \N__34497\
        );

    \I__5597\ : InMux
    port map (
            O => \N__34503\,
            I => \N__34497\
        );

    \I__5596\ : InMux
    port map (
            O => \N__34502\,
            I => \N__34494\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__34497\,
            I => \N__34491\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__34494\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__5593\ : Odrv12
    port map (
            O => \N__34491\,
            I => \c0.FRAME_MATCHER_state_29\
        );

    \I__5592\ : SRMux
    port map (
            O => \N__34486\,
            I => \N__34483\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__34483\,
            I => \N__34480\
        );

    \I__5590\ : Odrv12
    port map (
            O => \N__34480\,
            I => \c0.n21326\
        );

    \I__5589\ : InMux
    port map (
            O => \N__34477\,
            I => \N__34473\
        );

    \I__5588\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34470\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__34473\,
            I => \N__34467\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__34470\,
            I => \N__34464\
        );

    \I__5585\ : Span4Mux_v
    port map (
            O => \N__34467\,
            I => \N__34459\
        );

    \I__5584\ : Span4Mux_v
    port map (
            O => \N__34464\,
            I => \N__34459\
        );

    \I__5583\ : Odrv4
    port map (
            O => \N__34459\,
            I => \c0.n20658\
        );

    \I__5582\ : InMux
    port map (
            O => \N__34456\,
            I => \N__34449\
        );

    \I__5581\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34446\
        );

    \I__5580\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34438\
        );

    \I__5579\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34438\
        );

    \I__5578\ : InMux
    port map (
            O => \N__34452\,
            I => \N__34438\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__34449\,
            I => \N__34433\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__34446\,
            I => \N__34433\
        );

    \I__5575\ : InMux
    port map (
            O => \N__34445\,
            I => \N__34430\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__34438\,
            I => \N__34427\
        );

    \I__5573\ : Span4Mux_v
    port map (
            O => \N__34433\,
            I => \N__34421\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__34430\,
            I => \N__34421\
        );

    \I__5571\ : Span4Mux_h
    port map (
            O => \N__34427\,
            I => \N__34418\
        );

    \I__5570\ : InMux
    port map (
            O => \N__34426\,
            I => \N__34415\
        );

    \I__5569\ : Span4Mux_h
    port map (
            O => \N__34421\,
            I => \N__34412\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__34418\,
            I => \N__34409\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__34415\,
            I => \N__34406\
        );

    \I__5566\ : Odrv4
    port map (
            O => \N__34412\,
            I => \c0.n21152\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__34409\,
            I => \c0.n21152\
        );

    \I__5564\ : Odrv12
    port map (
            O => \N__34406\,
            I => \c0.n21152\
        );

    \I__5563\ : InMux
    port map (
            O => \N__34399\,
            I => \N__34395\
        );

    \I__5562\ : CascadeMux
    port map (
            O => \N__34398\,
            I => \N__34392\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__34395\,
            I => \N__34389\
        );

    \I__5560\ : InMux
    port map (
            O => \N__34392\,
            I => \N__34383\
        );

    \I__5559\ : Span4Mux_h
    port map (
            O => \N__34389\,
            I => \N__34380\
        );

    \I__5558\ : InMux
    port map (
            O => \N__34388\,
            I => \N__34373\
        );

    \I__5557\ : InMux
    port map (
            O => \N__34387\,
            I => \N__34373\
        );

    \I__5556\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34373\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__34383\,
            I => \c0.n21168\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__34380\,
            I => \c0.n21168\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__34373\,
            I => \c0.n21168\
        );

    \I__5552\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34363\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__34363\,
            I => \N__34359\
        );

    \I__5550\ : InMux
    port map (
            O => \N__34362\,
            I => \N__34356\
        );

    \I__5549\ : Span4Mux_h
    port map (
            O => \N__34359\,
            I => \N__34353\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__34356\,
            I => \c0.n12542\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__34353\,
            I => \c0.n12542\
        );

    \I__5546\ : InMux
    port map (
            O => \N__34348\,
            I => \N__34345\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__34345\,
            I => \N__34340\
        );

    \I__5544\ : InMux
    port map (
            O => \N__34344\,
            I => \N__34337\
        );

    \I__5543\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34334\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__34340\,
            I => \N__34329\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__34337\,
            I => \N__34329\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34326\
        );

    \I__5539\ : Span4Mux_h
    port map (
            O => \N__34329\,
            I => \N__34323\
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__34326\,
            I => \c0.n20180\
        );

    \I__5537\ : Odrv4
    port map (
            O => \N__34323\,
            I => \c0.n20180\
        );

    \I__5536\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34315\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__34315\,
            I => \c0.n23260\
        );

    \I__5534\ : CascadeMux
    port map (
            O => \N__34312\,
            I => \c0.n16_adj_4498_cascade_\
        );

    \I__5533\ : InMux
    port map (
            O => \N__34309\,
            I => \N__34303\
        );

    \I__5532\ : InMux
    port map (
            O => \N__34308\,
            I => \N__34303\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__34303\,
            I => \N__34298\
        );

    \I__5530\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34295\
        );

    \I__5529\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34292\
        );

    \I__5528\ : Span4Mux_h
    port map (
            O => \N__34298\,
            I => \N__34289\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__34295\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__34292\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__34289\,
            I => \c0.FRAME_MATCHER_state_22\
        );

    \I__5524\ : CascadeMux
    port map (
            O => \N__34282\,
            I => \c0.n14457_cascade_\
        );

    \I__5523\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34274\
        );

    \I__5522\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34269\
        );

    \I__5521\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34269\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__34274\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__34269\,
            I => \c0.FRAME_MATCHER_state_27\
        );

    \I__5518\ : SRMux
    port map (
            O => \N__34264\,
            I => \N__34261\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__34261\,
            I => \N__34258\
        );

    \I__5516\ : Span4Mux_h
    port map (
            O => \N__34258\,
            I => \N__34255\
        );

    \I__5515\ : Odrv4
    port map (
            O => \N__34255\,
            I => \c0.n21330\
        );

    \I__5514\ : CascadeMux
    port map (
            O => \N__34252\,
            I => \c0.n30_adj_4411_cascade_\
        );

    \I__5513\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34241\
        );

    \I__5512\ : InMux
    port map (
            O => \N__34248\,
            I => \N__34241\
        );

    \I__5511\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34238\
        );

    \I__5510\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34235\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__34241\,
            I => \N__34232\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__34238\,
            I => \N__34229\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__34235\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__5506\ : Odrv4
    port map (
            O => \N__34232\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__5505\ : Odrv4
    port map (
            O => \N__34229\,
            I => \c0.FRAME_MATCHER_state_8\
        );

    \I__5504\ : SRMux
    port map (
            O => \N__34222\,
            I => \N__34219\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__34219\,
            I => \N__34216\
        );

    \I__5502\ : Span4Mux_h
    port map (
            O => \N__34216\,
            I => \N__34213\
        );

    \I__5501\ : Odrv4
    port map (
            O => \N__34213\,
            I => \c0.n21344\
        );

    \I__5500\ : SRMux
    port map (
            O => \N__34210\,
            I => \N__34207\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__34207\,
            I => \N__34204\
        );

    \I__5498\ : Span4Mux_h
    port map (
            O => \N__34204\,
            I => \N__34201\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__34201\,
            I => \c0.n21336\
        );

    \I__5496\ : InMux
    port map (
            O => \N__34198\,
            I => \N__34194\
        );

    \I__5495\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34189\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__34194\,
            I => \N__34186\
        );

    \I__5493\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34183\
        );

    \I__5492\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34180\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__34189\,
            I => \N__34177\
        );

    \I__5490\ : Span4Mux_h
    port map (
            O => \N__34186\,
            I => \N__34172\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__34183\,
            I => \N__34172\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__34180\,
            I => data_in_2_3
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__34177\,
            I => data_in_2_3
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__34172\,
            I => data_in_2_3
        );

    \I__5485\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34161\
        );

    \I__5484\ : InMux
    port map (
            O => \N__34164\,
            I => \N__34158\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__34161\,
            I => \N__34153\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__34158\,
            I => \N__34150\
        );

    \I__5481\ : InMux
    port map (
            O => \N__34157\,
            I => \N__34147\
        );

    \I__5480\ : InMux
    port map (
            O => \N__34156\,
            I => \N__34144\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__34153\,
            I => \N__34141\
        );

    \I__5478\ : Odrv4
    port map (
            O => \N__34150\,
            I => data_in_2_1
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__34147\,
            I => data_in_2_1
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__34144\,
            I => data_in_2_1
        );

    \I__5475\ : Odrv4
    port map (
            O => \N__34141\,
            I => data_in_2_1
        );

    \I__5474\ : CascadeMux
    port map (
            O => \N__34132\,
            I => \c0.n13_adj_4388_cascade_\
        );

    \I__5473\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34126\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__34126\,
            I => \c0.n23135\
        );

    \I__5471\ : InMux
    port map (
            O => \N__34123\,
            I => \N__34120\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__34120\,
            I => \N__34116\
        );

    \I__5469\ : InMux
    port map (
            O => \N__34119\,
            I => \N__34113\
        );

    \I__5468\ : Span4Mux_h
    port map (
            O => \N__34116\,
            I => \N__34110\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__34113\,
            I => \quad_counter0.b_delay_counter_14\
        );

    \I__5466\ : Odrv4
    port map (
            O => \N__34110\,
            I => \quad_counter0.b_delay_counter_14\
        );

    \I__5465\ : InMux
    port map (
            O => \N__34105\,
            I => \N__34102\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__34102\,
            I => \N__34098\
        );

    \I__5463\ : InMux
    port map (
            O => \N__34101\,
            I => \N__34095\
        );

    \I__5462\ : Span4Mux_h
    port map (
            O => \N__34098\,
            I => \N__34092\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__34095\,
            I => \quad_counter0.b_delay_counter_7\
        );

    \I__5460\ : Odrv4
    port map (
            O => \N__34092\,
            I => \quad_counter0.b_delay_counter_7\
        );

    \I__5459\ : CascadeMux
    port map (
            O => \N__34087\,
            I => \N__34084\
        );

    \I__5458\ : InMux
    port map (
            O => \N__34084\,
            I => \N__34081\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__34081\,
            I => \N__34077\
        );

    \I__5456\ : InMux
    port map (
            O => \N__34080\,
            I => \N__34074\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__34077\,
            I => \N__34071\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__34074\,
            I => \quad_counter0.b_delay_counter_12\
        );

    \I__5453\ : Odrv4
    port map (
            O => \N__34071\,
            I => \quad_counter0.b_delay_counter_12\
        );

    \I__5452\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34063\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__34063\,
            I => \N__34059\
        );

    \I__5450\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34056\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__34059\,
            I => \N__34053\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__34056\,
            I => \quad_counter0.b_delay_counter_15\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__34053\,
            I => \quad_counter0.b_delay_counter_15\
        );

    \I__5446\ : InMux
    port map (
            O => \N__34048\,
            I => \N__34045\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__34045\,
            I => \N__34042\
        );

    \I__5444\ : Span4Mux_h
    port map (
            O => \N__34042\,
            I => \N__34039\
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__34039\,
            I => \quad_counter0.n27_adj_4200\
        );

    \I__5442\ : InMux
    port map (
            O => \N__34036\,
            I => \N__34033\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__34033\,
            I => \c0.n14457\
        );

    \I__5440\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34027\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__34027\,
            I => \N__34024\
        );

    \I__5438\ : Span4Mux_v
    port map (
            O => \N__34024\,
            I => \N__34020\
        );

    \I__5437\ : InMux
    port map (
            O => \N__34023\,
            I => \N__34017\
        );

    \I__5436\ : Span4Mux_h
    port map (
            O => \N__34020\,
            I => \N__34014\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__34017\,
            I => data_out_frame_8_0
        );

    \I__5434\ : Odrv4
    port map (
            O => \N__34014\,
            I => data_out_frame_8_0
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__34009\,
            I => \N__34006\
        );

    \I__5432\ : InMux
    port map (
            O => \N__34006\,
            I => \N__34000\
        );

    \I__5431\ : InMux
    port map (
            O => \N__34005\,
            I => \N__34000\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__34000\,
            I => data_out_frame_7_1
        );

    \I__5429\ : InMux
    port map (
            O => \N__33997\,
            I => \N__33994\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__33994\,
            I => \c0.n24093\
        );

    \I__5427\ : CascadeMux
    port map (
            O => \N__33991\,
            I => \c0.n5_adj_4518_cascade_\
        );

    \I__5426\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33985\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__33985\,
            I => \N__33982\
        );

    \I__5424\ : Span4Mux_h
    port map (
            O => \N__33982\,
            I => \N__33979\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__33979\,
            I => \c0.n23862\
        );

    \I__5422\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33972\
        );

    \I__5421\ : CascadeMux
    port map (
            O => \N__33975\,
            I => \N__33960\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__33972\,
            I => \N__33956\
        );

    \I__5419\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33949\
        );

    \I__5418\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33949\
        );

    \I__5417\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33949\
        );

    \I__5416\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33939\
        );

    \I__5415\ : InMux
    port map (
            O => \N__33967\,
            I => \N__33932\
        );

    \I__5414\ : InMux
    port map (
            O => \N__33966\,
            I => \N__33932\
        );

    \I__5413\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33927\
        );

    \I__5412\ : InMux
    port map (
            O => \N__33964\,
            I => \N__33927\
        );

    \I__5411\ : InMux
    port map (
            O => \N__33963\,
            I => \N__33924\
        );

    \I__5410\ : InMux
    port map (
            O => \N__33960\,
            I => \N__33919\
        );

    \I__5409\ : InMux
    port map (
            O => \N__33959\,
            I => \N__33919\
        );

    \I__5408\ : Span4Mux_v
    port map (
            O => \N__33956\,
            I => \N__33914\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__33949\,
            I => \N__33914\
        );

    \I__5406\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33907\
        );

    \I__5405\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33907\
        );

    \I__5404\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33907\
        );

    \I__5403\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33902\
        );

    \I__5402\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33902\
        );

    \I__5401\ : InMux
    port map (
            O => \N__33943\,
            I => \N__33899\
        );

    \I__5400\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33896\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__33939\,
            I => \N__33893\
        );

    \I__5398\ : InMux
    port map (
            O => \N__33938\,
            I => \N__33890\
        );

    \I__5397\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33883\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__33932\,
            I => \N__33870\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__33927\,
            I => \N__33870\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__33924\,
            I => \N__33870\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__33919\,
            I => \N__33870\
        );

    \I__5392\ : Span4Mux_v
    port map (
            O => \N__33914\,
            I => \N__33870\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__33907\,
            I => \N__33870\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__33902\,
            I => \N__33865\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33865\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__33896\,
            I => \N__33858\
        );

    \I__5387\ : Span4Mux_h
    port map (
            O => \N__33893\,
            I => \N__33858\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__33890\,
            I => \N__33855\
        );

    \I__5385\ : InMux
    port map (
            O => \N__33889\,
            I => \N__33845\
        );

    \I__5384\ : InMux
    port map (
            O => \N__33888\,
            I => \N__33845\
        );

    \I__5383\ : InMux
    port map (
            O => \N__33887\,
            I => \N__33845\
        );

    \I__5382\ : InMux
    port map (
            O => \N__33886\,
            I => \N__33845\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__33883\,
            I => \N__33838\
        );

    \I__5380\ : Span4Mux_v
    port map (
            O => \N__33870\,
            I => \N__33838\
        );

    \I__5379\ : Span4Mux_v
    port map (
            O => \N__33865\,
            I => \N__33838\
        );

    \I__5378\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33835\
        );

    \I__5377\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33832\
        );

    \I__5376\ : Span4Mux_h
    port map (
            O => \N__33858\,
            I => \N__33829\
        );

    \I__5375\ : Span4Mux_h
    port map (
            O => \N__33855\,
            I => \N__33826\
        );

    \I__5374\ : InMux
    port map (
            O => \N__33854\,
            I => \N__33823\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__33845\,
            I => \N__33816\
        );

    \I__5372\ : Sp12to4
    port map (
            O => \N__33838\,
            I => \N__33816\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__33835\,
            I => \N__33816\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__33832\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__5369\ : Odrv4
    port map (
            O => \N__33829\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__33826\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__33823\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__5366\ : Odrv12
    port map (
            O => \N__33816\,
            I => \c0.byte_transmit_counter_2\
        );

    \I__5365\ : InMux
    port map (
            O => \N__33805\,
            I => \N__33801\
        );

    \I__5364\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33798\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__33801\,
            I => \N__33795\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__33798\,
            I => data_out_frame_5_7
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__33795\,
            I => data_out_frame_5_7
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__33790\,
            I => \N__33787\
        );

    \I__5359\ : InMux
    port map (
            O => \N__33787\,
            I => \N__33784\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__33784\,
            I => \N__33781\
        );

    \I__5357\ : Span4Mux_h
    port map (
            O => \N__33781\,
            I => \N__33778\
        );

    \I__5356\ : Span4Mux_h
    port map (
            O => \N__33778\,
            I => \N__33775\
        );

    \I__5355\ : Odrv4
    port map (
            O => \N__33775\,
            I => \c0.n24054\
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__33772\,
            I => \N__33764\
        );

    \I__5353\ : CascadeMux
    port map (
            O => \N__33771\,
            I => \N__33760\
        );

    \I__5352\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33757\
        );

    \I__5351\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33749\
        );

    \I__5350\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33749\
        );

    \I__5349\ : InMux
    port map (
            O => \N__33767\,
            I => \N__33749\
        );

    \I__5348\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33744\
        );

    \I__5347\ : InMux
    port map (
            O => \N__33763\,
            I => \N__33744\
        );

    \I__5346\ : InMux
    port map (
            O => \N__33760\,
            I => \N__33741\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__33757\,
            I => \N__33738\
        );

    \I__5344\ : InMux
    port map (
            O => \N__33756\,
            I => \N__33735\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__33749\,
            I => \N__33731\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__33744\,
            I => \N__33722\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__33741\,
            I => \N__33722\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__33738\,
            I => \N__33722\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__33735\,
            I => \N__33722\
        );

    \I__5338\ : InMux
    port map (
            O => \N__33734\,
            I => \N__33719\
        );

    \I__5337\ : Span4Mux_h
    port map (
            O => \N__33731\,
            I => \N__33716\
        );

    \I__5336\ : Span4Mux_h
    port map (
            O => \N__33722\,
            I => \N__33713\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__33719\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__33716\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__33713\,
            I => \c0.tx.r_SM_Main_0\
        );

    \I__5332\ : InMux
    port map (
            O => \N__33706\,
            I => \N__33703\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__33703\,
            I => \N__33700\
        );

    \I__5330\ : Span4Mux_h
    port map (
            O => \N__33700\,
            I => \N__33697\
        );

    \I__5329\ : Odrv4
    port map (
            O => \N__33697\,
            I => \c0.tx.n7086\
        );

    \I__5328\ : CascadeMux
    port map (
            O => \N__33694\,
            I => \N__33673\
        );

    \I__5327\ : CascadeMux
    port map (
            O => \N__33693\,
            I => \N__33669\
        );

    \I__5326\ : CascadeMux
    port map (
            O => \N__33692\,
            I => \N__33665\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__33691\,
            I => \N__33660\
        );

    \I__5324\ : CascadeMux
    port map (
            O => \N__33690\,
            I => \N__33657\
        );

    \I__5323\ : CascadeMux
    port map (
            O => \N__33689\,
            I => \N__33653\
        );

    \I__5322\ : CascadeMux
    port map (
            O => \N__33688\,
            I => \N__33649\
        );

    \I__5321\ : CascadeMux
    port map (
            O => \N__33687\,
            I => \N__33645\
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__33686\,
            I => \N__33641\
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__33685\,
            I => \N__33637\
        );

    \I__5318\ : CascadeMux
    port map (
            O => \N__33684\,
            I => \N__33633\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__33683\,
            I => \N__33629\
        );

    \I__5316\ : CascadeMux
    port map (
            O => \N__33682\,
            I => \N__33625\
        );

    \I__5315\ : CascadeMux
    port map (
            O => \N__33681\,
            I => \N__33622\
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__33680\,
            I => \N__33619\
        );

    \I__5313\ : CascadeMux
    port map (
            O => \N__33679\,
            I => \N__33616\
        );

    \I__5312\ : CascadeMux
    port map (
            O => \N__33678\,
            I => \N__33613\
        );

    \I__5311\ : CascadeMux
    port map (
            O => \N__33677\,
            I => \N__33610\
        );

    \I__5310\ : CascadeMux
    port map (
            O => \N__33676\,
            I => \N__33607\
        );

    \I__5309\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33592\
        );

    \I__5308\ : InMux
    port map (
            O => \N__33672\,
            I => \N__33592\
        );

    \I__5307\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33592\
        );

    \I__5306\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33592\
        );

    \I__5305\ : InMux
    port map (
            O => \N__33665\,
            I => \N__33592\
        );

    \I__5304\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33592\
        );

    \I__5303\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33587\
        );

    \I__5302\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33587\
        );

    \I__5301\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33570\
        );

    \I__5300\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33570\
        );

    \I__5299\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33570\
        );

    \I__5298\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33570\
        );

    \I__5297\ : InMux
    port map (
            O => \N__33649\,
            I => \N__33570\
        );

    \I__5296\ : InMux
    port map (
            O => \N__33648\,
            I => \N__33570\
        );

    \I__5295\ : InMux
    port map (
            O => \N__33645\,
            I => \N__33570\
        );

    \I__5294\ : InMux
    port map (
            O => \N__33644\,
            I => \N__33570\
        );

    \I__5293\ : InMux
    port map (
            O => \N__33641\,
            I => \N__33553\
        );

    \I__5292\ : InMux
    port map (
            O => \N__33640\,
            I => \N__33553\
        );

    \I__5291\ : InMux
    port map (
            O => \N__33637\,
            I => \N__33553\
        );

    \I__5290\ : InMux
    port map (
            O => \N__33636\,
            I => \N__33553\
        );

    \I__5289\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33553\
        );

    \I__5288\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33553\
        );

    \I__5287\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33553\
        );

    \I__5286\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33553\
        );

    \I__5285\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33544\
        );

    \I__5284\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33544\
        );

    \I__5283\ : InMux
    port map (
            O => \N__33619\,
            I => \N__33544\
        );

    \I__5282\ : InMux
    port map (
            O => \N__33616\,
            I => \N__33544\
        );

    \I__5281\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33535\
        );

    \I__5280\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33535\
        );

    \I__5279\ : InMux
    port map (
            O => \N__33607\,
            I => \N__33535\
        );

    \I__5278\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33535\
        );

    \I__5277\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33532\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__33592\,
            I => \N__33527\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__33587\,
            I => \N__33527\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__33570\,
            I => \N__33522\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__33553\,
            I => \N__33522\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__33544\,
            I => \N__33517\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__33535\,
            I => \N__33517\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__33532\,
            I => \N__33514\
        );

    \I__5269\ : Span4Mux_v
    port map (
            O => \N__33527\,
            I => \N__33509\
        );

    \I__5268\ : Span4Mux_v
    port map (
            O => \N__33522\,
            I => \N__33509\
        );

    \I__5267\ : Span4Mux_h
    port map (
            O => \N__33517\,
            I => \N__33506\
        );

    \I__5266\ : Span4Mux_h
    port map (
            O => \N__33514\,
            I => \N__33499\
        );

    \I__5265\ : Span4Mux_h
    port map (
            O => \N__33509\,
            I => \N__33499\
        );

    \I__5264\ : Span4Mux_v
    port map (
            O => \N__33506\,
            I => \N__33499\
        );

    \I__5263\ : Odrv4
    port map (
            O => \N__33499\,
            I => \quad_counter0.n2227\
        );

    \I__5262\ : InMux
    port map (
            O => \N__33496\,
            I => \bfn_14_18_0_\
        );

    \I__5261\ : CascadeMux
    port map (
            O => \N__33493\,
            I => \c0.n14474_cascade_\
        );

    \I__5260\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33484\
        );

    \I__5259\ : InMux
    port map (
            O => \N__33489\,
            I => \N__33484\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__33484\,
            I => data_out_frame_9_1
        );

    \I__5257\ : CascadeMux
    port map (
            O => \N__33481\,
            I => \N__33478\
        );

    \I__5256\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33475\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__33475\,
            I => \N__33471\
        );

    \I__5254\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33468\
        );

    \I__5253\ : Span4Mux_v
    port map (
            O => \N__33471\,
            I => \N__33465\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__33468\,
            I => data_out_frame_8_1
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__33465\,
            I => data_out_frame_8_1
        );

    \I__5250\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33457\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__33457\,
            I => \N__33454\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__33454\,
            I => \N__33451\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__33451\,
            I => \c0.n24186\
        );

    \I__5246\ : InMux
    port map (
            O => \N__33448\,
            I => \N__33445\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__33445\,
            I => n2248
        );

    \I__5244\ : InMux
    port map (
            O => \N__33442\,
            I => \N__33439\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__33439\,
            I => n2240
        );

    \I__5242\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33433\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__33433\,
            I => \N__33429\
        );

    \I__5240\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33426\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__33429\,
            I => \N__33423\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__33426\,
            I => data_out_frame_7_7
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__33423\,
            I => data_out_frame_7_7
        );

    \I__5236\ : CascadeMux
    port map (
            O => \N__33418\,
            I => \N__33415\
        );

    \I__5235\ : InMux
    port map (
            O => \N__33415\,
            I => \N__33409\
        );

    \I__5234\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33409\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__33409\,
            I => data_out_frame_5_1
        );

    \I__5232\ : InMux
    port map (
            O => \N__33406\,
            I => \bfn_14_17_0_\
        );

    \I__5231\ : InMux
    port map (
            O => \N__33403\,
            I => \quad_counter0.n19604\
        );

    \I__5230\ : InMux
    port map (
            O => \N__33400\,
            I => \quad_counter0.n19605\
        );

    \I__5229\ : InMux
    port map (
            O => \N__33397\,
            I => \quad_counter0.n19606\
        );

    \I__5228\ : CascadeMux
    port map (
            O => \N__33394\,
            I => \N__33391\
        );

    \I__5227\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33388\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__33388\,
            I => \N__33383\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__33387\,
            I => \N__33380\
        );

    \I__5224\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33377\
        );

    \I__5223\ : Span4Mux_h
    port map (
            O => \N__33383\,
            I => \N__33373\
        );

    \I__5222\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33370\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__33377\,
            I => \N__33367\
        );

    \I__5220\ : CascadeMux
    port map (
            O => \N__33376\,
            I => \N__33363\
        );

    \I__5219\ : Sp12to4
    port map (
            O => \N__33373\,
            I => \N__33358\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__33370\,
            I => \N__33358\
        );

    \I__5217\ : Span4Mux_h
    port map (
            O => \N__33367\,
            I => \N__33355\
        );

    \I__5216\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33350\
        );

    \I__5215\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33350\
        );

    \I__5214\ : Odrv12
    port map (
            O => \N__33358\,
            I => encoder0_position_27
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__33355\,
            I => encoder0_position_27
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__33350\,
            I => encoder0_position_27
        );

    \I__5211\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33340\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__33340\,
            I => \N__33337\
        );

    \I__5209\ : Odrv12
    port map (
            O => \N__33337\,
            I => n2244
        );

    \I__5208\ : InMux
    port map (
            O => \N__33334\,
            I => \quad_counter0.n19607\
        );

    \I__5207\ : InMux
    port map (
            O => \N__33331\,
            I => \quad_counter0.n19608\
        );

    \I__5206\ : InMux
    port map (
            O => \N__33328\,
            I => \quad_counter0.n19609\
        );

    \I__5205\ : InMux
    port map (
            O => \N__33325\,
            I => \N__33322\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__33322\,
            I => \N__33319\
        );

    \I__5203\ : Span4Mux_v
    port map (
            O => \N__33319\,
            I => \N__33316\
        );

    \I__5202\ : Odrv4
    port map (
            O => \N__33316\,
            I => n2241
        );

    \I__5201\ : InMux
    port map (
            O => \N__33313\,
            I => \quad_counter0.n19610\
        );

    \I__5200\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33307\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__33307\,
            I => \N__33304\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__33304\,
            I => n2257
        );

    \I__5197\ : InMux
    port map (
            O => \N__33301\,
            I => \quad_counter0.n19594\
        );

    \I__5196\ : InMux
    port map (
            O => \N__33298\,
            I => \bfn_14_16_0_\
        );

    \I__5195\ : InMux
    port map (
            O => \N__33295\,
            I => \quad_counter0.n19596\
        );

    \I__5194\ : InMux
    port map (
            O => \N__33292\,
            I => \quad_counter0.n19597\
        );

    \I__5193\ : InMux
    port map (
            O => \N__33289\,
            I => \quad_counter0.n19598\
        );

    \I__5192\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33283\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__33283\,
            I => n2252
        );

    \I__5190\ : InMux
    port map (
            O => \N__33280\,
            I => \quad_counter0.n19599\
        );

    \I__5189\ : InMux
    port map (
            O => \N__33277\,
            I => \N__33274\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__33274\,
            I => \N__33271\
        );

    \I__5187\ : Odrv4
    port map (
            O => \N__33271\,
            I => n2251
        );

    \I__5186\ : InMux
    port map (
            O => \N__33268\,
            I => \quad_counter0.n19600\
        );

    \I__5185\ : InMux
    port map (
            O => \N__33265\,
            I => \quad_counter0.n19601\
        );

    \I__5184\ : InMux
    port map (
            O => \N__33262\,
            I => \quad_counter0.n19602\
        );

    \I__5183\ : InMux
    port map (
            O => \N__33259\,
            I => \quad_counter0.n19585\
        );

    \I__5182\ : InMux
    port map (
            O => \N__33256\,
            I => \quad_counter0.n19586\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__33253\,
            I => \N__33250\
        );

    \I__5180\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33246\
        );

    \I__5179\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33240\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__33246\,
            I => \N__33237\
        );

    \I__5177\ : CascadeMux
    port map (
            O => \N__33245\,
            I => \N__33234\
        );

    \I__5176\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33231\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__33243\,
            I => \N__33227\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__33240\,
            I => \N__33222\
        );

    \I__5173\ : Span4Mux_v
    port map (
            O => \N__33237\,
            I => \N__33222\
        );

    \I__5172\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33219\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__33231\,
            I => \N__33216\
        );

    \I__5170\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33213\
        );

    \I__5169\ : InMux
    port map (
            O => \N__33227\,
            I => \N__33210\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__33222\,
            I => encoder0_position_7
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__33219\,
            I => encoder0_position_7
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__33216\,
            I => encoder0_position_7
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__33213\,
            I => encoder0_position_7
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__33210\,
            I => encoder0_position_7
        );

    \I__5163\ : InMux
    port map (
            O => \N__33199\,
            I => \N__33196\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__33196\,
            I => n2264
        );

    \I__5161\ : InMux
    port map (
            O => \N__33193\,
            I => \bfn_14_15_0_\
        );

    \I__5160\ : InMux
    port map (
            O => \N__33190\,
            I => \quad_counter0.n19588\
        );

    \I__5159\ : InMux
    port map (
            O => \N__33187\,
            I => \quad_counter0.n19589\
        );

    \I__5158\ : InMux
    port map (
            O => \N__33184\,
            I => \quad_counter0.n19590\
        );

    \I__5157\ : InMux
    port map (
            O => \N__33181\,
            I => \quad_counter0.n19591\
        );

    \I__5156\ : InMux
    port map (
            O => \N__33178\,
            I => \quad_counter0.n19592\
        );

    \I__5155\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33172\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__33172\,
            I => \N__33169\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__33169\,
            I => n2258
        );

    \I__5152\ : InMux
    port map (
            O => \N__33166\,
            I => \quad_counter0.n19593\
        );

    \I__5151\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33151\
        );

    \I__5150\ : InMux
    port map (
            O => \N__33162\,
            I => \N__33151\
        );

    \I__5149\ : InMux
    port map (
            O => \N__33161\,
            I => \N__33151\
        );

    \I__5148\ : InMux
    port map (
            O => \N__33160\,
            I => \N__33151\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__33151\,
            I => \N__33148\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__33148\,
            I => \c0.n20160\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__33145\,
            I => \N__33142\
        );

    \I__5144\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33139\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__33139\,
            I => \N__33136\
        );

    \I__5142\ : Span4Mux_v
    port map (
            O => \N__33136\,
            I => \N__33133\
        );

    \I__5141\ : Span4Mux_v
    port map (
            O => \N__33133\,
            I => \N__33130\
        );

    \I__5140\ : Span4Mux_h
    port map (
            O => \N__33130\,
            I => \N__33127\
        );

    \I__5139\ : Odrv4
    port map (
            O => \N__33127\,
            I => \quad_counter0.count_direction\
        );

    \I__5138\ : InMux
    port map (
            O => \N__33124\,
            I => \quad_counter0.n19580\
        );

    \I__5137\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33118\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__33118\,
            I => n2270
        );

    \I__5135\ : InMux
    port map (
            O => \N__33115\,
            I => \quad_counter0.n19581\
        );

    \I__5134\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33109\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__33109\,
            I => n2269
        );

    \I__5132\ : InMux
    port map (
            O => \N__33106\,
            I => \quad_counter0.n19582\
        );

    \I__5131\ : InMux
    port map (
            O => \N__33103\,
            I => \N__33100\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__33100\,
            I => \N__33097\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__33097\,
            I => \N__33094\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__33094\,
            I => n2268
        );

    \I__5127\ : InMux
    port map (
            O => \N__33091\,
            I => \quad_counter0.n19583\
        );

    \I__5126\ : InMux
    port map (
            O => \N__33088\,
            I => \quad_counter0.n19584\
        );

    \I__5125\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33081\
        );

    \I__5124\ : CascadeMux
    port map (
            O => \N__33084\,
            I => \N__33078\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__33081\,
            I => \N__33075\
        );

    \I__5122\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33072\
        );

    \I__5121\ : Span4Mux_h
    port map (
            O => \N__33075\,
            I => \N__33069\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__33072\,
            I => \c0.n21943\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__33069\,
            I => \c0.n21943\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__33064\,
            I => \N__33061\
        );

    \I__5117\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33051\
        );

    \I__5116\ : InMux
    port map (
            O => \N__33060\,
            I => \N__33051\
        );

    \I__5115\ : InMux
    port map (
            O => \N__33059\,
            I => \N__33043\
        );

    \I__5114\ : InMux
    port map (
            O => \N__33058\,
            I => \N__33043\
        );

    \I__5113\ : InMux
    port map (
            O => \N__33057\,
            I => \N__33043\
        );

    \I__5112\ : InMux
    port map (
            O => \N__33056\,
            I => \N__33040\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__33037\
        );

    \I__5110\ : InMux
    port map (
            O => \N__33050\,
            I => \N__33034\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__33043\,
            I => \N__33031\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__33040\,
            I => \c0.n21196\
        );

    \I__5107\ : Odrv12
    port map (
            O => \N__33037\,
            I => \c0.n21196\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__33034\,
            I => \c0.n21196\
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__33031\,
            I => \c0.n21196\
        );

    \I__5104\ : CascadeMux
    port map (
            O => \N__33022\,
            I => \N__33019\
        );

    \I__5103\ : InMux
    port map (
            O => \N__33019\,
            I => \N__33014\
        );

    \I__5102\ : CascadeMux
    port map (
            O => \N__33018\,
            I => \N__33011\
        );

    \I__5101\ : CascadeMux
    port map (
            O => \N__33017\,
            I => \N__33007\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__33014\,
            I => \N__33004\
        );

    \I__5099\ : InMux
    port map (
            O => \N__33011\,
            I => \N__33001\
        );

    \I__5098\ : InMux
    port map (
            O => \N__33010\,
            I => \N__32998\
        );

    \I__5097\ : InMux
    port map (
            O => \N__33007\,
            I => \N__32995\
        );

    \I__5096\ : Span4Mux_h
    port map (
            O => \N__33004\,
            I => \N__32992\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__33001\,
            I => \N__32989\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__32998\,
            I => encoder1_position_25
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__32995\,
            I => encoder1_position_25
        );

    \I__5092\ : Odrv4
    port map (
            O => \N__32992\,
            I => encoder1_position_25
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__32989\,
            I => encoder1_position_25
        );

    \I__5090\ : CascadeMux
    port map (
            O => \N__32980\,
            I => \N__32976\
        );

    \I__5089\ : InMux
    port map (
            O => \N__32979\,
            I => \N__32972\
        );

    \I__5088\ : InMux
    port map (
            O => \N__32976\,
            I => \N__32969\
        );

    \I__5087\ : CascadeMux
    port map (
            O => \N__32975\,
            I => \N__32966\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__32972\,
            I => \N__32962\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__32969\,
            I => \N__32959\
        );

    \I__5084\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32956\
        );

    \I__5083\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32952\
        );

    \I__5082\ : Span4Mux_v
    port map (
            O => \N__32962\,
            I => \N__32945\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__32959\,
            I => \N__32945\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__32956\,
            I => \N__32945\
        );

    \I__5079\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32942\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__32952\,
            I => encoder1_position_11
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__32945\,
            I => encoder1_position_11
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__32942\,
            I => encoder1_position_11
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__32935\,
            I => \c0.n20232_cascade_\
        );

    \I__5074\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32928\
        );

    \I__5073\ : InMux
    port map (
            O => \N__32931\,
            I => \N__32925\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__32928\,
            I => \N__32920\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32920\
        );

    \I__5070\ : Span4Mux_h
    port map (
            O => \N__32920\,
            I => \N__32915\
        );

    \I__5069\ : InMux
    port map (
            O => \N__32919\,
            I => \N__32910\
        );

    \I__5068\ : InMux
    port map (
            O => \N__32918\,
            I => \N__32910\
        );

    \I__5067\ : Odrv4
    port map (
            O => \N__32915\,
            I => \c0.n21146\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__32910\,
            I => \c0.n21146\
        );

    \I__5065\ : CascadeMux
    port map (
            O => \N__32905\,
            I => \c0.n21146_cascade_\
        );

    \I__5064\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32897\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__32901\,
            I => \N__32894\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__32900\,
            I => \N__32889\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__32897\,
            I => \N__32886\
        );

    \I__5060\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32883\
        );

    \I__5059\ : InMux
    port map (
            O => \N__32893\,
            I => \N__32880\
        );

    \I__5058\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32877\
        );

    \I__5057\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32874\
        );

    \I__5056\ : Span4Mux_h
    port map (
            O => \N__32886\,
            I => \N__32871\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__32883\,
            I => \N__32868\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__32880\,
            I => encoder1_position_23
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__32877\,
            I => encoder1_position_23
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__32874\,
            I => encoder1_position_23
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__32871\,
            I => encoder1_position_23
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__32868\,
            I => encoder1_position_23
        );

    \I__5049\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32853\
        );

    \I__5048\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32849\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__32853\,
            I => \N__32846\
        );

    \I__5046\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32842\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__32849\,
            I => \N__32839\
        );

    \I__5044\ : Span4Mux_h
    port map (
            O => \N__32846\,
            I => \N__32836\
        );

    \I__5043\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32833\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__32842\,
            I => \c0.n20232\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__32839\,
            I => \c0.n20232\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__32836\,
            I => \c0.n20232\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__32833\,
            I => \c0.n20232\
        );

    \I__5038\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32820\
        );

    \I__5037\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32817\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__32820\,
            I => \N__32811\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__32817\,
            I => \N__32811\
        );

    \I__5034\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32808\
        );

    \I__5033\ : Span4Mux_h
    port map (
            O => \N__32811\,
            I => \N__32805\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__32808\,
            I => \c0.n20744\
        );

    \I__5031\ : Odrv4
    port map (
            O => \N__32805\,
            I => \c0.n20744\
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__32800\,
            I => \N__32796\
        );

    \I__5029\ : CascadeMux
    port map (
            O => \N__32799\,
            I => \N__32793\
        );

    \I__5028\ : InMux
    port map (
            O => \N__32796\,
            I => \N__32786\
        );

    \I__5027\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32781\
        );

    \I__5026\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32778\
        );

    \I__5025\ : InMux
    port map (
            O => \N__32791\,
            I => \N__32773\
        );

    \I__5024\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32773\
        );

    \I__5023\ : InMux
    port map (
            O => \N__32789\,
            I => \N__32770\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__32786\,
            I => \N__32767\
        );

    \I__5021\ : InMux
    port map (
            O => \N__32785\,
            I => \N__32764\
        );

    \I__5020\ : InMux
    port map (
            O => \N__32784\,
            I => \N__32761\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__32781\,
            I => \N__32758\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__32778\,
            I => \N__32753\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__32773\,
            I => \N__32753\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__32770\,
            I => encoder1_position_1
        );

    \I__5015\ : Odrv12
    port map (
            O => \N__32767\,
            I => encoder1_position_1
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__32764\,
            I => encoder1_position_1
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__32761\,
            I => encoder1_position_1
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__32758\,
            I => encoder1_position_1
        );

    \I__5011\ : Odrv12
    port map (
            O => \N__32753\,
            I => encoder1_position_1
        );

    \I__5010\ : CascadeMux
    port map (
            O => \N__32740\,
            I => \N__32735\
        );

    \I__5009\ : CascadeMux
    port map (
            O => \N__32739\,
            I => \N__32730\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__32738\,
            I => \N__32727\
        );

    \I__5007\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32721\
        );

    \I__5006\ : CascadeMux
    port map (
            O => \N__32734\,
            I => \N__32718\
        );

    \I__5005\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32715\
        );

    \I__5004\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32712\
        );

    \I__5003\ : InMux
    port map (
            O => \N__32727\,
            I => \N__32705\
        );

    \I__5002\ : InMux
    port map (
            O => \N__32726\,
            I => \N__32705\
        );

    \I__5001\ : InMux
    port map (
            O => \N__32725\,
            I => \N__32705\
        );

    \I__5000\ : CascadeMux
    port map (
            O => \N__32724\,
            I => \N__32701\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__32721\,
            I => \N__32697\
        );

    \I__4998\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32694\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__32715\,
            I => \N__32691\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__32712\,
            I => \N__32688\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__32705\,
            I => \N__32685\
        );

    \I__4994\ : InMux
    port map (
            O => \N__32704\,
            I => \N__32680\
        );

    \I__4993\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32680\
        );

    \I__4992\ : InMux
    port map (
            O => \N__32700\,
            I => \N__32677\
        );

    \I__4991\ : Span4Mux_v
    port map (
            O => \N__32697\,
            I => \N__32670\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__32694\,
            I => \N__32670\
        );

    \I__4989\ : Span4Mux_h
    port map (
            O => \N__32691\,
            I => \N__32670\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__32688\,
            I => \N__32667\
        );

    \I__4987\ : Sp12to4
    port map (
            O => \N__32685\,
            I => \N__32662\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__32680\,
            I => \N__32662\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__32677\,
            I => encoder1_position_5
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__32670\,
            I => encoder1_position_5
        );

    \I__4983\ : Odrv4
    port map (
            O => \N__32667\,
            I => encoder1_position_5
        );

    \I__4982\ : Odrv12
    port map (
            O => \N__32662\,
            I => encoder1_position_5
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__32653\,
            I => \c0.n22163_cascade_\
        );

    \I__4980\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32647\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__32647\,
            I => \c0.n20_adj_4505\
        );

    \I__4978\ : CascadeMux
    port map (
            O => \N__32644\,
            I => \c0.n19_adj_4506_cascade_\
        );

    \I__4977\ : InMux
    port map (
            O => \N__32641\,
            I => \N__32638\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__32638\,
            I => \N__32634\
        );

    \I__4975\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32631\
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__32634\,
            I => \c0.n21283\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__32631\,
            I => \c0.n21283\
        );

    \I__4972\ : InMux
    port map (
            O => \N__32626\,
            I => \N__32623\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__32623\,
            I => \N__32620\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__32620\,
            I => \c0.n6_adj_4508\
        );

    \I__4969\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32613\
        );

    \I__4968\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32610\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32607\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__32610\,
            I => \N__32604\
        );

    \I__4965\ : Span4Mux_h
    port map (
            O => \N__32607\,
            I => \N__32601\
        );

    \I__4964\ : Span4Mux_v
    port map (
            O => \N__32604\,
            I => \N__32598\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__32601\,
            I => \c0.n21116\
        );

    \I__4962\ : Odrv4
    port map (
            O => \N__32598\,
            I => \c0.n21116\
        );

    \I__4961\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32589\
        );

    \I__4960\ : InMux
    port map (
            O => \N__32592\,
            I => \N__32586\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__32589\,
            I => \N__32583\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__32586\,
            I => \N__32580\
        );

    \I__4957\ : Span4Mux_h
    port map (
            O => \N__32583\,
            I => \N__32577\
        );

    \I__4956\ : Odrv12
    port map (
            O => \N__32580\,
            I => \c0.n20819\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__32577\,
            I => \c0.n20819\
        );

    \I__4954\ : InMux
    port map (
            O => \N__32572\,
            I => \N__32569\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__32569\,
            I => \c0.n21_adj_4507\
        );

    \I__4952\ : CascadeMux
    port map (
            O => \N__32566\,
            I => \N__32562\
        );

    \I__4951\ : InMux
    port map (
            O => \N__32565\,
            I => \N__32558\
        );

    \I__4950\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32555\
        );

    \I__4949\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32549\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__32558\,
            I => \N__32544\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__32555\,
            I => \N__32544\
        );

    \I__4946\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32541\
        );

    \I__4945\ : InMux
    port map (
            O => \N__32553\,
            I => \N__32538\
        );

    \I__4944\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32535\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__32549\,
            I => \N__32526\
        );

    \I__4942\ : Span4Mux_h
    port map (
            O => \N__32544\,
            I => \N__32526\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__32541\,
            I => \N__32526\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__32538\,
            I => \N__32526\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__32535\,
            I => \N__32521\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__32526\,
            I => \N__32521\
        );

    \I__4937\ : Odrv4
    port map (
            O => \N__32521\,
            I => \c0.n20276\
        );

    \I__4936\ : InMux
    port map (
            O => \N__32518\,
            I => \N__32513\
        );

    \I__4935\ : InMux
    port map (
            O => \N__32517\,
            I => \N__32509\
        );

    \I__4934\ : InMux
    port map (
            O => \N__32516\,
            I => \N__32506\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__32513\,
            I => \N__32502\
        );

    \I__4932\ : InMux
    port map (
            O => \N__32512\,
            I => \N__32499\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__32509\,
            I => \N__32495\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__32506\,
            I => \N__32490\
        );

    \I__4929\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32487\
        );

    \I__4928\ : Span4Mux_v
    port map (
            O => \N__32502\,
            I => \N__32482\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__32499\,
            I => \N__32482\
        );

    \I__4926\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32479\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__32495\,
            I => \N__32476\
        );

    \I__4924\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32473\
        );

    \I__4923\ : InMux
    port map (
            O => \N__32493\,
            I => \N__32470\
        );

    \I__4922\ : Span4Mux_h
    port map (
            O => \N__32490\,
            I => \N__32465\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__32487\,
            I => \N__32465\
        );

    \I__4920\ : Span4Mux_v
    port map (
            O => \N__32482\,
            I => \N__32460\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__32479\,
            I => \N__32460\
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__32476\,
            I => \c0.n21122\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__32473\,
            I => \c0.n21122\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__32470\,
            I => \c0.n21122\
        );

    \I__4915\ : Odrv4
    port map (
            O => \N__32465\,
            I => \c0.n21122\
        );

    \I__4914\ : Odrv4
    port map (
            O => \N__32460\,
            I => \c0.n21122\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__32449\,
            I => \N__32443\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__32448\,
            I => \N__32439\
        );

    \I__4911\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32434\
        );

    \I__4910\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32434\
        );

    \I__4909\ : InMux
    port map (
            O => \N__32443\,
            I => \N__32431\
        );

    \I__4908\ : InMux
    port map (
            O => \N__32442\,
            I => \N__32428\
        );

    \I__4907\ : InMux
    port map (
            O => \N__32439\,
            I => \N__32425\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__32434\,
            I => \N__32422\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__32431\,
            I => \N__32417\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__32428\,
            I => \N__32414\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__32425\,
            I => \N__32411\
        );

    \I__4902\ : Span4Mux_h
    port map (
            O => \N__32422\,
            I => \N__32408\
        );

    \I__4901\ : InMux
    port map (
            O => \N__32421\,
            I => \N__32403\
        );

    \I__4900\ : InMux
    port map (
            O => \N__32420\,
            I => \N__32403\
        );

    \I__4899\ : Span4Mux_v
    port map (
            O => \N__32417\,
            I => \N__32398\
        );

    \I__4898\ : Span4Mux_h
    port map (
            O => \N__32414\,
            I => \N__32398\
        );

    \I__4897\ : Odrv4
    port map (
            O => \N__32411\,
            I => \c0.n21166\
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__32408\,
            I => \c0.n21166\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__32403\,
            I => \c0.n21166\
        );

    \I__4894\ : Odrv4
    port map (
            O => \N__32398\,
            I => \c0.n21166\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__32389\,
            I => \N__32386\
        );

    \I__4892\ : InMux
    port map (
            O => \N__32386\,
            I => \N__32381\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__32385\,
            I => \N__32377\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__32384\,
            I => \N__32374\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__32381\,
            I => \N__32368\
        );

    \I__4888\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32364\
        );

    \I__4887\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32361\
        );

    \I__4886\ : InMux
    port map (
            O => \N__32374\,
            I => \N__32358\
        );

    \I__4885\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32355\
        );

    \I__4884\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32352\
        );

    \I__4883\ : InMux
    port map (
            O => \N__32371\,
            I => \N__32349\
        );

    \I__4882\ : Span4Mux_v
    port map (
            O => \N__32368\,
            I => \N__32346\
        );

    \I__4881\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32343\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__32364\,
            I => \N__32334\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__32361\,
            I => \N__32334\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__32358\,
            I => \N__32334\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__32355\,
            I => \N__32334\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__32352\,
            I => \c0.n13480\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__32349\,
            I => \c0.n13480\
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__32346\,
            I => \c0.n13480\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__32343\,
            I => \c0.n13480\
        );

    \I__4872\ : Odrv4
    port map (
            O => \N__32334\,
            I => \c0.n13480\
        );

    \I__4871\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32320\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__32320\,
            I => \N__32317\
        );

    \I__4869\ : Span4Mux_h
    port map (
            O => \N__32317\,
            I => \N__32314\
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__32314\,
            I => \c0.n22078\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__32311\,
            I => \N__32306\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__32310\,
            I => \N__32303\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__32309\,
            I => \N__32299\
        );

    \I__4864\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32296\
        );

    \I__4863\ : InMux
    port map (
            O => \N__32303\,
            I => \N__32293\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__32302\,
            I => \N__32290\
        );

    \I__4861\ : InMux
    port map (
            O => \N__32299\,
            I => \N__32287\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32283\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__32293\,
            I => \N__32280\
        );

    \I__4858\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32277\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__32287\,
            I => \N__32274\
        );

    \I__4856\ : InMux
    port map (
            O => \N__32286\,
            I => \N__32270\
        );

    \I__4855\ : Span4Mux_v
    port map (
            O => \N__32283\,
            I => \N__32263\
        );

    \I__4854\ : Span4Mux_v
    port map (
            O => \N__32280\,
            I => \N__32263\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__32277\,
            I => \N__32263\
        );

    \I__4852\ : Span4Mux_h
    port map (
            O => \N__32274\,
            I => \N__32260\
        );

    \I__4851\ : InMux
    port map (
            O => \N__32273\,
            I => \N__32257\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__32270\,
            I => encoder1_position_9
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__32263\,
            I => encoder1_position_9
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__32260\,
            I => encoder1_position_9
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__32257\,
            I => encoder1_position_9
        );

    \I__4846\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32242\
        );

    \I__4845\ : InMux
    port map (
            O => \N__32247\,
            I => \N__32237\
        );

    \I__4844\ : InMux
    port map (
            O => \N__32246\,
            I => \N__32237\
        );

    \I__4843\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32234\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32228\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__32237\,
            I => \N__32228\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__32234\,
            I => \N__32225\
        );

    \I__4839\ : InMux
    port map (
            O => \N__32233\,
            I => \N__32222\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__32228\,
            I => \N__32219\
        );

    \I__4837\ : Odrv12
    port map (
            O => \N__32225\,
            I => \c0.n21112\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__32222\,
            I => \c0.n21112\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__32219\,
            I => \c0.n21112\
        );

    \I__4834\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32207\
        );

    \I__4833\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32201\
        );

    \I__4832\ : InMux
    port map (
            O => \N__32210\,
            I => \N__32198\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__32207\,
            I => \N__32195\
        );

    \I__4830\ : InMux
    port map (
            O => \N__32206\,
            I => \N__32190\
        );

    \I__4829\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32190\
        );

    \I__4828\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32187\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__32201\,
            I => \N__32179\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__32198\,
            I => \N__32179\
        );

    \I__4825\ : Span4Mux_h
    port map (
            O => \N__32195\,
            I => \N__32179\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__32190\,
            I => \N__32176\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__32187\,
            I => \N__32173\
        );

    \I__4822\ : InMux
    port map (
            O => \N__32186\,
            I => \N__32170\
        );

    \I__4821\ : Span4Mux_v
    port map (
            O => \N__32179\,
            I => \N__32167\
        );

    \I__4820\ : Span4Mux_h
    port map (
            O => \N__32176\,
            I => \N__32162\
        );

    \I__4819\ : Span4Mux_v
    port map (
            O => \N__32173\,
            I => \N__32162\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__32170\,
            I => \N__32159\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__32167\,
            I => \c0.n21253\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__32162\,
            I => \c0.n21253\
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__32159\,
            I => \c0.n21253\
        );

    \I__4814\ : CascadeMux
    port map (
            O => \N__32152\,
            I => \c0.n20180_cascade_\
        );

    \I__4813\ : InMux
    port map (
            O => \N__32149\,
            I => \N__32145\
        );

    \I__4812\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32142\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__32145\,
            I => \N__32136\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__32142\,
            I => \N__32136\
        );

    \I__4809\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32132\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__32136\,
            I => \N__32129\
        );

    \I__4807\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32126\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__32132\,
            I => \N__32123\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__32129\,
            I => \c0.data_out_frame_29__7__N_1144\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__32126\,
            I => \c0.data_out_frame_29__7__N_1144\
        );

    \I__4803\ : Odrv4
    port map (
            O => \N__32123\,
            I => \c0.data_out_frame_29__7__N_1144\
        );

    \I__4802\ : InMux
    port map (
            O => \N__32116\,
            I => \N__32110\
        );

    \I__4801\ : InMux
    port map (
            O => \N__32115\,
            I => \N__32106\
        );

    \I__4800\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32101\
        );

    \I__4799\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32101\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__32110\,
            I => \N__32097\
        );

    \I__4797\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32094\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__32106\,
            I => \N__32089\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__32101\,
            I => \N__32089\
        );

    \I__4794\ : InMux
    port map (
            O => \N__32100\,
            I => \N__32086\
        );

    \I__4793\ : Span4Mux_v
    port map (
            O => \N__32097\,
            I => \N__32083\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__32094\,
            I => \N__32080\
        );

    \I__4791\ : Span4Mux_h
    port map (
            O => \N__32089\,
            I => \N__32075\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__32086\,
            I => \N__32075\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__32083\,
            I => \c0.n20465\
        );

    \I__4788\ : Odrv12
    port map (
            O => \N__32080\,
            I => \c0.n20465\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__32075\,
            I => \c0.n20465\
        );

    \I__4786\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32065\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__32065\,
            I => \N__32061\
        );

    \I__4784\ : InMux
    port map (
            O => \N__32064\,
            I => \N__32058\
        );

    \I__4783\ : Span4Mux_v
    port map (
            O => \N__32061\,
            I => \N__32055\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__32058\,
            I => data_out_frame_13_7
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__32055\,
            I => data_out_frame_13_7
        );

    \I__4780\ : CascadeMux
    port map (
            O => \N__32050\,
            I => \N__32047\
        );

    \I__4779\ : InMux
    port map (
            O => \N__32047\,
            I => \N__32043\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__32046\,
            I => \N__32040\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__32043\,
            I => \N__32036\
        );

    \I__4776\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32030\
        );

    \I__4775\ : InMux
    port map (
            O => \N__32039\,
            I => \N__32030\
        );

    \I__4774\ : Span4Mux_h
    port map (
            O => \N__32036\,
            I => \N__32027\
        );

    \I__4773\ : InMux
    port map (
            O => \N__32035\,
            I => \N__32024\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__32030\,
            I => \N__32021\
        );

    \I__4771\ : Odrv4
    port map (
            O => \N__32027\,
            I => \c0.n21056\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__32024\,
            I => \c0.n21056\
        );

    \I__4769\ : Odrv4
    port map (
            O => \N__32021\,
            I => \c0.n21056\
        );

    \I__4768\ : InMux
    port map (
            O => \N__32014\,
            I => \N__32010\
        );

    \I__4767\ : InMux
    port map (
            O => \N__32013\,
            I => \N__32007\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__32010\,
            I => \c0.n22177\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__32007\,
            I => \c0.n22177\
        );

    \I__4764\ : InMux
    port map (
            O => \N__32002\,
            I => \N__31999\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__31999\,
            I => \c0.n22072\
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__31996\,
            I => \c0.n22072_cascade_\
        );

    \I__4761\ : InMux
    port map (
            O => \N__31993\,
            I => \N__31990\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__31990\,
            I => \N__31985\
        );

    \I__4759\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31982\
        );

    \I__4758\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31979\
        );

    \I__4757\ : Span4Mux_h
    port map (
            O => \N__31985\,
            I => \N__31974\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31974\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__31979\,
            I => \c0.n22073\
        );

    \I__4754\ : Odrv4
    port map (
            O => \N__31974\,
            I => \c0.n22073\
        );

    \I__4753\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31965\
        );

    \I__4752\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31961\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__31965\,
            I => \N__31958\
        );

    \I__4750\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31953\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__31961\,
            I => \N__31948\
        );

    \I__4748\ : Span4Mux_v
    port map (
            O => \N__31958\,
            I => \N__31948\
        );

    \I__4747\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31943\
        );

    \I__4746\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31943\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__31953\,
            I => \N__31940\
        );

    \I__4744\ : Span4Mux_v
    port map (
            O => \N__31948\,
            I => \N__31935\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__31943\,
            I => \N__31935\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__31940\,
            I => \c0.n20175\
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__31935\,
            I => \c0.n20175\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__31930\,
            I => \c0.n20249_cascade_\
        );

    \I__4739\ : InMux
    port map (
            O => \N__31927\,
            I => \N__31923\
        );

    \I__4738\ : InMux
    port map (
            O => \N__31926\,
            I => \N__31919\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__31923\,
            I => \N__31916\
        );

    \I__4736\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31913\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__31919\,
            I => \N__31909\
        );

    \I__4734\ : Span4Mux_v
    port map (
            O => \N__31916\,
            I => \N__31904\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__31913\,
            I => \N__31904\
        );

    \I__4732\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31901\
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__31909\,
            I => \c0.n12528\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__31904\,
            I => \c0.n12528\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__31901\,
            I => \c0.n12528\
        );

    \I__4728\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31887\
        );

    \I__4727\ : InMux
    port map (
            O => \N__31893\,
            I => \N__31887\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__31892\,
            I => \N__31883\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__31887\,
            I => \N__31878\
        );

    \I__4724\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31872\
        );

    \I__4723\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31872\
        );

    \I__4722\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31867\
        );

    \I__4721\ : InMux
    port map (
            O => \N__31881\,
            I => \N__31867\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__31878\,
            I => \N__31864\
        );

    \I__4719\ : InMux
    port map (
            O => \N__31877\,
            I => \N__31861\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__31872\,
            I => \c0.n21065\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__31867\,
            I => \c0.n21065\
        );

    \I__4716\ : Odrv4
    port map (
            O => \N__31864\,
            I => \c0.n21065\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__31861\,
            I => \c0.n21065\
        );

    \I__4714\ : InMux
    port map (
            O => \N__31852\,
            I => \N__31849\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__31849\,
            I => \N__31846\
        );

    \I__4712\ : Span4Mux_h
    port map (
            O => \N__31846\,
            I => \N__31843\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__31843\,
            I => \c0.n21842\
        );

    \I__4710\ : InMux
    port map (
            O => \N__31840\,
            I => \N__31835\
        );

    \I__4709\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31832\
        );

    \I__4708\ : CascadeMux
    port map (
            O => \N__31838\,
            I => \N__31829\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__31835\,
            I => \N__31824\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__31832\,
            I => \N__31824\
        );

    \I__4705\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31821\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__31824\,
            I => \N__31818\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__31821\,
            I => \c0.n20230\
        );

    \I__4702\ : Odrv4
    port map (
            O => \N__31818\,
            I => \c0.n20230\
        );

    \I__4701\ : InMux
    port map (
            O => \N__31813\,
            I => \N__31810\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__31810\,
            I => \N__31807\
        );

    \I__4699\ : Span12Mux_v
    port map (
            O => \N__31807\,
            I => \N__31804\
        );

    \I__4698\ : Odrv12
    port map (
            O => \N__31804\,
            I => \c0.n6_adj_4394\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__31801\,
            I => \c0.n6_adj_4497_cascade_\
        );

    \I__4696\ : InMux
    port map (
            O => \N__31798\,
            I => \N__31794\
        );

    \I__4695\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31791\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__31794\,
            I => \N__31788\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__31791\,
            I => \N__31785\
        );

    \I__4692\ : Span4Mux_h
    port map (
            O => \N__31788\,
            I => \N__31782\
        );

    \I__4691\ : Odrv4
    port map (
            O => \N__31785\,
            I => \c0.n20151\
        );

    \I__4690\ : Odrv4
    port map (
            O => \N__31782\,
            I => \c0.n20151\
        );

    \I__4689\ : InMux
    port map (
            O => \N__31777\,
            I => \N__31774\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__31774\,
            I => \c0.data_out_frame_29_6\
        );

    \I__4687\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31767\
        );

    \I__4686\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31764\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__31767\,
            I => \N__31761\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__31764\,
            I => \N__31758\
        );

    \I__4683\ : Span4Mux_h
    port map (
            O => \N__31761\,
            I => \N__31754\
        );

    \I__4682\ : Span4Mux_v
    port map (
            O => \N__31758\,
            I => \N__31751\
        );

    \I__4681\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31748\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__31754\,
            I => \c0.n21848\
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__31751\,
            I => \c0.n21848\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__31748\,
            I => \c0.n21848\
        );

    \I__4677\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31738\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__31738\,
            I => \N__31735\
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__31735\,
            I => \c0.n20253\
        );

    \I__4674\ : CascadeMux
    port map (
            O => \N__31732\,
            I => \c0.n21852_cascade_\
        );

    \I__4673\ : InMux
    port map (
            O => \N__31729\,
            I => \N__31723\
        );

    \I__4672\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31723\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__31723\,
            I => \c0.n22346\
        );

    \I__4670\ : InMux
    port map (
            O => \N__31720\,
            I => \N__31714\
        );

    \I__4669\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31714\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__31714\,
            I => \N__31711\
        );

    \I__4667\ : Odrv12
    port map (
            O => \N__31711\,
            I => \c0.n22126\
        );

    \I__4666\ : InMux
    port map (
            O => \N__31708\,
            I => \N__31704\
        );

    \I__4665\ : InMux
    port map (
            O => \N__31707\,
            I => \N__31701\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__31704\,
            I => \c0.n20298\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__31701\,
            I => \c0.n20298\
        );

    \I__4662\ : CascadeMux
    port map (
            O => \N__31696\,
            I => \c0.n10_adj_4512_cascade_\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__31693\,
            I => \N__31689\
        );

    \I__4660\ : InMux
    port map (
            O => \N__31692\,
            I => \N__31684\
        );

    \I__4659\ : InMux
    port map (
            O => \N__31689\,
            I => \N__31679\
        );

    \I__4658\ : InMux
    port map (
            O => \N__31688\,
            I => \N__31676\
        );

    \I__4657\ : InMux
    port map (
            O => \N__31687\,
            I => \N__31673\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__31684\,
            I => \N__31670\
        );

    \I__4655\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31667\
        );

    \I__4654\ : InMux
    port map (
            O => \N__31682\,
            I => \N__31664\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__31679\,
            I => \N__31657\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__31676\,
            I => \N__31657\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__31673\,
            I => \N__31657\
        );

    \I__4650\ : Span4Mux_v
    port map (
            O => \N__31670\,
            I => \N__31653\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__31667\,
            I => \N__31646\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__31664\,
            I => \N__31646\
        );

    \I__4647\ : Span4Mux_h
    port map (
            O => \N__31657\,
            I => \N__31646\
        );

    \I__4646\ : InMux
    port map (
            O => \N__31656\,
            I => \N__31643\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__31653\,
            I => \c0.n10496\
        );

    \I__4644\ : Odrv4
    port map (
            O => \N__31646\,
            I => \c0.n10496\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__31643\,
            I => \c0.n10496\
        );

    \I__4642\ : InMux
    port map (
            O => \N__31636\,
            I => \N__31627\
        );

    \I__4641\ : InMux
    port map (
            O => \N__31635\,
            I => \N__31624\
        );

    \I__4640\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31618\
        );

    \I__4639\ : InMux
    port map (
            O => \N__31633\,
            I => \N__31618\
        );

    \I__4638\ : InMux
    port map (
            O => \N__31632\,
            I => \N__31613\
        );

    \I__4637\ : InMux
    port map (
            O => \N__31631\,
            I => \N__31613\
        );

    \I__4636\ : InMux
    port map (
            O => \N__31630\,
            I => \N__31610\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__31627\,
            I => \N__31607\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__31624\,
            I => \N__31604\
        );

    \I__4633\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31601\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__31618\,
            I => \N__31594\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__31613\,
            I => \N__31594\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__31610\,
            I => \N__31594\
        );

    \I__4629\ : Span4Mux_h
    port map (
            O => \N__31607\,
            I => \N__31587\
        );

    \I__4628\ : Span4Mux_v
    port map (
            O => \N__31604\,
            I => \N__31587\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__31601\,
            I => \N__31587\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__31594\,
            I => \c0.n20274\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__31587\,
            I => \c0.n20274\
        );

    \I__4624\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31579\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__31579\,
            I => \N__31576\
        );

    \I__4622\ : Span4Mux_v
    port map (
            O => \N__31576\,
            I => \N__31573\
        );

    \I__4621\ : Odrv4
    port map (
            O => \N__31573\,
            I => \c0.n21231\
        );

    \I__4620\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31566\
        );

    \I__4619\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31562\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__31566\,
            I => \N__31558\
        );

    \I__4617\ : InMux
    port map (
            O => \N__31565\,
            I => \N__31555\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__31562\,
            I => \N__31552\
        );

    \I__4615\ : InMux
    port map (
            O => \N__31561\,
            I => \N__31549\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__31558\,
            I => \c0.n22736\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__31555\,
            I => \c0.n22736\
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__31552\,
            I => \c0.n22736\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__31549\,
            I => \c0.n22736\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__31540\,
            I => \c0.n21162_cascade_\
        );

    \I__4609\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31531\
        );

    \I__4608\ : InMux
    port map (
            O => \N__31536\,
            I => \N__31531\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__31531\,
            I => \c0.n12526\
        );

    \I__4606\ : InMux
    port map (
            O => \N__31528\,
            I => \N__31522\
        );

    \I__4605\ : InMux
    port map (
            O => \N__31527\,
            I => \N__31522\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__31522\,
            I => \c0.n20201\
        );

    \I__4603\ : CascadeMux
    port map (
            O => \N__31519\,
            I => \N__31516\
        );

    \I__4602\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31510\
        );

    \I__4601\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31510\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__31510\,
            I => \N__31507\
        );

    \I__4599\ : Odrv4
    port map (
            O => \N__31507\,
            I => \c0.n21876\
        );

    \I__4598\ : CascadeMux
    port map (
            O => \N__31504\,
            I => \N__31501\
        );

    \I__4597\ : InMux
    port map (
            O => \N__31501\,
            I => \N__31498\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__31498\,
            I => \N__31495\
        );

    \I__4595\ : Span4Mux_v
    port map (
            O => \N__31495\,
            I => \N__31492\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__31492\,
            I => \c0.n24119\
        );

    \I__4593\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31486\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__31486\,
            I => \N__31482\
        );

    \I__4591\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31479\
        );

    \I__4590\ : Span4Mux_h
    port map (
            O => \N__31482\,
            I => \N__31476\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__31479\,
            I => \N__31473\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__31476\,
            I => \c0.n21050\
        );

    \I__4587\ : Odrv12
    port map (
            O => \N__31473\,
            I => \c0.n21050\
        );

    \I__4586\ : InMux
    port map (
            O => \N__31468\,
            I => \N__31465\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__31465\,
            I => \c0.n6_adj_4402\
        );

    \I__4584\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31459\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__31459\,
            I => \N__31454\
        );

    \I__4582\ : InMux
    port map (
            O => \N__31458\,
            I => \N__31451\
        );

    \I__4581\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31448\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__31454\,
            I => \c0.n22188\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__31451\,
            I => \c0.n22188\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__31448\,
            I => \c0.n22188\
        );

    \I__4577\ : CascadeMux
    port map (
            O => \N__31441\,
            I => \c0.n20658_cascade_\
        );

    \I__4576\ : InMux
    port map (
            O => \N__31438\,
            I => \N__31435\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__31435\,
            I => \N__31431\
        );

    \I__4574\ : InMux
    port map (
            O => \N__31434\,
            I => \N__31428\
        );

    \I__4573\ : Span4Mux_h
    port map (
            O => \N__31431\,
            I => \N__31425\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__31428\,
            I => \c0.n22166\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__31425\,
            I => \c0.n22166\
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__31420\,
            I => \N__31412\
        );

    \I__4569\ : CascadeMux
    port map (
            O => \N__31419\,
            I => \N__31409\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__31418\,
            I => \N__31406\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__31417\,
            I => \N__31401\
        );

    \I__4566\ : CascadeMux
    port map (
            O => \N__31416\,
            I => \N__31398\
        );

    \I__4565\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31391\
        );

    \I__4564\ : InMux
    port map (
            O => \N__31412\,
            I => \N__31391\
        );

    \I__4563\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31391\
        );

    \I__4562\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31386\
        );

    \I__4561\ : InMux
    port map (
            O => \N__31405\,
            I => \N__31386\
        );

    \I__4560\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31383\
        );

    \I__4559\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31378\
        );

    \I__4558\ : InMux
    port map (
            O => \N__31398\,
            I => \N__31378\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__31391\,
            I => \N__31374\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__31386\,
            I => \N__31367\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__31383\,
            I => \N__31367\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__31378\,
            I => \N__31367\
        );

    \I__4553\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31364\
        );

    \I__4552\ : Span12Mux_h
    port map (
            O => \N__31374\,
            I => \N__31361\
        );

    \I__4551\ : Span4Mux_v
    port map (
            O => \N__31367\,
            I => \N__31358\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__31364\,
            I => \c0.n10467\
        );

    \I__4549\ : Odrv12
    port map (
            O => \N__31361\,
            I => \c0.n10467\
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__31358\,
            I => \c0.n10467\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__31351\,
            I => \N__31345\
        );

    \I__4546\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31342\
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__31349\,
            I => \N__31338\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__31348\,
            I => \N__31334\
        );

    \I__4543\ : InMux
    port map (
            O => \N__31345\,
            I => \N__31331\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__31342\,
            I => \N__31328\
        );

    \I__4541\ : InMux
    port map (
            O => \N__31341\,
            I => \N__31325\
        );

    \I__4540\ : InMux
    port map (
            O => \N__31338\,
            I => \N__31322\
        );

    \I__4539\ : InMux
    port map (
            O => \N__31337\,
            I => \N__31319\
        );

    \I__4538\ : InMux
    port map (
            O => \N__31334\,
            I => \N__31316\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__31331\,
            I => \N__31313\
        );

    \I__4536\ : Span4Mux_v
    port map (
            O => \N__31328\,
            I => \N__31310\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__31325\,
            I => \c0.n22180\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__31322\,
            I => \c0.n22180\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__31319\,
            I => \c0.n22180\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__31316\,
            I => \c0.n22180\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__31313\,
            I => \c0.n22180\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__31310\,
            I => \c0.n22180\
        );

    \I__4529\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31289\
        );

    \I__4528\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31289\
        );

    \I__4527\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31286\
        );

    \I__4526\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31282\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__31289\,
            I => \N__31277\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__31286\,
            I => \N__31277\
        );

    \I__4523\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31274\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__31282\,
            I => \N__31269\
        );

    \I__4521\ : Span4Mux_v
    port map (
            O => \N__31277\,
            I => \N__31266\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__31274\,
            I => \N__31263\
        );

    \I__4519\ : InMux
    port map (
            O => \N__31273\,
            I => \N__31258\
        );

    \I__4518\ : InMux
    port map (
            O => \N__31272\,
            I => \N__31258\
        );

    \I__4517\ : Span4Mux_h
    port map (
            O => \N__31269\,
            I => \N__31253\
        );

    \I__4516\ : Span4Mux_v
    port map (
            O => \N__31266\,
            I => \N__31249\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__31263\,
            I => \N__31244\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__31258\,
            I => \N__31244\
        );

    \I__4513\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31241\
        );

    \I__4512\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31238\
        );

    \I__4511\ : Span4Mux_v
    port map (
            O => \N__31253\,
            I => \N__31235\
        );

    \I__4510\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31232\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__31249\,
            I => \c0.n20330\
        );

    \I__4508\ : Odrv4
    port map (
            O => \N__31244\,
            I => \c0.n20330\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__31241\,
            I => \c0.n20330\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__31238\,
            I => \c0.n20330\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__31235\,
            I => \c0.n20330\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__31232\,
            I => \c0.n20330\
        );

    \I__4503\ : CascadeMux
    port map (
            O => \N__31219\,
            I => \N__31214\
        );

    \I__4502\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31210\
        );

    \I__4501\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31203\
        );

    \I__4500\ : InMux
    port map (
            O => \N__31214\,
            I => \N__31203\
        );

    \I__4499\ : InMux
    port map (
            O => \N__31213\,
            I => \N__31200\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__31210\,
            I => \N__31197\
        );

    \I__4497\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31194\
        );

    \I__4496\ : InMux
    port map (
            O => \N__31208\,
            I => \N__31191\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__31203\,
            I => \N__31185\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31185\
        );

    \I__4493\ : Span4Mux_v
    port map (
            O => \N__31197\,
            I => \N__31182\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31177\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__31191\,
            I => \N__31177\
        );

    \I__4490\ : InMux
    port map (
            O => \N__31190\,
            I => \N__31174\
        );

    \I__4489\ : Span4Mux_h
    port map (
            O => \N__31185\,
            I => \N__31171\
        );

    \I__4488\ : Span4Mux_h
    port map (
            O => \N__31182\,
            I => \N__31166\
        );

    \I__4487\ : Span4Mux_v
    port map (
            O => \N__31177\,
            I => \N__31166\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__31174\,
            I => \c0.n10434\
        );

    \I__4485\ : Odrv4
    port map (
            O => \N__31171\,
            I => \c0.n10434\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__31166\,
            I => \c0.n10434\
        );

    \I__4483\ : InMux
    port map (
            O => \N__31159\,
            I => \N__31153\
        );

    \I__4482\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31153\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__31153\,
            I => \N__31148\
        );

    \I__4480\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31145\
        );

    \I__4479\ : InMux
    port map (
            O => \N__31151\,
            I => \N__31142\
        );

    \I__4478\ : Span4Mux_h
    port map (
            O => \N__31148\,
            I => \N__31139\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__31145\,
            I => \c0.n10513\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__31142\,
            I => \c0.n10513\
        );

    \I__4475\ : Odrv4
    port map (
            O => \N__31139\,
            I => \c0.n10513\
        );

    \I__4474\ : InMux
    port map (
            O => \N__31132\,
            I => \N__31123\
        );

    \I__4473\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31123\
        );

    \I__4472\ : InMux
    port map (
            O => \N__31130\,
            I => \N__31120\
        );

    \I__4471\ : InMux
    port map (
            O => \N__31129\,
            I => \N__31115\
        );

    \I__4470\ : InMux
    port map (
            O => \N__31128\,
            I => \N__31115\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__31123\,
            I => \N__31110\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__31120\,
            I => \N__31110\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__31115\,
            I => \N__31107\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__31110\,
            I => \c0.n21189\
        );

    \I__4465\ : Odrv4
    port map (
            O => \N__31107\,
            I => \c0.n21189\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__31102\,
            I => \N__31099\
        );

    \I__4463\ : InMux
    port map (
            O => \N__31099\,
            I => \N__31096\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__31096\,
            I => \c0.n21135\
        );

    \I__4461\ : InMux
    port map (
            O => \N__31093\,
            I => \N__31090\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__31090\,
            I => \N__31085\
        );

    \I__4459\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31082\
        );

    \I__4458\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31079\
        );

    \I__4457\ : Odrv12
    port map (
            O => \N__31085\,
            I => \c0.n21219\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__31082\,
            I => \c0.n21219\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__31079\,
            I => \c0.n21219\
        );

    \I__4454\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31067\
        );

    \I__4453\ : InMux
    port map (
            O => \N__31071\,
            I => \N__31064\
        );

    \I__4452\ : InMux
    port map (
            O => \N__31070\,
            I => \N__31061\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__31067\,
            I => \c0.n21811\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__31064\,
            I => \c0.n21811\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__31061\,
            I => \c0.n21811\
        );

    \I__4448\ : CascadeMux
    port map (
            O => \N__31054\,
            I => \c0.n21135_cascade_\
        );

    \I__4447\ : InMux
    port map (
            O => \N__31051\,
            I => \c0.tx.n19545\
        );

    \I__4446\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31044\
        );

    \I__4445\ : InMux
    port map (
            O => \N__31047\,
            I => \N__31039\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__31044\,
            I => \N__31036\
        );

    \I__4443\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31031\
        );

    \I__4442\ : InMux
    port map (
            O => \N__31042\,
            I => \N__31031\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__31039\,
            I => \r_Clock_Count_7\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__31036\,
            I => \r_Clock_Count_7\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__31031\,
            I => \r_Clock_Count_7\
        );

    \I__4438\ : InMux
    port map (
            O => \N__31024\,
            I => \N__31021\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__31021\,
            I => \N__31018\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__31018\,
            I => n314
        );

    \I__4435\ : InMux
    port map (
            O => \N__31015\,
            I => \c0.tx.n19546\
        );

    \I__4434\ : InMux
    port map (
            O => \N__31012\,
            I => \bfn_13_22_0_\
        );

    \I__4433\ : InMux
    port map (
            O => \N__31009\,
            I => \N__31006\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__31006\,
            I => \c0.n12878\
        );

    \I__4431\ : SRMux
    port map (
            O => \N__31003\,
            I => \N__31000\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__31000\,
            I => \N__30997\
        );

    \I__4429\ : Span4Mux_h
    port map (
            O => \N__30997\,
            I => \N__30994\
        );

    \I__4428\ : Span4Mux_h
    port map (
            O => \N__30994\,
            I => \N__30991\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__30991\,
            I => \c0.n21360\
        );

    \I__4426\ : SRMux
    port map (
            O => \N__30988\,
            I => \N__30985\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__30985\,
            I => \c0.n21356\
        );

    \I__4424\ : InMux
    port map (
            O => \N__30982\,
            I => \N__30978\
        );

    \I__4423\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30975\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__30978\,
            I => \N__30972\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__30975\,
            I => \c0.n22317\
        );

    \I__4420\ : Odrv4
    port map (
            O => \N__30972\,
            I => \c0.n22317\
        );

    \I__4419\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30964\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__30964\,
            I => \c0.n6_adj_4305\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__30961\,
            I => \c0.tx.n6_cascade_\
        );

    \I__4416\ : InMux
    port map (
            O => \N__30958\,
            I => \N__30955\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__30955\,
            I => \c0.tx.n31\
        );

    \I__4414\ : CascadeMux
    port map (
            O => \N__30952\,
            I => \c0.tx.n31_cascade_\
        );

    \I__4413\ : InMux
    port map (
            O => \N__30949\,
            I => \N__30946\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__30946\,
            I => \c0.tx.n47\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__30943\,
            I => \N__30940\
        );

    \I__4410\ : InMux
    port map (
            O => \N__30940\,
            I => \N__30937\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__30937\,
            I => \c0.tx.n10\
        );

    \I__4408\ : InMux
    port map (
            O => \N__30934\,
            I => \N__30930\
        );

    \I__4407\ : InMux
    port map (
            O => \N__30933\,
            I => \N__30926\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__30930\,
            I => \N__30923\
        );

    \I__4405\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30920\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__30926\,
            I => \N__30915\
        );

    \I__4403\ : Span4Mux_v
    port map (
            O => \N__30923\,
            I => \N__30915\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__30920\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__4401\ : Odrv4
    port map (
            O => \N__30915\,
            I => \c0.tx.r_Clock_Count_0\
        );

    \I__4400\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30907\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__30907\,
            I => \N__30904\
        );

    \I__4398\ : Odrv12
    port map (
            O => \N__30904\,
            I => \c0.tx.n23960\
        );

    \I__4397\ : InMux
    port map (
            O => \N__30901\,
            I => \bfn_13_21_0_\
        );

    \I__4396\ : InMux
    port map (
            O => \N__30898\,
            I => \N__30893\
        );

    \I__4395\ : InMux
    port map (
            O => \N__30897\,
            I => \N__30890\
        );

    \I__4394\ : InMux
    port map (
            O => \N__30896\,
            I => \N__30887\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__30893\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__30890\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__30887\,
            I => \c0.tx.r_Clock_Count_1\
        );

    \I__4390\ : InMux
    port map (
            O => \N__30880\,
            I => \N__30877\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__30877\,
            I => \c0.tx.n23961\
        );

    \I__4388\ : InMux
    port map (
            O => \N__30874\,
            I => \c0.tx.n19540\
        );

    \I__4387\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30866\
        );

    \I__4386\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30863\
        );

    \I__4385\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30860\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__30866\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__30863\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__30860\,
            I => \c0.tx.r_Clock_Count_2\
        );

    \I__4381\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30850\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__30850\,
            I => \c0.tx.n23958\
        );

    \I__4379\ : InMux
    port map (
            O => \N__30847\,
            I => \c0.tx.n19541\
        );

    \I__4378\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30839\
        );

    \I__4377\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30836\
        );

    \I__4376\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30833\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__30839\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__30836\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__30833\,
            I => \c0.tx.r_Clock_Count_3\
        );

    \I__4372\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30823\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__30823\,
            I => \c0.tx.n23963\
        );

    \I__4370\ : InMux
    port map (
            O => \N__30820\,
            I => \c0.tx.n19542\
        );

    \I__4369\ : InMux
    port map (
            O => \N__30817\,
            I => \N__30813\
        );

    \I__4368\ : InMux
    port map (
            O => \N__30816\,
            I => \N__30810\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__30813\,
            I => \N__30804\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__30810\,
            I => \N__30804\
        );

    \I__4365\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30801\
        );

    \I__4364\ : Span4Mux_v
    port map (
            O => \N__30804\,
            I => \N__30798\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__30801\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__30798\,
            I => \c0.tx.r_Clock_Count_4\
        );

    \I__4361\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30790\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__30790\,
            I => \N__30787\
        );

    \I__4359\ : Odrv12
    port map (
            O => \N__30787\,
            I => \c0.tx.n23953\
        );

    \I__4358\ : InMux
    port map (
            O => \N__30784\,
            I => \c0.tx.n19543\
        );

    \I__4357\ : InMux
    port map (
            O => \N__30781\,
            I => \N__30775\
        );

    \I__4356\ : InMux
    port map (
            O => \N__30780\,
            I => \N__30772\
        );

    \I__4355\ : InMux
    port map (
            O => \N__30779\,
            I => \N__30767\
        );

    \I__4354\ : InMux
    port map (
            O => \N__30778\,
            I => \N__30767\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__30775\,
            I => \r_Clock_Count_5\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__30772\,
            I => \r_Clock_Count_5\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__30767\,
            I => \r_Clock_Count_5\
        );

    \I__4350\ : InMux
    port map (
            O => \N__30760\,
            I => \N__30757\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__30757\,
            I => n316
        );

    \I__4348\ : InMux
    port map (
            O => \N__30754\,
            I => \c0.tx.n19544\
        );

    \I__4347\ : CascadeMux
    port map (
            O => \N__30751\,
            I => \o_Tx_Serial_N_3783_cascade_\
        );

    \I__4346\ : InMux
    port map (
            O => \N__30748\,
            I => \N__30745\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__30745\,
            I => \N__30742\
        );

    \I__4344\ : Span4Mux_v
    port map (
            O => \N__30742\,
            I => \N__30739\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__30739\,
            I => \c0.tx.n12\
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__30736\,
            I => \N__30732\
        );

    \I__4341\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30722\
        );

    \I__4340\ : InMux
    port map (
            O => \N__30732\,
            I => \N__30722\
        );

    \I__4339\ : InMux
    port map (
            O => \N__30731\,
            I => \N__30722\
        );

    \I__4338\ : InMux
    port map (
            O => \N__30730\,
            I => \N__30715\
        );

    \I__4337\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30715\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__30722\,
            I => \N__30712\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__30721\,
            I => \N__30708\
        );

    \I__4334\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30700\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__30715\,
            I => \N__30697\
        );

    \I__4332\ : Span4Mux_h
    port map (
            O => \N__30712\,
            I => \N__30694\
        );

    \I__4331\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30691\
        );

    \I__4330\ : InMux
    port map (
            O => \N__30708\,
            I => \N__30684\
        );

    \I__4329\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30684\
        );

    \I__4328\ : InMux
    port map (
            O => \N__30706\,
            I => \N__30684\
        );

    \I__4327\ : InMux
    port map (
            O => \N__30705\,
            I => \N__30677\
        );

    \I__4326\ : InMux
    port map (
            O => \N__30704\,
            I => \N__30677\
        );

    \I__4325\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30677\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__30700\,
            I => \r_SM_Main_1_adj_4550\
        );

    \I__4323\ : Odrv12
    port map (
            O => \N__30697\,
            I => \r_SM_Main_1_adj_4550\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__30694\,
            I => \r_SM_Main_1_adj_4550\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__30691\,
            I => \r_SM_Main_1_adj_4550\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__30684\,
            I => \r_SM_Main_1_adj_4550\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__30677\,
            I => \r_SM_Main_1_adj_4550\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__30664\,
            I => \c0.tx.n6_adj_4214_cascade_\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__30661\,
            I => \N__30657\
        );

    \I__4316\ : InMux
    port map (
            O => \N__30660\,
            I => \N__30654\
        );

    \I__4315\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30651\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__30654\,
            I => \N__30645\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__30651\,
            I => \N__30645\
        );

    \I__4312\ : InMux
    port map (
            O => \N__30650\,
            I => \N__30639\
        );

    \I__4311\ : Span4Mux_h
    port map (
            O => \N__30645\,
            I => \N__30636\
        );

    \I__4310\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30629\
        );

    \I__4309\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30629\
        );

    \I__4308\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30629\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__30639\,
            I => \c0.tx.n16630\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__30636\,
            I => \c0.tx.n16630\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__30629\,
            I => \c0.tx.n16630\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__30622\,
            I => \n8_cascade_\
        );

    \I__4303\ : InMux
    port map (
            O => \N__30619\,
            I => \N__30615\
        );

    \I__4302\ : InMux
    port map (
            O => \N__30618\,
            I => \N__30612\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__30615\,
            I => \N__30608\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__30612\,
            I => \N__30605\
        );

    \I__4299\ : InMux
    port map (
            O => \N__30611\,
            I => \N__30602\
        );

    \I__4298\ : Span12Mux_h
    port map (
            O => \N__30608\,
            I => \N__30597\
        );

    \I__4297\ : Sp12to4
    port map (
            O => \N__30605\,
            I => \N__30597\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__30602\,
            I => data_in_0_2
        );

    \I__4295\ : Odrv12
    port map (
            O => \N__30597\,
            I => data_in_0_2
        );

    \I__4294\ : InMux
    port map (
            O => \N__30592\,
            I => \N__30588\
        );

    \I__4293\ : InMux
    port map (
            O => \N__30591\,
            I => \N__30585\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__30588\,
            I => \c0.n13006\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__30585\,
            I => \c0.n13006\
        );

    \I__4290\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30576\
        );

    \I__4289\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30573\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__30576\,
            I => \c0.n21767\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__30573\,
            I => \c0.n21767\
        );

    \I__4286\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30565\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__30565\,
            I => \N__30562\
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__30562\,
            I => \c0.tx.n14296\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__30559\,
            I => \N__30554\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__30558\,
            I => \N__30551\
        );

    \I__4281\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30547\
        );

    \I__4280\ : InMux
    port map (
            O => \N__30554\,
            I => \N__30544\
        );

    \I__4279\ : InMux
    port map (
            O => \N__30551\,
            I => \N__30541\
        );

    \I__4278\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30538\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__30547\,
            I => \N__30535\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__30544\,
            I => data_in_1_0
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__30541\,
            I => data_in_1_0
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__30538\,
            I => data_in_1_0
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__30535\,
            I => data_in_1_0
        );

    \I__4272\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30522\
        );

    \I__4271\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30519\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__30522\,
            I => data_in_0_0
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__30519\,
            I => data_in_0_0
        );

    \I__4268\ : CascadeMux
    port map (
            O => \N__30514\,
            I => \N__30510\
        );

    \I__4267\ : InMux
    port map (
            O => \N__30513\,
            I => \N__30505\
        );

    \I__4266\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30505\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__30505\,
            I => data_in_0_4
        );

    \I__4264\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30499\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__30499\,
            I => \N__30495\
        );

    \I__4262\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30491\
        );

    \I__4261\ : Span4Mux_v
    port map (
            O => \N__30495\,
            I => \N__30488\
        );

    \I__4260\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30485\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__30491\,
            I => data_in_1_7
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__30488\,
            I => data_in_1_7
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__30485\,
            I => data_in_1_7
        );

    \I__4256\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30475\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__30475\,
            I => \c0.n10_adj_4494\
        );

    \I__4254\ : CascadeMux
    port map (
            O => \N__30472\,
            I => \N__30469\
        );

    \I__4253\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30466\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__30466\,
            I => \N__30463\
        );

    \I__4251\ : Odrv4
    port map (
            O => \N__30463\,
            I => \c0.n16_adj_4476\
        );

    \I__4250\ : InMux
    port map (
            O => \N__30460\,
            I => \N__30457\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__30457\,
            I => \c0.n17_adj_4477\
        );

    \I__4248\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30447\
        );

    \I__4247\ : CascadeMux
    port map (
            O => \N__30453\,
            I => \N__30444\
        );

    \I__4246\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30436\
        );

    \I__4245\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30436\
        );

    \I__4244\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30436\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__30447\,
            I => \N__30433\
        );

    \I__4242\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30427\
        );

    \I__4241\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30427\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__30436\,
            I => \N__30424\
        );

    \I__4239\ : Span4Mux_h
    port map (
            O => \N__30433\,
            I => \N__30421\
        );

    \I__4238\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30418\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__30427\,
            I => \r_Bit_Index_0_adj_4553\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__30424\,
            I => \r_Bit_Index_0_adj_4553\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__30421\,
            I => \r_Bit_Index_0_adj_4553\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__30418\,
            I => \r_Bit_Index_0_adj_4553\
        );

    \I__4233\ : InMux
    port map (
            O => \N__30409\,
            I => \N__30406\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__30406\,
            I => \N__30403\
        );

    \I__4231\ : Odrv4
    port map (
            O => \N__30403\,
            I => n24192
        );

    \I__4230\ : InMux
    port map (
            O => \N__30400\,
            I => \N__30397\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30394\
        );

    \I__4228\ : Span4Mux_h
    port map (
            O => \N__30394\,
            I => \N__30391\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__30391\,
            I => n24198
        );

    \I__4226\ : InMux
    port map (
            O => \N__30388\,
            I => \N__30385\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__30385\,
            I => \N__30381\
        );

    \I__4224\ : InMux
    port map (
            O => \N__30384\,
            I => \N__30378\
        );

    \I__4223\ : Span4Mux_h
    port map (
            O => \N__30381\,
            I => \N__30375\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__30378\,
            I => data_out_frame_6_4
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__30375\,
            I => data_out_frame_6_4
        );

    \I__4220\ : InMux
    port map (
            O => \N__30370\,
            I => \N__30367\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__30367\,
            I => \N__30363\
        );

    \I__4218\ : InMux
    port map (
            O => \N__30366\,
            I => \N__30360\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__30363\,
            I => \c0.n13003\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__30360\,
            I => \c0.n13003\
        );

    \I__4215\ : InMux
    port map (
            O => \N__30355\,
            I => \N__30352\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__30352\,
            I => \c0.n19_adj_4367\
        );

    \I__4213\ : CascadeMux
    port map (
            O => \N__30349\,
            I => \c0.n20_adj_4362_cascade_\
        );

    \I__4212\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30343\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__30343\,
            I => \c0.n23834\
        );

    \I__4210\ : InMux
    port map (
            O => \N__30340\,
            I => \N__30335\
        );

    \I__4209\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30332\
        );

    \I__4208\ : InMux
    port map (
            O => \N__30338\,
            I => \N__30329\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__30335\,
            I => \N__30325\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__30332\,
            I => \N__30322\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__30329\,
            I => \N__30319\
        );

    \I__4204\ : InMux
    port map (
            O => \N__30328\,
            I => \N__30316\
        );

    \I__4203\ : Span4Mux_v
    port map (
            O => \N__30325\,
            I => \N__30313\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__30322\,
            I => \N__30310\
        );

    \I__4201\ : Odrv12
    port map (
            O => \N__30319\,
            I => data_in_1_2
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__30316\,
            I => data_in_1_2
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__30313\,
            I => data_in_1_2
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__30310\,
            I => data_in_1_2
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__30301\,
            I => \N__30296\
        );

    \I__4196\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30293\
        );

    \I__4195\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30288\
        );

    \I__4194\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30288\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__30293\,
            I => data_in_0_5
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__30288\,
            I => data_in_0_5
        );

    \I__4191\ : InMux
    port map (
            O => \N__30283\,
            I => \N__30280\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__30280\,
            I => \N__30274\
        );

    \I__4189\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30269\
        );

    \I__4188\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30269\
        );

    \I__4187\ : InMux
    port map (
            O => \N__30277\,
            I => \N__30266\
        );

    \I__4186\ : Odrv12
    port map (
            O => \N__30274\,
            I => data_in_1_6
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__30269\,
            I => data_in_1_6
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__30266\,
            I => data_in_1_6
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__30259\,
            I => \c0.n17_adj_4479_cascade_\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__30256\,
            I => \N__30253\
        );

    \I__4181\ : InMux
    port map (
            O => \N__30253\,
            I => \N__30249\
        );

    \I__4180\ : InMux
    port map (
            O => \N__30252\,
            I => \N__30246\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__30249\,
            I => \c0.n13023\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__30246\,
            I => \c0.n13023\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__30241\,
            I => \c0.n21914_cascade_\
        );

    \I__4176\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30235\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__30235\,
            I => \c0.n21_adj_4320\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__30232\,
            I => \N__30228\
        );

    \I__4173\ : InMux
    port map (
            O => \N__30231\,
            I => \N__30225\
        );

    \I__4172\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30222\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__30225\,
            I => \N__30219\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__30222\,
            I => data_out_frame_8_4
        );

    \I__4169\ : Odrv12
    port map (
            O => \N__30219\,
            I => data_out_frame_8_4
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__30214\,
            I => \N__30211\
        );

    \I__4167\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30208\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__30208\,
            I => \N__30205\
        );

    \I__4165\ : Span4Mux_h
    port map (
            O => \N__30205\,
            I => \N__30202\
        );

    \I__4164\ : Span4Mux_h
    port map (
            O => \N__30202\,
            I => \N__30199\
        );

    \I__4163\ : Odrv4
    port map (
            O => \N__30199\,
            I => \c0.n23880\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__4161\ : InMux
    port map (
            O => \N__30193\,
            I => \N__30187\
        );

    \I__4160\ : InMux
    port map (
            O => \N__30192\,
            I => \N__30187\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__30187\,
            I => data_out_frame_9_4
        );

    \I__4158\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30181\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__30181\,
            I => \N__30178\
        );

    \I__4156\ : Odrv4
    port map (
            O => \N__30178\,
            I => n2178
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__30175\,
            I => \N__30172\
        );

    \I__4154\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30168\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__30171\,
            I => \N__30165\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__30168\,
            I => \N__30160\
        );

    \I__4151\ : InMux
    port map (
            O => \N__30165\,
            I => \N__30157\
        );

    \I__4150\ : InMux
    port map (
            O => \N__30164\,
            I => \N__30154\
        );

    \I__4149\ : InMux
    port map (
            O => \N__30163\,
            I => \N__30151\
        );

    \I__4148\ : Span4Mux_h
    port map (
            O => \N__30160\,
            I => \N__30148\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__30157\,
            I => \N__30145\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__30154\,
            I => \N__30142\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__30151\,
            I => encoder1_position_27
        );

    \I__4144\ : Odrv4
    port map (
            O => \N__30148\,
            I => encoder1_position_27
        );

    \I__4143\ : Odrv12
    port map (
            O => \N__30145\,
            I => encoder1_position_27
        );

    \I__4142\ : Odrv12
    port map (
            O => \N__30142\,
            I => encoder1_position_27
        );

    \I__4141\ : InMux
    port map (
            O => \N__30133\,
            I => \N__30130\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__30130\,
            I => \N__30126\
        );

    \I__4139\ : InMux
    port map (
            O => \N__30129\,
            I => \N__30123\
        );

    \I__4138\ : Span4Mux_v
    port map (
            O => \N__30126\,
            I => \N__30120\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__30123\,
            I => data_out_frame_10_2
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__30120\,
            I => data_out_frame_10_2
        );

    \I__4135\ : InMux
    port map (
            O => \N__30115\,
            I => \N__30112\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__30112\,
            I => \N__30108\
        );

    \I__4133\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30105\
        );

    \I__4132\ : Span4Mux_v
    port map (
            O => \N__30108\,
            I => \N__30102\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__30105\,
            I => data_out_frame_5_4
        );

    \I__4130\ : Odrv4
    port map (
            O => \N__30102\,
            I => data_out_frame_5_4
        );

    \I__4129\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30094\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__30094\,
            I => \N__30091\
        );

    \I__4127\ : Sp12to4
    port map (
            O => \N__30091\,
            I => \N__30088\
        );

    \I__4126\ : Span12Mux_v
    port map (
            O => \N__30088\,
            I => \N__30085\
        );

    \I__4125\ : Odrv12
    port map (
            O => \N__30085\,
            I => \c0.n11\
        );

    \I__4124\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30079\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__30079\,
            I => \N__30076\
        );

    \I__4122\ : Odrv12
    port map (
            O => \N__30076\,
            I => \c0.n14_adj_4329\
        );

    \I__4121\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30070\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__30070\,
            I => \N__30067\
        );

    \I__4119\ : Span4Mux_h
    port map (
            O => \N__30067\,
            I => \N__30064\
        );

    \I__4118\ : Odrv4
    port map (
            O => \N__30064\,
            I => n2198
        );

    \I__4117\ : InMux
    port map (
            O => \N__30061\,
            I => \N__30058\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__30058\,
            I => \N__30055\
        );

    \I__4115\ : Span4Mux_h
    port map (
            O => \N__30055\,
            I => \N__30052\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__30052\,
            I => n2192
        );

    \I__4113\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30046\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__30046\,
            I => \N__30043\
        );

    \I__4111\ : Span4Mux_v
    port map (
            O => \N__30043\,
            I => \N__30040\
        );

    \I__4110\ : Sp12to4
    port map (
            O => \N__30040\,
            I => \N__30037\
        );

    \I__4109\ : Odrv12
    port map (
            O => \N__30037\,
            I => n2186
        );

    \I__4108\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30031\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__30031\,
            I => \N__30026\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__30030\,
            I => \N__30022\
        );

    \I__4105\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30019\
        );

    \I__4104\ : Span4Mux_v
    port map (
            O => \N__30026\,
            I => \N__30016\
        );

    \I__4103\ : InMux
    port map (
            O => \N__30025\,
            I => \N__30011\
        );

    \I__4102\ : InMux
    port map (
            O => \N__30022\,
            I => \N__30011\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__30019\,
            I => encoder1_position_19
        );

    \I__4100\ : Odrv4
    port map (
            O => \N__30016\,
            I => encoder1_position_19
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__30011\,
            I => encoder1_position_19
        );

    \I__4098\ : InMux
    port map (
            O => \N__30004\,
            I => \N__30001\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__30001\,
            I => \c0.n19_adj_4319\
        );

    \I__4096\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29995\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__29995\,
            I => \c0.n23557\
        );

    \I__4094\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29989\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__29989\,
            I => \N__29986\
        );

    \I__4092\ : Span4Mux_h
    port map (
            O => \N__29986\,
            I => \N__29983\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__29983\,
            I => n2180
        );

    \I__4090\ : InMux
    port map (
            O => \N__29980\,
            I => \N__29968\
        );

    \I__4089\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29968\
        );

    \I__4088\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29968\
        );

    \I__4087\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29968\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__29968\,
            I => \c0.n20767\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__29965\,
            I => \c0.n20767_cascade_\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__29962\,
            I => \N__29959\
        );

    \I__4083\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29954\
        );

    \I__4082\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29951\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__29957\,
            I => \N__29948\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__29954\,
            I => \N__29944\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__29951\,
            I => \N__29941\
        );

    \I__4078\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29938\
        );

    \I__4077\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29934\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__29944\,
            I => \N__29929\
        );

    \I__4075\ : Span4Mux_h
    port map (
            O => \N__29941\,
            I => \N__29929\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__29938\,
            I => \N__29926\
        );

    \I__4073\ : InMux
    port map (
            O => \N__29937\,
            I => \N__29923\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__29934\,
            I => encoder1_position_24
        );

    \I__4071\ : Odrv4
    port map (
            O => \N__29929\,
            I => encoder1_position_24
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__29926\,
            I => encoder1_position_24
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__29923\,
            I => encoder1_position_24
        );

    \I__4068\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29911\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__29911\,
            I => \N__29908\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__29908\,
            I => \N__29905\
        );

    \I__4065\ : Odrv4
    port map (
            O => \N__29905\,
            I => n2195
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__29902\,
            I => \N__29899\
        );

    \I__4063\ : InMux
    port map (
            O => \N__29899\,
            I => \N__29895\
        );

    \I__4062\ : InMux
    port map (
            O => \N__29898\,
            I => \N__29892\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__29895\,
            I => data_out_frame_9_6
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__29892\,
            I => data_out_frame_9_6
        );

    \I__4059\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29884\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__29884\,
            I => \N__29880\
        );

    \I__4057\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29877\
        );

    \I__4056\ : Span4Mux_h
    port map (
            O => \N__29880\,
            I => \N__29874\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__29877\,
            I => \N__29869\
        );

    \I__4054\ : Span4Mux_h
    port map (
            O => \N__29874\,
            I => \N__29869\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__29869\,
            I => data_out_frame_13_6
        );

    \I__4052\ : InMux
    port map (
            O => \N__29866\,
            I => \N__29863\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__29863\,
            I => \N__29860\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__29860\,
            I => \N__29857\
        );

    \I__4049\ : Odrv4
    port map (
            O => \N__29857\,
            I => n2194
        );

    \I__4048\ : InMux
    port map (
            O => \N__29854\,
            I => \N__29847\
        );

    \I__4047\ : InMux
    port map (
            O => \N__29853\,
            I => \N__29844\
        );

    \I__4046\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29837\
        );

    \I__4045\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29837\
        );

    \I__4044\ : InMux
    port map (
            O => \N__29850\,
            I => \N__29837\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__29847\,
            I => \c0.n21175\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__29844\,
            I => \c0.n21175\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__29837\,
            I => \c0.n21175\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__29830\,
            I => \N__29826\
        );

    \I__4039\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29821\
        );

    \I__4038\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29816\
        );

    \I__4037\ : InMux
    port map (
            O => \N__29825\,
            I => \N__29816\
        );

    \I__4036\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29813\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__29821\,
            I => \c0.n21156\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__29816\,
            I => \c0.n21156\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__29813\,
            I => \c0.n21156\
        );

    \I__4032\ : InMux
    port map (
            O => \N__29806\,
            I => \N__29801\
        );

    \I__4031\ : InMux
    port map (
            O => \N__29805\,
            I => \N__29796\
        );

    \I__4030\ : InMux
    port map (
            O => \N__29804\,
            I => \N__29796\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__29801\,
            I => \N__29791\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__29796\,
            I => \N__29791\
        );

    \I__4027\ : Odrv4
    port map (
            O => \N__29791\,
            I => \c0.n12554\
        );

    \I__4026\ : InMux
    port map (
            O => \N__29788\,
            I => \N__29785\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__29785\,
            I => \N__29782\
        );

    \I__4024\ : Span4Mux_h
    port map (
            O => \N__29782\,
            I => \N__29777\
        );

    \I__4023\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29772\
        );

    \I__4022\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29772\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__29777\,
            I => \c0.n20931\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__29772\,
            I => \c0.n20931\
        );

    \I__4019\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29761\
        );

    \I__4018\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29758\
        );

    \I__4017\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29753\
        );

    \I__4016\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29753\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__29761\,
            I => \c0.n22991\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__29758\,
            I => \c0.n22991\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__29753\,
            I => \c0.n22991\
        );

    \I__4012\ : CascadeMux
    port map (
            O => \N__29746\,
            I => \c0.n21189_cascade_\
        );

    \I__4011\ : InMux
    port map (
            O => \N__29743\,
            I => \N__29739\
        );

    \I__4010\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29736\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__29739\,
            I => \N__29733\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__29736\,
            I => \c0.n21058\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__29733\,
            I => \c0.n21058\
        );

    \I__4006\ : InMux
    port map (
            O => \N__29728\,
            I => \N__29722\
        );

    \I__4005\ : InMux
    port map (
            O => \N__29727\,
            I => \N__29722\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29718\
        );

    \I__4003\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29715\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__29718\,
            I => \c0.n21192\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__29715\,
            I => \c0.n21192\
        );

    \I__4000\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29707\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__29707\,
            I => \N__29702\
        );

    \I__3998\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29699\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__29705\,
            I => \N__29696\
        );

    \I__3996\ : Span4Mux_v
    port map (
            O => \N__29702\,
            I => \N__29692\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__29699\,
            I => \N__29689\
        );

    \I__3994\ : InMux
    port map (
            O => \N__29696\,
            I => \N__29684\
        );

    \I__3993\ : InMux
    port map (
            O => \N__29695\,
            I => \N__29684\
        );

    \I__3992\ : Span4Mux_v
    port map (
            O => \N__29692\,
            I => \N__29679\
        );

    \I__3991\ : Span4Mux_v
    port map (
            O => \N__29689\,
            I => \N__29679\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__29684\,
            I => \N__29676\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__29679\,
            I => \c0.n13349\
        );

    \I__3988\ : Odrv12
    port map (
            O => \N__29676\,
            I => \c0.n13349\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__29671\,
            I => \c0.n13480_cascade_\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__29668\,
            I => \c0.n21122_cascade_\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__29665\,
            I => \N__29661\
        );

    \I__3984\ : InMux
    port map (
            O => \N__29664\,
            I => \N__29656\
        );

    \I__3983\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29652\
        );

    \I__3982\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29647\
        );

    \I__3981\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29647\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__29656\,
            I => \N__29644\
        );

    \I__3979\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29641\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__29652\,
            I => \N__29636\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__29647\,
            I => \N__29631\
        );

    \I__3976\ : Span4Mux_v
    port map (
            O => \N__29644\,
            I => \N__29631\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__29641\,
            I => \N__29628\
        );

    \I__3974\ : InMux
    port map (
            O => \N__29640\,
            I => \N__29623\
        );

    \I__3973\ : InMux
    port map (
            O => \N__29639\,
            I => \N__29623\
        );

    \I__3972\ : Span4Mux_v
    port map (
            O => \N__29636\,
            I => \N__29618\
        );

    \I__3971\ : Span4Mux_h
    port map (
            O => \N__29631\,
            I => \N__29618\
        );

    \I__3970\ : Odrv4
    port map (
            O => \N__29628\,
            I => encoder1_position_14
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__29623\,
            I => encoder1_position_14
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__29618\,
            I => encoder1_position_14
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__29611\,
            I => \c0.n6_adj_4509_cascade_\
        );

    \I__3966\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29605\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__29605\,
            I => \c0.n22393\
        );

    \I__3964\ : InMux
    port map (
            O => \N__29602\,
            I => \N__29597\
        );

    \I__3963\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29594\
        );

    \I__3962\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29591\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__29597\,
            I => \c0.n10498\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__29594\,
            I => \c0.n10498\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__29591\,
            I => \c0.n10498\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__29584\,
            I => \c0.n22393_cascade_\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__29581\,
            I => \c0.n14_adj_4510_cascade_\
        );

    \I__3956\ : InMux
    port map (
            O => \N__29578\,
            I => \N__29570\
        );

    \I__3955\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29570\
        );

    \I__3954\ : InMux
    port map (
            O => \N__29576\,
            I => \N__29565\
        );

    \I__3953\ : InMux
    port map (
            O => \N__29575\,
            I => \N__29565\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__29570\,
            I => \N__29559\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__29565\,
            I => \N__29556\
        );

    \I__3950\ : InMux
    port map (
            O => \N__29564\,
            I => \N__29553\
        );

    \I__3949\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29550\
        );

    \I__3948\ : InMux
    port map (
            O => \N__29562\,
            I => \N__29547\
        );

    \I__3947\ : Span4Mux_h
    port map (
            O => \N__29559\,
            I => \N__29544\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__29556\,
            I => \N__29537\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__29553\,
            I => \N__29537\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__29550\,
            I => \N__29537\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__29547\,
            I => \c0.n10462\
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__29544\,
            I => \c0.n10462\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__29537\,
            I => \c0.n10462\
        );

    \I__3940\ : InMux
    port map (
            O => \N__29530\,
            I => \N__29524\
        );

    \I__3939\ : InMux
    port map (
            O => \N__29529\,
            I => \N__29524\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29521\
        );

    \I__3937\ : Span4Mux_h
    port map (
            O => \N__29521\,
            I => \N__29517\
        );

    \I__3936\ : InMux
    port map (
            O => \N__29520\,
            I => \N__29514\
        );

    \I__3935\ : Odrv4
    port map (
            O => \N__29517\,
            I => \c0.n21150\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__29514\,
            I => \c0.n21150\
        );

    \I__3933\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29506\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__29506\,
            I => \c0.n10_adj_4511\
        );

    \I__3931\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29500\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__29500\,
            I => \c0.n10_adj_4330\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__29497\,
            I => \c0.n21192_cascade_\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__29494\,
            I => \c0.n20931_cascade_\
        );

    \I__3927\ : InMux
    port map (
            O => \N__29491\,
            I => \N__29488\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__29488\,
            I => \c0.n22151\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__29485\,
            I => \c0.n22151_cascade_\
        );

    \I__3924\ : CascadeMux
    port map (
            O => \N__29482\,
            I => \c0.n6_adj_4397_cascade_\
        );

    \I__3923\ : InMux
    port map (
            O => \N__29479\,
            I => \N__29476\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__29476\,
            I => \c0.data_out_frame_28_0\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__29473\,
            I => \N__29470\
        );

    \I__3920\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29467\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__29467\,
            I => \N__29463\
        );

    \I__3918\ : InMux
    port map (
            O => \N__29466\,
            I => \N__29460\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__29463\,
            I => \c0.n22018\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__29460\,
            I => \c0.n22018\
        );

    \I__3915\ : InMux
    port map (
            O => \N__29455\,
            I => \N__29452\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__29452\,
            I => \c0.data_out_frame_29_5\
        );

    \I__3913\ : InMux
    port map (
            O => \N__29449\,
            I => \N__29446\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__29446\,
            I => \c0.data_out_frame_28_5\
        );

    \I__3911\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29440\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29437\
        );

    \I__3909\ : Span4Mux_h
    port map (
            O => \N__29437\,
            I => \N__29434\
        );

    \I__3908\ : Sp12to4
    port map (
            O => \N__29434\,
            I => \N__29431\
        );

    \I__3907\ : Span12Mux_v
    port map (
            O => \N__29431\,
            I => \N__29428\
        );

    \I__3906\ : Odrv12
    port map (
            O => \N__29428\,
            I => \c0.n26_adj_4347\
        );

    \I__3905\ : InMux
    port map (
            O => \N__29425\,
            I => \N__29420\
        );

    \I__3904\ : InMux
    port map (
            O => \N__29424\,
            I => \N__29417\
        );

    \I__3903\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29413\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29408\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__29417\,
            I => \N__29405\
        );

    \I__3900\ : InMux
    port map (
            O => \N__29416\,
            I => \N__29402\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__29413\,
            I => \N__29399\
        );

    \I__3898\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29394\
        );

    \I__3897\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29394\
        );

    \I__3896\ : Span4Mux_v
    port map (
            O => \N__29408\,
            I => \N__29389\
        );

    \I__3895\ : Span4Mux_v
    port map (
            O => \N__29405\,
            I => \N__29389\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__29402\,
            I => \c0.n20376\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__29399\,
            I => \c0.n20376\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__29394\,
            I => \c0.n20376\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__29389\,
            I => \c0.n20376\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__29380\,
            I => \c0.n22018_cascade_\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__29377\,
            I => \N__29374\
        );

    \I__3888\ : InMux
    port map (
            O => \N__29374\,
            I => \N__29371\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__29371\,
            I => \N__29368\
        );

    \I__3886\ : Span4Mux_h
    port map (
            O => \N__29368\,
            I => \N__29365\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__29365\,
            I => \c0.n21946\
        );

    \I__3884\ : CascadeMux
    port map (
            O => \N__29362\,
            I => \c0.n21946_cascade_\
        );

    \I__3883\ : InMux
    port map (
            O => \N__29359\,
            I => \N__29355\
        );

    \I__3882\ : InMux
    port map (
            O => \N__29358\,
            I => \N__29350\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__29355\,
            I => \N__29347\
        );

    \I__3880\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29344\
        );

    \I__3879\ : InMux
    port map (
            O => \N__29353\,
            I => \N__29341\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__29350\,
            I => \N__29338\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__29347\,
            I => \N__29335\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__29344\,
            I => \N__29332\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__29341\,
            I => \N__29327\
        );

    \I__3874\ : Span4Mux_h
    port map (
            O => \N__29338\,
            I => \N__29327\
        );

    \I__3873\ : Odrv4
    port map (
            O => \N__29335\,
            I => \c0.n12532\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__29332\,
            I => \c0.n12532\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__29327\,
            I => \c0.n12532\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__29320\,
            I => \c0.n12491_cascade_\
        );

    \I__3869\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29314\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__29314\,
            I => \c0.data_out_frame_28_6\
        );

    \I__3867\ : InMux
    port map (
            O => \N__29311\,
            I => \N__29308\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__29308\,
            I => \N__29305\
        );

    \I__3865\ : Span4Mux_v
    port map (
            O => \N__29305\,
            I => \N__29302\
        );

    \I__3864\ : Span4Mux_v
    port map (
            O => \N__29302\,
            I => \N__29299\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__29299\,
            I => \c0.n26_adj_4351\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__29296\,
            I => \c0.n7_adj_4307_cascade_\
        );

    \I__3861\ : InMux
    port map (
            O => \N__29293\,
            I => \N__29289\
        );

    \I__3860\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29286\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__29289\,
            I => \N__29283\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__29286\,
            I => \N__29280\
        );

    \I__3857\ : Span4Mux_h
    port map (
            O => \N__29283\,
            I => \N__29277\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__29280\,
            I => \data_out_frame_29__3__N_1662\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__29277\,
            I => \data_out_frame_29__3__N_1662\
        );

    \I__3854\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29267\
        );

    \I__3853\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29264\
        );

    \I__3852\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29261\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__29267\,
            I => \c0.n22024\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__29264\,
            I => \c0.n22024\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__29261\,
            I => \c0.n22024\
        );

    \I__3848\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29251\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29248\
        );

    \I__3846\ : Odrv12
    port map (
            O => \N__29248\,
            I => \c0.data_out_frame_29_4\
        );

    \I__3845\ : SRMux
    port map (
            O => \N__29245\,
            I => \N__29242\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__29242\,
            I => \N__29239\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__29239\,
            I => \N__29236\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__29236\,
            I => \c0.n21376\
        );

    \I__3841\ : SRMux
    port map (
            O => \N__29233\,
            I => \N__29230\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__29230\,
            I => \c0.n21362\
        );

    \I__3839\ : CascadeMux
    port map (
            O => \N__29227\,
            I => \N__29224\
        );

    \I__3838\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29221\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__29221\,
            I => \N__29218\
        );

    \I__3836\ : Odrv4
    port map (
            O => \N__29218\,
            I => \c0.n21128\
        );

    \I__3835\ : InMux
    port map (
            O => \N__29215\,
            I => \N__29212\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__29212\,
            I => \c0.n12_adj_4516\
        );

    \I__3833\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29206\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__29206\,
            I => \c0.n9_adj_4339\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__29203\,
            I => \c0.tx.n16631_cascade_\
        );

    \I__3830\ : InMux
    port map (
            O => \N__29200\,
            I => \N__29194\
        );

    \I__3829\ : InMux
    port map (
            O => \N__29199\,
            I => \N__29194\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__29194\,
            I => \N__29189\
        );

    \I__3827\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29186\
        );

    \I__3826\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29183\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__29189\,
            I => \N__29180\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__29186\,
            I => n14442
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__29183\,
            I => n14442
        );

    \I__3822\ : Odrv4
    port map (
            O => \N__29180\,
            I => n14442
        );

    \I__3821\ : SRMux
    port map (
            O => \N__29173\,
            I => \N__29170\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__29170\,
            I => \N__29167\
        );

    \I__3819\ : Odrv4
    port map (
            O => \N__29167\,
            I => \c0.n21370\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__29164\,
            I => \c0.n10_adj_4231_cascade_\
        );

    \I__3817\ : InMux
    port map (
            O => \N__29161\,
            I => \N__29158\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__29158\,
            I => \c0.n14\
        );

    \I__3815\ : InMux
    port map (
            O => \N__29155\,
            I => \N__29149\
        );

    \I__3814\ : InMux
    port map (
            O => \N__29154\,
            I => \N__29146\
        );

    \I__3813\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29139\
        );

    \I__3812\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29139\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__29149\,
            I => \N__29136\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__29146\,
            I => \N__29132\
        );

    \I__3809\ : InMux
    port map (
            O => \N__29145\,
            I => \N__29127\
        );

    \I__3808\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29127\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__29139\,
            I => \N__29124\
        );

    \I__3806\ : Span4Mux_v
    port map (
            O => \N__29136\,
            I => \N__29121\
        );

    \I__3805\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29118\
        );

    \I__3804\ : Span12Mux_s11_h
    port map (
            O => \N__29132\,
            I => \N__29114\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__29127\,
            I => \N__29111\
        );

    \I__3802\ : Span4Mux_h
    port map (
            O => \N__29124\,
            I => \N__29108\
        );

    \I__3801\ : Span4Mux_v
    port map (
            O => \N__29121\,
            I => \N__29103\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__29118\,
            I => \N__29103\
        );

    \I__3799\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29100\
        );

    \I__3798\ : Odrv12
    port map (
            O => \N__29114\,
            I => n9539
        );

    \I__3797\ : Odrv12
    port map (
            O => \N__29111\,
            I => n9539
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__29108\,
            I => n9539
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__29103\,
            I => n9539
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__29100\,
            I => n9539
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__29089\,
            I => \N__29085\
        );

    \I__3792\ : InMux
    port map (
            O => \N__29088\,
            I => \N__29082\
        );

    \I__3791\ : InMux
    port map (
            O => \N__29085\,
            I => \N__29079\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__29082\,
            I => data_out_frame_10_0
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__29079\,
            I => data_out_frame_10_0
        );

    \I__3788\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29071\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__29071\,
            I => \N__29065\
        );

    \I__3786\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29062\
        );

    \I__3785\ : InMux
    port map (
            O => \N__29069\,
            I => \N__29057\
        );

    \I__3784\ : InMux
    port map (
            O => \N__29068\,
            I => \N__29057\
        );

    \I__3783\ : Odrv4
    port map (
            O => \N__29065\,
            I => data_in_3_3
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__29062\,
            I => data_in_3_3
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__29057\,
            I => data_in_3_3
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__29050\,
            I => \N__29046\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__29049\,
            I => \N__29043\
        );

    \I__3778\ : InMux
    port map (
            O => \N__29046\,
            I => \N__29039\
        );

    \I__3777\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29036\
        );

    \I__3776\ : InMux
    port map (
            O => \N__29042\,
            I => \N__29033\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__29039\,
            I => \N__29029\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__29036\,
            I => \N__29024\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__29033\,
            I => \N__29024\
        );

    \I__3772\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29021\
        );

    \I__3771\ : Span4Mux_h
    port map (
            O => \N__29029\,
            I => \N__29016\
        );

    \I__3770\ : Span4Mux_h
    port map (
            O => \N__29024\,
            I => \N__29016\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__29021\,
            I => encoder1_position_18
        );

    \I__3768\ : Odrv4
    port map (
            O => \N__29016\,
            I => encoder1_position_18
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__29011\,
            I => \N__29007\
        );

    \I__3766\ : InMux
    port map (
            O => \N__29010\,
            I => \N__29004\
        );

    \I__3765\ : InMux
    port map (
            O => \N__29007\,
            I => \N__29001\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__29004\,
            I => data_out_frame_11_2
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__29001\,
            I => data_out_frame_11_2
        );

    \I__3762\ : InMux
    port map (
            O => \N__28996\,
            I => \N__28993\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__28993\,
            I => \N__28990\
        );

    \I__3760\ : Span4Mux_v
    port map (
            O => \N__28990\,
            I => \N__28987\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__28987\,
            I => \c0.n24177\
        );

    \I__3758\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28980\
        );

    \I__3757\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28977\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__28980\,
            I => \N__28974\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__28977\,
            I => \N__28969\
        );

    \I__3754\ : Span4Mux_h
    port map (
            O => \N__28974\,
            I => \N__28969\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__28969\,
            I => data_out_frame_5_0
        );

    \I__3752\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28962\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__28965\,
            I => \N__28959\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__28962\,
            I => \N__28955\
        );

    \I__3749\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28951\
        );

    \I__3748\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28948\
        );

    \I__3747\ : Span4Mux_v
    port map (
            O => \N__28955\,
            I => \N__28945\
        );

    \I__3746\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28942\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28939\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__28948\,
            I => encoder1_position_29
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__28945\,
            I => encoder1_position_29
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__28942\,
            I => encoder1_position_29
        );

    \I__3741\ : Odrv12
    port map (
            O => \N__28939\,
            I => encoder1_position_29
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__28930\,
            I => \N__28926\
        );

    \I__3739\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28923\
        );

    \I__3738\ : InMux
    port map (
            O => \N__28926\,
            I => \N__28920\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__28923\,
            I => \N__28917\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__28920\,
            I => data_out_frame_10_5
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__28917\,
            I => data_out_frame_10_5
        );

    \I__3734\ : InMux
    port map (
            O => \N__28912\,
            I => \N__28908\
        );

    \I__3733\ : InMux
    port map (
            O => \N__28911\,
            I => \N__28905\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__28908\,
            I => data_out_frame_12_3
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__28905\,
            I => data_out_frame_12_3
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__28900\,
            I => \c0.n7_adj_4492_cascade_\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__28897\,
            I => \N__28893\
        );

    \I__3728\ : InMux
    port map (
            O => \N__28896\,
            I => \N__28890\
        );

    \I__3727\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28885\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__28890\,
            I => \N__28882\
        );

    \I__3725\ : InMux
    port map (
            O => \N__28889\,
            I => \N__28877\
        );

    \I__3724\ : InMux
    port map (
            O => \N__28888\,
            I => \N__28877\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__28885\,
            I => data_in_1_5
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__28882\,
            I => data_in_1_5
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__28877\,
            I => data_in_1_5
        );

    \I__3720\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28867\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__28867\,
            I => \c0.n9_adj_4493\
        );

    \I__3718\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28861\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__28861\,
            I => \c0.n23600\
        );

    \I__3716\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28849\
        );

    \I__3715\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28849\
        );

    \I__3714\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28849\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__28849\,
            I => data_in_0_6
        );

    \I__3712\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28840\
        );

    \I__3711\ : InMux
    port map (
            O => \N__28845\,
            I => \N__28837\
        );

    \I__3710\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28832\
        );

    \I__3709\ : InMux
    port map (
            O => \N__28843\,
            I => \N__28832\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__28840\,
            I => \N__28825\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__28837\,
            I => \N__28825\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__28832\,
            I => \N__28825\
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__28825\,
            I => data_in_2_2
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__28822\,
            I => \N__28819\
        );

    \I__3703\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28815\
        );

    \I__3702\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28812\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__28815\,
            I => \N__28806\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__28812\,
            I => \N__28806\
        );

    \I__3699\ : InMux
    port map (
            O => \N__28811\,
            I => \N__28803\
        );

    \I__3698\ : Span4Mux_v
    port map (
            O => \N__28806\,
            I => \N__28800\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__28803\,
            I => data_in_0_3
        );

    \I__3696\ : Odrv4
    port map (
            O => \N__28800\,
            I => data_in_0_3
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__28795\,
            I => \c0.n14_adj_4495_cascade_\
        );

    \I__3694\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28789\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__28789\,
            I => \c0.n15_adj_4496\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__28786\,
            I => \N__28783\
        );

    \I__3691\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28778\
        );

    \I__3690\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28775\
        );

    \I__3689\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28772\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__28778\,
            I => \N__28767\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__28775\,
            I => \N__28762\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__28772\,
            I => \N__28762\
        );

    \I__3685\ : InMux
    port map (
            O => \N__28771\,
            I => \N__28759\
        );

    \I__3684\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28756\
        );

    \I__3683\ : Span4Mux_h
    port map (
            O => \N__28767\,
            I => \N__28753\
        );

    \I__3682\ : Span4Mux_v
    port map (
            O => \N__28762\,
            I => \N__28750\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__28759\,
            I => encoder1_position_31
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__28756\,
            I => encoder1_position_31
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__28753\,
            I => encoder1_position_31
        );

    \I__3678\ : Odrv4
    port map (
            O => \N__28750\,
            I => encoder1_position_31
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__28741\,
            I => \N__28737\
        );

    \I__3676\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28734\
        );

    \I__3675\ : InMux
    port map (
            O => \N__28737\,
            I => \N__28731\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__28734\,
            I => \N__28728\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__28731\,
            I => data_out_frame_10_7
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__28728\,
            I => data_out_frame_10_7
        );

    \I__3671\ : InMux
    port map (
            O => \N__28723\,
            I => \N__28719\
        );

    \I__3670\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28716\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__28719\,
            I => \N__28713\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__28716\,
            I => data_out_frame_8_7
        );

    \I__3667\ : Odrv4
    port map (
            O => \N__28713\,
            I => data_out_frame_8_7
        );

    \I__3666\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28705\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28701\
        );

    \I__3664\ : InMux
    port map (
            O => \N__28704\,
            I => \N__28698\
        );

    \I__3663\ : Span4Mux_v
    port map (
            O => \N__28701\,
            I => \N__28695\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__28698\,
            I => data_out_frame_11_7
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__28695\,
            I => data_out_frame_11_7
        );

    \I__3660\ : InMux
    port map (
            O => \N__28690\,
            I => \N__28687\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__28687\,
            I => \N__28684\
        );

    \I__3658\ : Span4Mux_v
    port map (
            O => \N__28684\,
            I => \N__28681\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__28681\,
            I => n2181
        );

    \I__3656\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28675\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__28675\,
            I => \N__28672\
        );

    \I__3654\ : Span4Mux_h
    port map (
            O => \N__28672\,
            I => \N__28669\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__28669\,
            I => \c0.n22224\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__28666\,
            I => \c0.n22224_cascade_\
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__28663\,
            I => \c0.n13349_cascade_\
        );

    \I__3650\ : InMux
    port map (
            O => \N__28660\,
            I => \N__28657\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__28657\,
            I => \N__28654\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__28654\,
            I => \c0.n6_adj_4334\
        );

    \I__3647\ : InMux
    port map (
            O => \N__28651\,
            I => \N__28648\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__28648\,
            I => \N__28645\
        );

    \I__3645\ : Span4Mux_h
    port map (
            O => \N__28645\,
            I => \N__28642\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__28642\,
            I => n24104
        );

    \I__3643\ : InMux
    port map (
            O => \N__28639\,
            I => \N__28636\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__28636\,
            I => \c0.n22405\
        );

    \I__3641\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28630\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__28630\,
            I => \c0.n22102\
        );

    \I__3639\ : CascadeMux
    port map (
            O => \N__28627\,
            I => \c0.n22361_cascade_\
        );

    \I__3638\ : InMux
    port map (
            O => \N__28624\,
            I => \N__28621\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__28621\,
            I => \N__28618\
        );

    \I__3636\ : Odrv4
    port map (
            O => \N__28618\,
            I => \c0.n10_adj_4314\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__28615\,
            I => \N__28612\
        );

    \I__3634\ : InMux
    port map (
            O => \N__28612\,
            I => \N__28607\
        );

    \I__3633\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28603\
        );

    \I__3632\ : InMux
    port map (
            O => \N__28610\,
            I => \N__28600\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__28607\,
            I => \N__28597\
        );

    \I__3630\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28594\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__28603\,
            I => \N__28591\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__28600\,
            I => encoder1_position_21
        );

    \I__3627\ : Odrv12
    port map (
            O => \N__28597\,
            I => encoder1_position_21
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__28594\,
            I => encoder1_position_21
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__28591\,
            I => encoder1_position_21
        );

    \I__3624\ : InMux
    port map (
            O => \N__28582\,
            I => \N__28579\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__28579\,
            I => \N__28576\
        );

    \I__3622\ : Span4Mux_v
    port map (
            O => \N__28576\,
            I => \N__28573\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__28573\,
            I => \N__28570\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__28570\,
            I => \c0.n24153\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__28567\,
            I => \N__28563\
        );

    \I__3618\ : InMux
    port map (
            O => \N__28566\,
            I => \N__28558\
        );

    \I__3617\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28558\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__28558\,
            I => data_out_frame_8_6
        );

    \I__3615\ : InMux
    port map (
            O => \N__28555\,
            I => \N__28552\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__28552\,
            I => \N__28549\
        );

    \I__3613\ : Span4Mux_h
    port map (
            O => \N__28549\,
            I => \N__28546\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__28546\,
            I => \c0.n24156\
        );

    \I__3611\ : InMux
    port map (
            O => \N__28543\,
            I => \N__28540\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__28540\,
            I => \N__28536\
        );

    \I__3609\ : InMux
    port map (
            O => \N__28539\,
            I => \N__28533\
        );

    \I__3608\ : Span4Mux_h
    port map (
            O => \N__28536\,
            I => \N__28530\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__28533\,
            I => data_out_frame_12_6
        );

    \I__3606\ : Odrv4
    port map (
            O => \N__28530\,
            I => data_out_frame_12_6
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__28525\,
            I => \N__28522\
        );

    \I__3604\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28518\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__28521\,
            I => \N__28515\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__28518\,
            I => \N__28512\
        );

    \I__3601\ : InMux
    port map (
            O => \N__28515\,
            I => \N__28509\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__28512\,
            I => \N__28506\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__28509\,
            I => data_out_frame_11_3
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__28506\,
            I => data_out_frame_11_3
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__28501\,
            I => \c0.n21110_cascade_\
        );

    \I__3596\ : InMux
    port map (
            O => \N__28498\,
            I => \N__28495\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__28495\,
            I => \N__28492\
        );

    \I__3594\ : Odrv12
    port map (
            O => \N__28492\,
            I => \c0.n14_adj_4514\
        );

    \I__3593\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28482\
        );

    \I__3592\ : InMux
    port map (
            O => \N__28488\,
            I => \N__28482\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__28487\,
            I => \N__28478\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__28482\,
            I => \N__28475\
        );

    \I__3589\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28471\
        );

    \I__3588\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28467\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__28475\,
            I => \N__28464\
        );

    \I__3586\ : InMux
    port map (
            O => \N__28474\,
            I => \N__28461\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__28471\,
            I => \N__28458\
        );

    \I__3584\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28455\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__28467\,
            I => \N__28452\
        );

    \I__3582\ : Span4Mux_h
    port map (
            O => \N__28464\,
            I => \N__28447\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__28461\,
            I => \N__28447\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__28458\,
            I => encoder1_position_22
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__28455\,
            I => encoder1_position_22
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__28452\,
            I => encoder1_position_22
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__28447\,
            I => encoder1_position_22
        );

    \I__3576\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28435\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__28435\,
            I => \N__28432\
        );

    \I__3574\ : Span4Mux_h
    port map (
            O => \N__28432\,
            I => \N__28429\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__28429\,
            I => n2201
        );

    \I__3572\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28423\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__28423\,
            I => \N__28419\
        );

    \I__3570\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28416\
        );

    \I__3569\ : Span4Mux_h
    port map (
            O => \N__28419\,
            I => \N__28413\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__28416\,
            I => \N__28410\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__28413\,
            I => \c0.n22277\
        );

    \I__3566\ : Odrv12
    port map (
            O => \N__28410\,
            I => \c0.n22277\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__28405\,
            I => \c0.n22102_cascade_\
        );

    \I__3564\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28399\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__28399\,
            I => \c0.n22293\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__28396\,
            I => \c0.n15_adj_4325_cascade_\
        );

    \I__3561\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28384\
        );

    \I__3560\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28384\
        );

    \I__3559\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28384\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__28384\,
            I => \N__28381\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__28381\,
            I => \c0.n21041\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__28378\,
            I => \c0.n21041_cascade_\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__28375\,
            I => \c0.n6_adj_4313_cascade_\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__28372\,
            I => \c0.n21156_cascade_\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__28369\,
            I => \c0.n21175_cascade_\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__28366\,
            I => \c0.n20276_cascade_\
        );

    \I__3551\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28360\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__28360\,
            I => \c0.n22066\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__28357\,
            I => \N__28353\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__28356\,
            I => \N__28349\
        );

    \I__3547\ : InMux
    port map (
            O => \N__28353\,
            I => \N__28346\
        );

    \I__3546\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28339\
        );

    \I__3545\ : InMux
    port map (
            O => \N__28349\,
            I => \N__28339\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__28346\,
            I => \N__28335\
        );

    \I__3543\ : InMux
    port map (
            O => \N__28345\,
            I => \N__28329\
        );

    \I__3542\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28329\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__28339\,
            I => \N__28326\
        );

    \I__3540\ : InMux
    port map (
            O => \N__28338\,
            I => \N__28322\
        );

    \I__3539\ : Span4Mux_h
    port map (
            O => \N__28335\,
            I => \N__28318\
        );

    \I__3538\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28315\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__28329\,
            I => \N__28312\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__28326\,
            I => \N__28308\
        );

    \I__3535\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28305\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__28322\,
            I => \N__28302\
        );

    \I__3533\ : InMux
    port map (
            O => \N__28321\,
            I => \N__28299\
        );

    \I__3532\ : Span4Mux_v
    port map (
            O => \N__28318\,
            I => \N__28292\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__28315\,
            I => \N__28292\
        );

    \I__3530\ : Span4Mux_h
    port map (
            O => \N__28312\,
            I => \N__28292\
        );

    \I__3529\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28289\
        );

    \I__3528\ : Span4Mux_h
    port map (
            O => \N__28308\,
            I => \N__28286\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__28305\,
            I => encoder1_position_3
        );

    \I__3526\ : Odrv4
    port map (
            O => \N__28302\,
            I => encoder1_position_3
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__28299\,
            I => encoder1_position_3
        );

    \I__3524\ : Odrv4
    port map (
            O => \N__28292\,
            I => encoder1_position_3
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__28289\,
            I => encoder1_position_3
        );

    \I__3522\ : Odrv4
    port map (
            O => \N__28286\,
            I => encoder1_position_3
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__28273\,
            I => \c0.n21071_cascade_\
        );

    \I__3520\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28266\
        );

    \I__3519\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28263\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__28266\,
            I => \N__28258\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__28263\,
            I => \N__28258\
        );

    \I__3516\ : Odrv4
    port map (
            O => \N__28258\,
            I => \data_out_frame_29__2__N_1749\
        );

    \I__3515\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28252\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__28252\,
            I => \c0.n17_adj_4501\
        );

    \I__3513\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28246\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__28246\,
            I => \c0.data_out_frame_29_0\
        );

    \I__3511\ : InMux
    port map (
            O => \N__28243\,
            I => \N__28240\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28237\
        );

    \I__3509\ : Span4Mux_v
    port map (
            O => \N__28237\,
            I => \N__28234\
        );

    \I__3508\ : Span4Mux_v
    port map (
            O => \N__28234\,
            I => \N__28231\
        );

    \I__3507\ : Span4Mux_v
    port map (
            O => \N__28231\,
            I => \N__28228\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__28228\,
            I => \c0.n26_adj_4423\
        );

    \I__3505\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28222\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__28222\,
            I => \c0.n16_adj_4500\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__28219\,
            I => \N__28215\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__28218\,
            I => \N__28212\
        );

    \I__3501\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28209\
        );

    \I__3500\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28206\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__28209\,
            I => \N__28203\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__28206\,
            I => \N__28200\
        );

    \I__3497\ : Span4Mux_h
    port map (
            O => \N__28203\,
            I => \N__28195\
        );

    \I__3496\ : Span4Mux_h
    port map (
            O => \N__28200\,
            I => \N__28195\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__28195\,
            I => \c0.n10422\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__28192\,
            I => \c0.n14_adj_4340_cascade_\
        );

    \I__3493\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28186\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__28186\,
            I => \c0.n20320\
        );

    \I__3491\ : CascadeMux
    port map (
            O => \N__28183\,
            I => \c0.n20320_cascade_\
        );

    \I__3490\ : CascadeMux
    port map (
            O => \N__28180\,
            I => \c0.n22180_cascade_\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__28177\,
            I => \c0.n10498_cascade_\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__28174\,
            I => \c0.n20253_cascade_\
        );

    \I__3487\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28166\
        );

    \I__3486\ : InMux
    port map (
            O => \N__28170\,
            I => \N__28161\
        );

    \I__3485\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28161\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__28166\,
            I => \N__28156\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__28161\,
            I => \N__28156\
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__28156\,
            I => \c0.n21229\
        );

    \I__3481\ : InMux
    port map (
            O => \N__28153\,
            I => \N__28150\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__28150\,
            I => \c0.n15_adj_4513\
        );

    \I__3479\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28144\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__28144\,
            I => \quad_counter0.n28_adj_4202\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__28141\,
            I => \quad_counter0.n27_adj_4204_cascade_\
        );

    \I__3476\ : InMux
    port map (
            O => \N__28138\,
            I => \N__28135\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__28135\,
            I => \quad_counter0.n25_adj_4205\
        );

    \I__3474\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28126\
        );

    \I__3473\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28126\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__28126\,
            I => n9821
        );

    \I__3471\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28119\
        );

    \I__3470\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28116\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__28119\,
            I => \quad_counter0.a_delay_counter_12\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__28116\,
            I => \quad_counter0.a_delay_counter_12\
        );

    \I__3467\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28107\
        );

    \I__3466\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28104\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__28107\,
            I => \quad_counter0.a_delay_counter_13\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__28104\,
            I => \quad_counter0.a_delay_counter_13\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__28099\,
            I => \N__28095\
        );

    \I__3462\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28092\
        );

    \I__3461\ : InMux
    port map (
            O => \N__28095\,
            I => \N__28089\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__28092\,
            I => \quad_counter0.a_delay_counter_6\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__28089\,
            I => \quad_counter0.a_delay_counter_6\
        );

    \I__3458\ : InMux
    port map (
            O => \N__28084\,
            I => \N__28080\
        );

    \I__3457\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28077\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__28080\,
            I => \quad_counter0.a_delay_counter_9\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__28077\,
            I => \quad_counter0.a_delay_counter_9\
        );

    \I__3454\ : InMux
    port map (
            O => \N__28072\,
            I => \N__28069\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__28069\,
            I => \quad_counter0.n26_adj_4203\
        );

    \I__3452\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28062\
        );

    \I__3451\ : InMux
    port map (
            O => \N__28065\,
            I => \N__28059\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__28062\,
            I => \N__28056\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__28059\,
            I => \N__28053\
        );

    \I__3448\ : Span4Mux_v
    port map (
            O => \N__28056\,
            I => \N__28050\
        );

    \I__3447\ : Span4Mux_v
    port map (
            O => \N__28053\,
            I => \N__28047\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__28050\,
            I => \data_out_frame_28__3__N_1881\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__28047\,
            I => \data_out_frame_28__3__N_1881\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__28042\,
            I => \N__28039\
        );

    \I__3443\ : InMux
    port map (
            O => \N__28039\,
            I => \N__28036\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__28036\,
            I => \N__28032\
        );

    \I__3441\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28029\
        );

    \I__3440\ : Span4Mux_h
    port map (
            O => \N__28032\,
            I => \N__28026\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__28029\,
            I => \N__28023\
        );

    \I__3438\ : Span4Mux_v
    port map (
            O => \N__28026\,
            I => \N__28020\
        );

    \I__3437\ : Span4Mux_h
    port map (
            O => \N__28023\,
            I => \N__28017\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__28020\,
            I => \c0.n20257\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__28017\,
            I => \c0.n20257\
        );

    \I__3434\ : InMux
    port map (
            O => \N__28012\,
            I => \N__28009\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__28009\,
            I => \c0.n21062\
        );

    \I__3432\ : InMux
    port map (
            O => \N__28006\,
            I => \N__28003\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__28003\,
            I => \N__28000\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__28000\,
            I => \c0.data_out_frame_28_1\
        );

    \I__3429\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27994\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__27994\,
            I => \c0.data_out_frame_29_1\
        );

    \I__3427\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27988\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__27988\,
            I => \N__27985\
        );

    \I__3425\ : Span4Mux_v
    port map (
            O => \N__27985\,
            I => \N__27982\
        );

    \I__3424\ : Span4Mux_v
    port map (
            O => \N__27982\,
            I => \N__27979\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__27979\,
            I => \c0.n26_adj_4519\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__27976\,
            I => \c0.n12542_cascade_\
        );

    \I__3421\ : InMux
    port map (
            O => \N__27973\,
            I => \N__27966\
        );

    \I__3420\ : InMux
    port map (
            O => \N__27972\,
            I => \N__27966\
        );

    \I__3419\ : InMux
    port map (
            O => \N__27971\,
            I => \N__27963\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__27966\,
            I => \quad_counter0.B_delayed\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__27963\,
            I => \quad_counter0.B_delayed\
        );

    \I__3416\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27954\
        );

    \I__3415\ : InMux
    port map (
            O => \N__27957\,
            I => \N__27951\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__27954\,
            I => \quad_counter0.a_delay_counter_3\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__27951\,
            I => \quad_counter0.a_delay_counter_3\
        );

    \I__3412\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27942\
        );

    \I__3411\ : InMux
    port map (
            O => \N__27945\,
            I => \N__27939\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__27942\,
            I => \quad_counter0.a_delay_counter_8\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__27939\,
            I => \quad_counter0.a_delay_counter_8\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__27934\,
            I => \N__27930\
        );

    \I__3407\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27927\
        );

    \I__3406\ : InMux
    port map (
            O => \N__27930\,
            I => \N__27924\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__27927\,
            I => \quad_counter0.a_delay_counter_2\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__27924\,
            I => \quad_counter0.a_delay_counter_2\
        );

    \I__3403\ : InMux
    port map (
            O => \N__27919\,
            I => \N__27915\
        );

    \I__3402\ : InMux
    port map (
            O => \N__27918\,
            I => \N__27912\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__27915\,
            I => \quad_counter0.a_delay_counter_1\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__27912\,
            I => \quad_counter0.a_delay_counter_1\
        );

    \I__3399\ : InMux
    port map (
            O => \N__27907\,
            I => \N__27903\
        );

    \I__3398\ : InMux
    port map (
            O => \N__27906\,
            I => \N__27900\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__27903\,
            I => \quad_counter0.a_delay_counter_5\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__27900\,
            I => \quad_counter0.a_delay_counter_5\
        );

    \I__3395\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27891\
        );

    \I__3394\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27888\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__27891\,
            I => \quad_counter0.a_delay_counter_11\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__27888\,
            I => \quad_counter0.a_delay_counter_11\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__27883\,
            I => \N__27879\
        );

    \I__3390\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27876\
        );

    \I__3389\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27873\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__27876\,
            I => \quad_counter0.a_delay_counter_4\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__27873\,
            I => \quad_counter0.a_delay_counter_4\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__27868\,
            I => \N__27865\
        );

    \I__3385\ : InMux
    port map (
            O => \N__27865\,
            I => \N__27860\
        );

    \I__3384\ : InMux
    port map (
            O => \N__27864\,
            I => \N__27855\
        );

    \I__3383\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27852\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__27860\,
            I => \N__27849\
        );

    \I__3381\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27844\
        );

    \I__3380\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27844\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__27855\,
            I => \N__27841\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__27852\,
            I => \A_filtered\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__27849\,
            I => \A_filtered\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__27844\,
            I => \A_filtered\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__27841\,
            I => \A_filtered\
        );

    \I__3374\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27826\
        );

    \I__3373\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27826\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__27826\,
            I => \N__27821\
        );

    \I__3371\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27818\
        );

    \I__3370\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27815\
        );

    \I__3369\ : Span4Mux_h
    port map (
            O => \N__27821\,
            I => \N__27808\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__27818\,
            I => \N__27808\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__27815\,
            I => \N__27808\
        );

    \I__3366\ : Span4Mux_v
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__3365\ : Sp12to4
    port map (
            O => \N__27805\,
            I => \N__27802\
        );

    \I__3364\ : Odrv12
    port map (
            O => \N__27802\,
            I => \PIN_7_c\
        );

    \I__3363\ : CascadeMux
    port map (
            O => \N__27799\,
            I => \N__27796\
        );

    \I__3362\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27790\
        );

    \I__3361\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27790\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__27790\,
            I => \N__27786\
        );

    \I__3359\ : InMux
    port map (
            O => \N__27789\,
            I => \N__27783\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__27786\,
            I => \N__27780\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__27783\,
            I => \N__27777\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__27780\,
            I => \quadA_delayed\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__27777\,
            I => \quadA_delayed\
        );

    \I__3354\ : CEMux
    port map (
            O => \N__27772\,
            I => \N__27769\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__27769\,
            I => \N__27765\
        );

    \I__3352\ : CEMux
    port map (
            O => \N__27768\,
            I => \N__27762\
        );

    \I__3351\ : Span4Mux_h
    port map (
            O => \N__27765\,
            I => \N__27759\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__27762\,
            I => \N__27756\
        );

    \I__3349\ : Span4Mux_h
    port map (
            O => \N__27759\,
            I => \N__27753\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__27756\,
            I => n14421
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__27753\,
            I => n14421
        );

    \I__3346\ : SRMux
    port map (
            O => \N__27748\,
            I => \N__27743\
        );

    \I__3345\ : SRMux
    port map (
            O => \N__27747\,
            I => \N__27740\
        );

    \I__3344\ : InMux
    port map (
            O => \N__27746\,
            I => \N__27737\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__27743\,
            I => \N__27734\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__27740\,
            I => \N__27729\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__27737\,
            I => \N__27729\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__27734\,
            I => \a_delay_counter_15__N_4124\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__27729\,
            I => \a_delay_counter_15__N_4124\
        );

    \I__3338\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27721\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__27721\,
            I => n39
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__27718\,
            I => \n14421_cascade_\
        );

    \I__3335\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27710\
        );

    \I__3334\ : InMux
    port map (
            O => \N__27714\,
            I => \N__27707\
        );

    \I__3333\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27704\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__27710\,
            I => a_delay_counter_0
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__27707\,
            I => a_delay_counter_0
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__27704\,
            I => a_delay_counter_0
        );

    \I__3329\ : InMux
    port map (
            O => \N__27697\,
            I => \N__27693\
        );

    \I__3328\ : InMux
    port map (
            O => \N__27696\,
            I => \N__27690\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__27693\,
            I => \quad_counter0.a_delay_counter_14\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__27690\,
            I => \quad_counter0.a_delay_counter_14\
        );

    \I__3325\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27681\
        );

    \I__3324\ : InMux
    port map (
            O => \N__27684\,
            I => \N__27678\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__27681\,
            I => \quad_counter0.a_delay_counter_15\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__27678\,
            I => \quad_counter0.a_delay_counter_15\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__27673\,
            I => \N__27669\
        );

    \I__3320\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27666\
        );

    \I__3319\ : InMux
    port map (
            O => \N__27669\,
            I => \N__27663\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__27666\,
            I => \quad_counter0.a_delay_counter_7\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__27663\,
            I => \quad_counter0.a_delay_counter_7\
        );

    \I__3316\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27654\
        );

    \I__3315\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27651\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__27654\,
            I => \quad_counter0.a_delay_counter_10\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__27651\,
            I => \quad_counter0.a_delay_counter_10\
        );

    \I__3312\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27642\
        );

    \I__3311\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27639\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__27642\,
            I => \quad_counter0.b_delay_counter_3\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__27639\,
            I => \quad_counter0.b_delay_counter_3\
        );

    \I__3308\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27630\
        );

    \I__3307\ : InMux
    port map (
            O => \N__27633\,
            I => \N__27627\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__27630\,
            I => \quad_counter0.b_delay_counter_9\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__27627\,
            I => \quad_counter0.b_delay_counter_9\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__27622\,
            I => \N__27618\
        );

    \I__3303\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27615\
        );

    \I__3302\ : InMux
    port map (
            O => \N__27618\,
            I => \N__27612\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__27615\,
            I => \quad_counter0.b_delay_counter_4\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__27612\,
            I => \quad_counter0.b_delay_counter_4\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__27607\,
            I => \N__27603\
        );

    \I__3298\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27599\
        );

    \I__3297\ : InMux
    port map (
            O => \N__27603\,
            I => \N__27596\
        );

    \I__3296\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27593\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__27599\,
            I => \N__27590\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__27596\,
            I => b_delay_counter_0
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__27593\,
            I => b_delay_counter_0
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__27590\,
            I => b_delay_counter_0
        );

    \I__3291\ : InMux
    port map (
            O => \N__27583\,
            I => \N__27580\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__27580\,
            I => \N__27575\
        );

    \I__3289\ : InMux
    port map (
            O => \N__27579\,
            I => \N__27569\
        );

    \I__3288\ : InMux
    port map (
            O => \N__27578\,
            I => \N__27569\
        );

    \I__3287\ : Span4Mux_v
    port map (
            O => \N__27575\,
            I => \N__27566\
        );

    \I__3286\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27563\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__27569\,
            I => \N__27560\
        );

    \I__3284\ : Span4Mux_h
    port map (
            O => \N__27566\,
            I => \N__27555\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__27563\,
            I => \N__27555\
        );

    \I__3282\ : Sp12to4
    port map (
            O => \N__27560\,
            I => \N__27552\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__27555\,
            I => \N__27549\
        );

    \I__3280\ : Span12Mux_v
    port map (
            O => \N__27552\,
            I => \N__27546\
        );

    \I__3279\ : Span4Mux_v
    port map (
            O => \N__27549\,
            I => \N__27543\
        );

    \I__3278\ : Odrv12
    port map (
            O => \N__27546\,
            I => \PIN_8_c\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__27543\,
            I => \PIN_8_c\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__27538\,
            I => \N__27535\
        );

    \I__3275\ : InMux
    port map (
            O => \N__27535\,
            I => \N__27532\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__27532\,
            I => \N__27527\
        );

    \I__3273\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27522\
        );

    \I__3272\ : InMux
    port map (
            O => \N__27530\,
            I => \N__27522\
        );

    \I__3271\ : Span4Mux_v
    port map (
            O => \N__27527\,
            I => \N__27519\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__27522\,
            I => \N__27516\
        );

    \I__3269\ : Span4Mux_h
    port map (
            O => \N__27519\,
            I => \N__27513\
        );

    \I__3268\ : Span4Mux_v
    port map (
            O => \N__27516\,
            I => \N__27510\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__27513\,
            I => \quadB_delayed\
        );

    \I__3266\ : Odrv4
    port map (
            O => \N__27510\,
            I => \quadB_delayed\
        );

    \I__3265\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27496\
        );

    \I__3264\ : InMux
    port map (
            O => \N__27504\,
            I => \N__27496\
        );

    \I__3263\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27496\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__27496\,
            I => \B_filtered\
        );

    \I__3261\ : InMux
    port map (
            O => \N__27493\,
            I => \N__27489\
        );

    \I__3260\ : InMux
    port map (
            O => \N__27492\,
            I => \N__27486\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__27489\,
            I => \quad_counter0.b_delay_counter_13\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__27486\,
            I => \quad_counter0.b_delay_counter_13\
        );

    \I__3257\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27477\
        );

    \I__3256\ : InMux
    port map (
            O => \N__27480\,
            I => \N__27474\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__27477\,
            I => \quad_counter0.b_delay_counter_1\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__27474\,
            I => \quad_counter0.b_delay_counter_1\
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__27469\,
            I => \N__27465\
        );

    \I__3252\ : InMux
    port map (
            O => \N__27468\,
            I => \N__27462\
        );

    \I__3251\ : InMux
    port map (
            O => \N__27465\,
            I => \N__27459\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__27462\,
            I => \quad_counter0.b_delay_counter_2\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__27459\,
            I => \quad_counter0.b_delay_counter_2\
        );

    \I__3248\ : InMux
    port map (
            O => \N__27454\,
            I => \N__27450\
        );

    \I__3247\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27447\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__27450\,
            I => \quad_counter0.b_delay_counter_5\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__27447\,
            I => \quad_counter0.b_delay_counter_5\
        );

    \I__3244\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27438\
        );

    \I__3243\ : InMux
    port map (
            O => \N__27441\,
            I => \N__27435\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__27438\,
            I => \quad_counter0.b_delay_counter_11\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__27435\,
            I => \quad_counter0.b_delay_counter_11\
        );

    \I__3240\ : InMux
    port map (
            O => \N__27430\,
            I => \N__27426\
        );

    \I__3239\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27423\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__27426\,
            I => \quad_counter0.b_delay_counter_10\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__27423\,
            I => \quad_counter0.b_delay_counter_10\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__27418\,
            I => \N__27414\
        );

    \I__3235\ : InMux
    port map (
            O => \N__27417\,
            I => \N__27411\
        );

    \I__3234\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27408\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__27411\,
            I => \quad_counter0.b_delay_counter_8\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__27408\,
            I => \quad_counter0.b_delay_counter_8\
        );

    \I__3231\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27399\
        );

    \I__3230\ : InMux
    port map (
            O => \N__27402\,
            I => \N__27396\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__27399\,
            I => \quad_counter0.b_delay_counter_6\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__27396\,
            I => \quad_counter0.b_delay_counter_6\
        );

    \I__3227\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27388\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__27388\,
            I => \quad_counter0.n28_adj_4198\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__27385\,
            I => \quad_counter0.n26_adj_4199_cascade_\
        );

    \I__3224\ : InMux
    port map (
            O => \N__27382\,
            I => \N__27379\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__27379\,
            I => \quad_counter0.n25_adj_4201\
        );

    \I__3222\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27373\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__27373\,
            I => \N__27369\
        );

    \I__3220\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27366\
        );

    \I__3219\ : Span4Mux_h
    port map (
            O => \N__27369\,
            I => \N__27363\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__27366\,
            I => n12909
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__27363\,
            I => n12909
        );

    \I__3216\ : InMux
    port map (
            O => \N__27358\,
            I => \N__27355\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__27355\,
            I => \quad_counter0.A_delayed\
        );

    \I__3214\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27349\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__27349\,
            I => \N__27346\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__27346\,
            I => n10_adj_4535
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__27343\,
            I => \N__27339\
        );

    \I__3210\ : CascadeMux
    port map (
            O => \N__27342\,
            I => \N__27335\
        );

    \I__3209\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27331\
        );

    \I__3208\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27326\
        );

    \I__3207\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27323\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__27334\,
            I => \N__27319\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__27331\,
            I => \N__27316\
        );

    \I__3204\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27311\
        );

    \I__3203\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27311\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__27326\,
            I => \N__27305\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__27323\,
            I => \N__27302\
        );

    \I__3200\ : InMux
    port map (
            O => \N__27322\,
            I => \N__27297\
        );

    \I__3199\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27297\
        );

    \I__3198\ : Span4Mux_v
    port map (
            O => \N__27316\,
            I => \N__27292\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__27311\,
            I => \N__27292\
        );

    \I__3196\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27289\
        );

    \I__3195\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27286\
        );

    \I__3194\ : InMux
    port map (
            O => \N__27308\,
            I => \N__27283\
        );

    \I__3193\ : Span4Mux_h
    port map (
            O => \N__27305\,
            I => \N__27280\
        );

    \I__3192\ : Span4Mux_h
    port map (
            O => \N__27302\,
            I => \N__27277\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__27297\,
            I => \N__27272\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__27292\,
            I => \N__27272\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__27289\,
            I => \N__27269\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__27286\,
            I => byte_transmit_counter_5
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__27283\,
            I => byte_transmit_counter_5
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__27280\,
            I => byte_transmit_counter_5
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__27277\,
            I => byte_transmit_counter_5
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__27272\,
            I => byte_transmit_counter_5
        );

    \I__3183\ : Odrv12
    port map (
            O => \N__27269\,
            I => byte_transmit_counter_5
        );

    \I__3182\ : InMux
    port map (
            O => \N__27256\,
            I => \N__27250\
        );

    \I__3181\ : InMux
    port map (
            O => \N__27255\,
            I => \N__27250\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__27250\,
            I => \r_Tx_Data_1\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__27247\,
            I => \N__27242\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__27246\,
            I => \N__27239\
        );

    \I__3177\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27232\
        );

    \I__3176\ : InMux
    port map (
            O => \N__27242\,
            I => \N__27232\
        );

    \I__3175\ : InMux
    port map (
            O => \N__27239\,
            I => \N__27232\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__27232\,
            I => data_in_0_7
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__27229\,
            I => \N__27225\
        );

    \I__3172\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27222\
        );

    \I__3171\ : InMux
    port map (
            O => \N__27225\,
            I => \N__27219\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__27222\,
            I => \N__27214\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__27219\,
            I => \N__27214\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__27214\,
            I => data_out_frame_5_3
        );

    \I__3167\ : InMux
    port map (
            O => \N__27211\,
            I => \N__27207\
        );

    \I__3166\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27204\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__27207\,
            I => \N__27201\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__27204\,
            I => data_out_frame_6_3
        );

    \I__3163\ : Odrv12
    port map (
            O => \N__27201\,
            I => data_out_frame_6_3
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__27196\,
            I => \N__27193\
        );

    \I__3161\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27190\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__27190\,
            I => \N__27187\
        );

    \I__3159\ : Span4Mux_h
    port map (
            O => \N__27187\,
            I => \N__27184\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__27184\,
            I => \c0.n5\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__27181\,
            I => \N__27177\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__27180\,
            I => \N__27174\
        );

    \I__3155\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27171\
        );

    \I__3154\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27168\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27165\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__27168\,
            I => \N__27160\
        );

    \I__3151\ : Span4Mux_h
    port map (
            O => \N__27165\,
            I => \N__27160\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__27160\,
            I => data_out_frame_5_5
        );

    \I__3149\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27153\
        );

    \I__3148\ : InMux
    port map (
            O => \N__27156\,
            I => \N__27150\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__27153\,
            I => \N__27147\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__27150\,
            I => data_out_frame_11_0
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__27147\,
            I => data_out_frame_11_0
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__27142\,
            I => \c0.n24165_cascade_\
        );

    \I__3143\ : InMux
    port map (
            O => \N__27139\,
            I => \N__27136\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__27136\,
            I => \c0.n24168\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__27133\,
            I => \N__27130\
        );

    \I__3140\ : InMux
    port map (
            O => \N__27130\,
            I => \N__27127\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__27127\,
            I => \c0.n11_adj_4218\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__27124\,
            I => \N__27120\
        );

    \I__3137\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27115\
        );

    \I__3136\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27115\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__27115\,
            I => data_out_frame_11_5
        );

    \I__3134\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27109\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__27109\,
            I => \N__27105\
        );

    \I__3132\ : InMux
    port map (
            O => \N__27108\,
            I => \N__27102\
        );

    \I__3131\ : Span4Mux_v
    port map (
            O => \N__27105\,
            I => \N__27099\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__27102\,
            I => data_out_frame_9_5
        );

    \I__3129\ : Odrv4
    port map (
            O => \N__27099\,
            I => data_out_frame_9_5
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__27094\,
            I => \c0.n24141_cascade_\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__27091\,
            I => \N__27088\
        );

    \I__3126\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27082\
        );

    \I__3125\ : InMux
    port map (
            O => \N__27087\,
            I => \N__27082\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__27082\,
            I => data_out_frame_8_5
        );

    \I__3123\ : InMux
    port map (
            O => \N__27079\,
            I => \N__27076\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__27076\,
            I => \N__27073\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__27073\,
            I => \c0.n24144\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__27070\,
            I => \N__27067\
        );

    \I__3119\ : InMux
    port map (
            O => \N__27067\,
            I => \N__27063\
        );

    \I__3118\ : InMux
    port map (
            O => \N__27066\,
            I => \N__27060\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__27063\,
            I => \r_Tx_Data_7\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__27060\,
            I => \r_Tx_Data_7\
        );

    \I__3115\ : InMux
    port map (
            O => \N__27055\,
            I => \N__27051\
        );

    \I__3114\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27048\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__27051\,
            I => \r_Tx_Data_3\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__27048\,
            I => \r_Tx_Data_3\
        );

    \I__3111\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27037\
        );

    \I__3110\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27029\
        );

    \I__3109\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27029\
        );

    \I__3108\ : InMux
    port map (
            O => \N__27040\,
            I => \N__27029\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__27037\,
            I => \N__27026\
        );

    \I__3106\ : InMux
    port map (
            O => \N__27036\,
            I => \N__27023\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__27029\,
            I => \r_Bit_Index_2_adj_4551\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__27026\,
            I => \r_Bit_Index_2_adj_4551\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__27023\,
            I => \r_Bit_Index_2_adj_4551\
        );

    \I__3102\ : InMux
    port map (
            O => \N__27016\,
            I => \N__27013\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__27013\,
            I => \N__27010\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__27010\,
            I => \N__27006\
        );

    \I__3099\ : InMux
    port map (
            O => \N__27009\,
            I => \N__27003\
        );

    \I__3098\ : Span4Mux_h
    port map (
            O => \N__27006\,
            I => \N__27000\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__27003\,
            I => \N__26997\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__27000\,
            I => n4_adj_4554
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__26997\,
            I => n4_adj_4554
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__26992\,
            I => \n24189_cascade_\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__26989\,
            I => \N__26984\
        );

    \I__3092\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26979\
        );

    \I__3091\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26979\
        );

    \I__3090\ : InMux
    port map (
            O => \N__26984\,
            I => \N__26975\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__26979\,
            I => \N__26972\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__26978\,
            I => \N__26967\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__26975\,
            I => \N__26963\
        );

    \I__3086\ : Span4Mux_h
    port map (
            O => \N__26972\,
            I => \N__26960\
        );

    \I__3085\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26953\
        );

    \I__3084\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26953\
        );

    \I__3083\ : InMux
    port map (
            O => \N__26967\,
            I => \N__26953\
        );

    \I__3082\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26950\
        );

    \I__3081\ : Span4Mux_v
    port map (
            O => \N__26963\,
            I => \N__26947\
        );

    \I__3080\ : Odrv4
    port map (
            O => \N__26960\,
            I => \r_Bit_Index_1_adj_4552\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__26953\,
            I => \r_Bit_Index_1_adj_4552\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__26950\,
            I => \r_Bit_Index_1_adj_4552\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__26947\,
            I => \r_Bit_Index_1_adj_4552\
        );

    \I__3076\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26935\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__26935\,
            I => \c0.n6_adj_4392\
        );

    \I__3074\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26928\
        );

    \I__3073\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26925\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__26928\,
            I => \N__26922\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__26925\,
            I => \N__26917\
        );

    \I__3070\ : Span4Mux_h
    port map (
            O => \N__26922\,
            I => \N__26917\
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__26917\,
            I => \c0.byte_transmit_counter_6\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__26914\,
            I => \c0.n23574_cascade_\
        );

    \I__3067\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26907\
        );

    \I__3066\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26904\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__26907\,
            I => \N__26901\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__26904\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__3063\ : Odrv12
    port map (
            O => \N__26901\,
            I => \c0.byte_transmit_counter_7\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__26896\,
            I => \c0.n38_adj_4387_cascade_\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__26893\,
            I => \N__26890\
        );

    \I__3060\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26886\
        );

    \I__3059\ : InMux
    port map (
            O => \N__26889\,
            I => \N__26883\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__26886\,
            I => \N__26880\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__26883\,
            I => data_out_frame_5_2
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__26880\,
            I => data_out_frame_5_2
        );

    \I__3055\ : InMux
    port map (
            O => \N__26875\,
            I => \N__26870\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__26874\,
            I => \N__26867\
        );

    \I__3053\ : InMux
    port map (
            O => \N__26873\,
            I => \N__26860\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__26870\,
            I => \N__26857\
        );

    \I__3051\ : InMux
    port map (
            O => \N__26867\,
            I => \N__26854\
        );

    \I__3050\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26851\
        );

    \I__3049\ : InMux
    port map (
            O => \N__26865\,
            I => \N__26848\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__26864\,
            I => \N__26845\
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__26863\,
            I => \N__26842\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__26860\,
            I => \N__26839\
        );

    \I__3045\ : Span4Mux_v
    port map (
            O => \N__26857\,
            I => \N__26834\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__26854\,
            I => \N__26834\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__26851\,
            I => \N__26831\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__26848\,
            I => \N__26828\
        );

    \I__3041\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26825\
        );

    \I__3040\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26822\
        );

    \I__3039\ : Span4Mux_h
    port map (
            O => \N__26839\,
            I => \N__26819\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__26834\,
            I => \N__26814\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__26831\,
            I => \N__26814\
        );

    \I__3036\ : Span4Mux_h
    port map (
            O => \N__26828\,
            I => \N__26811\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__26825\,
            I => \N__26806\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__26822\,
            I => \N__26806\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__26819\,
            I => n23768
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__26814\,
            I => n23768
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__26811\,
            I => n23768
        );

    \I__3030\ : Odrv12
    port map (
            O => \N__26806\,
            I => n23768
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__26797\,
            I => \N__26793\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__26796\,
            I => \N__26785\
        );

    \I__3027\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26776\
        );

    \I__3026\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26771\
        );

    \I__3025\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26771\
        );

    \I__3024\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26766\
        );

    \I__3023\ : InMux
    port map (
            O => \N__26789\,
            I => \N__26766\
        );

    \I__3022\ : InMux
    port map (
            O => \N__26788\,
            I => \N__26761\
        );

    \I__3021\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26761\
        );

    \I__3020\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26756\
        );

    \I__3019\ : InMux
    port map (
            O => \N__26783\,
            I => \N__26756\
        );

    \I__3018\ : InMux
    port map (
            O => \N__26782\,
            I => \N__26749\
        );

    \I__3017\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26749\
        );

    \I__3016\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26749\
        );

    \I__3015\ : InMux
    port map (
            O => \N__26779\,
            I => \N__26746\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__26776\,
            I => \N__26739\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__26771\,
            I => \N__26736\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__26766\,
            I => \N__26733\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__26761\,
            I => \N__26730\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__26756\,
            I => \N__26723\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26723\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26723\
        );

    \I__3007\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26720\
        );

    \I__3006\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26715\
        );

    \I__3005\ : InMux
    port map (
            O => \N__26743\,
            I => \N__26715\
        );

    \I__3004\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26712\
        );

    \I__3003\ : Span4Mux_h
    port map (
            O => \N__26739\,
            I => \N__26709\
        );

    \I__3002\ : Span4Mux_h
    port map (
            O => \N__26736\,
            I => \N__26704\
        );

    \I__3001\ : Span4Mux_h
    port map (
            O => \N__26733\,
            I => \N__26704\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__26730\,
            I => \N__26701\
        );

    \I__2999\ : Span4Mux_v
    port map (
            O => \N__26723\,
            I => \N__26696\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__26720\,
            I => \N__26696\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__26715\,
            I => byte_transmit_counter_4
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__26712\,
            I => byte_transmit_counter_4
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__26709\,
            I => byte_transmit_counter_4
        );

    \I__2994\ : Odrv4
    port map (
            O => \N__26704\,
            I => byte_transmit_counter_4
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__26701\,
            I => byte_transmit_counter_4
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__26696\,
            I => byte_transmit_counter_4
        );

    \I__2991\ : InMux
    port map (
            O => \N__26683\,
            I => \N__26680\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__26680\,
            I => n23864
        );

    \I__2989\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26674\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__26674\,
            I => \N__26670\
        );

    \I__2987\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26667\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__26670\,
            I => \N__26664\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__26667\,
            I => data_out_frame_5_6
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__26664\,
            I => data_out_frame_5_6
        );

    \I__2983\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26655\
        );

    \I__2982\ : InMux
    port map (
            O => \N__26658\,
            I => \N__26652\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__26655\,
            I => \N__26649\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__26652\,
            I => data_out_frame_13_3
        );

    \I__2979\ : Odrv4
    port map (
            O => \N__26649\,
            I => data_out_frame_13_3
        );

    \I__2978\ : InMux
    port map (
            O => \N__26644\,
            I => \N__26641\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__26641\,
            I => n2184
        );

    \I__2976\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26635\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__26635\,
            I => n2182
        );

    \I__2974\ : InMux
    port map (
            O => \N__26632\,
            I => \N__26629\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__26629\,
            I => n2176
        );

    \I__2972\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26623\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__26623\,
            I => \N__26619\
        );

    \I__2970\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26616\
        );

    \I__2969\ : Span4Mux_v
    port map (
            O => \N__26619\,
            I => \N__26613\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__26616\,
            I => data_out_frame_29_3
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__26613\,
            I => data_out_frame_29_3
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__26608\,
            I => \N__26604\
        );

    \I__2965\ : InMux
    port map (
            O => \N__26607\,
            I => \N__26601\
        );

    \I__2964\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26598\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__26601\,
            I => \N__26595\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__26598\,
            I => data_out_frame_28_3
        );

    \I__2961\ : Odrv12
    port map (
            O => \N__26595\,
            I => data_out_frame_28_3
        );

    \I__2960\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26587\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__26587\,
            I => \N__26584\
        );

    \I__2958\ : Odrv4
    port map (
            O => \N__26584\,
            I => \c0.n26\
        );

    \I__2957\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26578\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__26578\,
            I => n2175
        );

    \I__2955\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26572\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__26572\,
            I => \N__26568\
        );

    \I__2953\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26565\
        );

    \I__2952\ : Span4Mux_h
    port map (
            O => \N__26568\,
            I => \N__26562\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__26565\,
            I => data_out_frame_7_5
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__26562\,
            I => data_out_frame_7_5
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__26557\,
            I => \N__26554\
        );

    \I__2948\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26551\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__26551\,
            I => \N__26548\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__26548\,
            I => \N__26545\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__26545\,
            I => \c0.n5_adj_4346\
        );

    \I__2944\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26538\
        );

    \I__2943\ : InMux
    port map (
            O => \N__26541\,
            I => \N__26535\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__26538\,
            I => \N__26532\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__26535\,
            I => \N__26527\
        );

    \I__2940\ : Span4Mux_v
    port map (
            O => \N__26532\,
            I => \N__26527\
        );

    \I__2939\ : Odrv4
    port map (
            O => \N__26527\,
            I => data_out_frame_9_7
        );

    \I__2938\ : IoInMux
    port map (
            O => \N__26524\,
            I => \N__26521\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__26521\,
            I => \N__26518\
        );

    \I__2936\ : IoSpan4Mux
    port map (
            O => \N__26518\,
            I => \N__26514\
        );

    \I__2935\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26511\
        );

    \I__2934\ : Span4Mux_s0_h
    port map (
            O => \N__26514\,
            I => \N__26508\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__26511\,
            I => \N__26505\
        );

    \I__2932\ : Span4Mux_s3_v
    port map (
            O => \N__26508\,
            I => \N__26500\
        );

    \I__2931\ : Span4Mux_s3_v
    port map (
            O => \N__26505\,
            I => \N__26500\
        );

    \I__2930\ : Sp12to4
    port map (
            O => \N__26500\,
            I => \N__26497\
        );

    \I__2929\ : Span12Mux_s10_h
    port map (
            O => \N__26497\,
            I => \N__26494\
        );

    \I__2928\ : Span12Mux_v
    port map (
            O => \N__26494\,
            I => \N__26490\
        );

    \I__2927\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26487\
        );

    \I__2926\ : Odrv12
    port map (
            O => \N__26490\,
            I => tx_o
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__26487\,
            I => tx_o
        );

    \I__2924\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26478\
        );

    \I__2923\ : InMux
    port map (
            O => \N__26481\,
            I => \N__26475\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__26478\,
            I => \N__26472\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__26475\,
            I => \N__26467\
        );

    \I__2920\ : Span4Mux_h
    port map (
            O => \N__26472\,
            I => \N__26467\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__26467\,
            I => \c0.data_out_frame_29__7__N_850\
        );

    \I__2918\ : InMux
    port map (
            O => \N__26464\,
            I => \N__26461\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__26461\,
            I => \N__26457\
        );

    \I__2916\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26454\
        );

    \I__2915\ : Span4Mux_v
    port map (
            O => \N__26457\,
            I => \N__26451\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__26454\,
            I => data_out_frame_11_4
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__26451\,
            I => data_out_frame_11_4
        );

    \I__2912\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26443\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__26443\,
            I => \N__26440\
        );

    \I__2910\ : Span4Mux_h
    port map (
            O => \N__26440\,
            I => \N__26437\
        );

    \I__2909\ : Odrv4
    port map (
            O => \N__26437\,
            I => \c0.n23881\
        );

    \I__2908\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26431\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__26431\,
            I => n2189
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__26428\,
            I => \N__26424\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__26427\,
            I => \N__26420\
        );

    \I__2904\ : InMux
    port map (
            O => \N__26424\,
            I => \N__26414\
        );

    \I__2903\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26411\
        );

    \I__2902\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26408\
        );

    \I__2901\ : InMux
    port map (
            O => \N__26419\,
            I => \N__26403\
        );

    \I__2900\ : InMux
    port map (
            O => \N__26418\,
            I => \N__26403\
        );

    \I__2899\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26400\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__26414\,
            I => \N__26397\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__26411\,
            I => \N__26394\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__26408\,
            I => \N__26389\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__26403\,
            I => \N__26389\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__26400\,
            I => encoder1_position_16
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__26397\,
            I => encoder1_position_16
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__26394\,
            I => encoder1_position_16
        );

    \I__2891\ : Odrv4
    port map (
            O => \N__26389\,
            I => encoder1_position_16
        );

    \I__2890\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26374\
        );

    \I__2889\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26374\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__26374\,
            I => data_out_frame_10_4
        );

    \I__2887\ : InMux
    port map (
            O => \N__26371\,
            I => \N__26368\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__26368\,
            I => \N__26365\
        );

    \I__2885\ : Span4Mux_v
    port map (
            O => \N__26365\,
            I => \N__26361\
        );

    \I__2884\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26358\
        );

    \I__2883\ : Span4Mux_v
    port map (
            O => \N__26361\,
            I => \N__26355\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__26358\,
            I => data_out_frame_7_2
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__26355\,
            I => data_out_frame_7_2
        );

    \I__2880\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26347\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__26347\,
            I => n2188
        );

    \I__2878\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26341\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__26341\,
            I => n2204
        );

    \I__2876\ : CascadeMux
    port map (
            O => \N__26338\,
            I => \c0.n6_adj_4310_cascade_\
        );

    \I__2875\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26329\
        );

    \I__2874\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26329\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__26329\,
            I => \c0.n22037\
        );

    \I__2872\ : InMux
    port map (
            O => \N__26326\,
            I => \N__26321\
        );

    \I__2871\ : InMux
    port map (
            O => \N__26325\,
            I => \N__26315\
        );

    \I__2870\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26315\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__26321\,
            I => \N__26312\
        );

    \I__2868\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26307\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__26315\,
            I => \N__26304\
        );

    \I__2866\ : Span4Mux_v
    port map (
            O => \N__26312\,
            I => \N__26301\
        );

    \I__2865\ : InMux
    port map (
            O => \N__26311\,
            I => \N__26298\
        );

    \I__2864\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26295\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__26307\,
            I => \N__26292\
        );

    \I__2862\ : Span4Mux_h
    port map (
            O => \N__26304\,
            I => \N__26289\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__26301\,
            I => encoder1_position_15
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__26298\,
            I => encoder1_position_15
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__26295\,
            I => encoder1_position_15
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__26292\,
            I => encoder1_position_15
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__26289\,
            I => encoder1_position_15
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__26278\,
            I => \N__26275\
        );

    \I__2855\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26269\
        );

    \I__2854\ : InMux
    port map (
            O => \N__26274\,
            I => \N__26269\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__26269\,
            I => data_out_frame_12_7
        );

    \I__2852\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26263\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__26263\,
            I => \N__26260\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__26260\,
            I => \N__26257\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__26257\,
            I => \c0.n11_adj_4360\
        );

    \I__2848\ : InMux
    port map (
            O => \N__26254\,
            I => \N__26251\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__26251\,
            I => n2197
        );

    \I__2846\ : InMux
    port map (
            O => \N__26248\,
            I => \N__26245\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__26245\,
            I => \N__26242\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__26242\,
            I => \c0.n5_adj_4227\
        );

    \I__2843\ : InMux
    port map (
            O => \N__26239\,
            I => \N__26233\
        );

    \I__2842\ : InMux
    port map (
            O => \N__26238\,
            I => \N__26233\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__26233\,
            I => data_out_frame_7_4
        );

    \I__2840\ : InMux
    port map (
            O => \N__26230\,
            I => \N__26227\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__26227\,
            I => \c0.n22116\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__26224\,
            I => \N__26221\
        );

    \I__2837\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26218\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__26218\,
            I => \N__26215\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__26215\,
            I => \c0.n6_adj_4308\
        );

    \I__2834\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26208\
        );

    \I__2833\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26205\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__26208\,
            I => \N__26200\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__26205\,
            I => \N__26200\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__26200\,
            I => data_out_frame_13_0
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__26197\,
            I => \N__26194\
        );

    \I__2828\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26191\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__26191\,
            I => \N__26188\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__26188\,
            I => \N__26185\
        );

    \I__2825\ : Span4Mux_v
    port map (
            O => \N__26185\,
            I => \N__26182\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__26182\,
            I => \c0.n11_adj_4424\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__26179\,
            I => \c0.n6_adj_4335_cascade_\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__26176\,
            I => \c0.n21229_cascade_\
        );

    \I__2821\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26170\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__26170\,
            I => \N__26167\
        );

    \I__2819\ : Span4Mux_v
    port map (
            O => \N__26167\,
            I => \N__26164\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__26164\,
            I => n2193
        );

    \I__2817\ : InMux
    port map (
            O => \N__26161\,
            I => \N__26158\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__26158\,
            I => \N__26155\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__26155\,
            I => \c0.n6_adj_4309\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__26152\,
            I => \N__26149\
        );

    \I__2813\ : InMux
    port map (
            O => \N__26149\,
            I => \N__26145\
        );

    \I__2812\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26142\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__26145\,
            I => data_out_frame_29_2
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__26142\,
            I => data_out_frame_29_2
        );

    \I__2809\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26134\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__26134\,
            I => \N__26131\
        );

    \I__2807\ : Span4Mux_v
    port map (
            O => \N__26131\,
            I => \N__26128\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__26128\,
            I => n2196
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__26125\,
            I => \c0.n13079_cascade_\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__26122\,
            I => \c0.n21305_cascade_\
        );

    \I__2803\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26116\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__26116\,
            I => \c0.data_out_frame_28_2\
        );

    \I__2801\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26110\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__26110\,
            I => \N__26107\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__26107\,
            I => \c0.n6_adj_4515\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__26104\,
            I => \c0.n12532_cascade_\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__26101\,
            I => \c0.n22126_cascade_\
        );

    \I__2796\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26095\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__26095\,
            I => \N__26092\
        );

    \I__2794\ : Span4Mux_v
    port map (
            O => \N__26092\,
            I => \N__26089\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__26089\,
            I => \c0.data_out_frame_28_4\
        );

    \I__2792\ : InMux
    port map (
            O => \N__26086\,
            I => \N__26082\
        );

    \I__2791\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26079\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__26082\,
            I => \N__26076\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__26079\,
            I => \quad_counter1.a_delay_counter_12\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__26076\,
            I => \quad_counter1.a_delay_counter_12\
        );

    \I__2787\ : InMux
    port map (
            O => \N__26071\,
            I => \N__26067\
        );

    \I__2786\ : InMux
    port map (
            O => \N__26070\,
            I => \N__26064\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__26067\,
            I => \quad_counter1.a_delay_counter_13\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__26064\,
            I => \quad_counter1.a_delay_counter_13\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__26059\,
            I => \N__26055\
        );

    \I__2782\ : InMux
    port map (
            O => \N__26058\,
            I => \N__26052\
        );

    \I__2781\ : InMux
    port map (
            O => \N__26055\,
            I => \N__26049\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__26052\,
            I => \quad_counter1.a_delay_counter_9\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__26049\,
            I => \quad_counter1.a_delay_counter_9\
        );

    \I__2778\ : InMux
    port map (
            O => \N__26044\,
            I => \N__26040\
        );

    \I__2777\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26037\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__26040\,
            I => \quad_counter1.a_delay_counter_6\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__26037\,
            I => \quad_counter1.a_delay_counter_6\
        );

    \I__2774\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__26029\,
            I => \N__26026\
        );

    \I__2772\ : Span4Mux_v
    port map (
            O => \N__26026\,
            I => \N__26023\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__26023\,
            I => \quad_counter1.n26\
        );

    \I__2770\ : SRMux
    port map (
            O => \N__26020\,
            I => \N__26017\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__26017\,
            I => \N__26013\
        );

    \I__2768\ : SRMux
    port map (
            O => \N__26016\,
            I => \N__26010\
        );

    \I__2767\ : Span4Mux_v
    port map (
            O => \N__26013\,
            I => \N__26005\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__26010\,
            I => \N__26005\
        );

    \I__2765\ : Sp12to4
    port map (
            O => \N__26005\,
            I => \N__26001\
        );

    \I__2764\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25998\
        );

    \I__2763\ : Odrv12
    port map (
            O => \N__26001\,
            I => \a_delay_counter_15__N_4124_adj_4547\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__25998\,
            I => \a_delay_counter_15__N_4124_adj_4547\
        );

    \I__2761\ : InMux
    port map (
            O => \N__25993\,
            I => \N__25988\
        );

    \I__2760\ : InMux
    port map (
            O => \N__25992\,
            I => \N__25983\
        );

    \I__2759\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25983\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__25988\,
            I => \N__25980\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__25983\,
            I => \N__25977\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__25980\,
            I => \N__25974\
        );

    \I__2755\ : Span4Mux_v
    port map (
            O => \N__25977\,
            I => \N__25971\
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__25974\,
            I => \quadA_delayed_adj_4542\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__25971\,
            I => \quadA_delayed_adj_4542\
        );

    \I__2752\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25960\
        );

    \I__2751\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25960\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__25960\,
            I => \N__25956\
        );

    \I__2749\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25953\
        );

    \I__2748\ : Span4Mux_v
    port map (
            O => \N__25956\,
            I => \N__25950\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__25953\,
            I => \N__25947\
        );

    \I__2746\ : Span4Mux_h
    port map (
            O => \N__25950\,
            I => \N__25943\
        );

    \I__2745\ : Span4Mux_v
    port map (
            O => \N__25947\,
            I => \N__25940\
        );

    \I__2744\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25937\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__25943\,
            I => \N__25934\
        );

    \I__2742\ : Sp12to4
    port map (
            O => \N__25940\,
            I => \N__25929\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__25937\,
            I => \N__25929\
        );

    \I__2740\ : Sp12to4
    port map (
            O => \N__25934\,
            I => \N__25924\
        );

    \I__2739\ : Span12Mux_h
    port map (
            O => \N__25929\,
            I => \N__25924\
        );

    \I__2738\ : Odrv12
    port map (
            O => \N__25924\,
            I => \PIN_12_c\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__25921\,
            I => \a_delay_counter_15__N_4124_adj_4547_cascade_\
        );

    \I__2736\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25915\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__25915\,
            I => \N__25912\
        );

    \I__2734\ : Span4Mux_h
    port map (
            O => \N__25912\,
            I => \N__25909\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__25909\,
            I => n9818
        );

    \I__2732\ : CEMux
    port map (
            O => \N__25906\,
            I => \N__25901\
        );

    \I__2731\ : CEMux
    port map (
            O => \N__25905\,
            I => \N__25898\
        );

    \I__2730\ : InMux
    port map (
            O => \N__25904\,
            I => \N__25895\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__25901\,
            I => n14228
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__25898\,
            I => n14228
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__25895\,
            I => n14228
        );

    \I__2726\ : InMux
    port map (
            O => \N__25888\,
            I => \quad_counter0.n19502\
        );

    \I__2725\ : InMux
    port map (
            O => \N__25885\,
            I => \N__25882\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__25882\,
            I => \c0.n24_adj_4502\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__25879\,
            I => \c0.n18_adj_4414_cascade_\
        );

    \I__2722\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25873\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__25873\,
            I => \c0.n13360\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__25870\,
            I => \c0.n23550_cascade_\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__25867\,
            I => \c0.n22_adj_4503_cascade_\
        );

    \I__2718\ : InMux
    port map (
            O => \N__25864\,
            I => \N__25861\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__25861\,
            I => \c0.n26_adj_4504\
        );

    \I__2716\ : InMux
    port map (
            O => \N__25858\,
            I => \N__25855\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__25855\,
            I => \N__25852\
        );

    \I__2714\ : Span4Mux_h
    port map (
            O => \N__25852\,
            I => \N__25849\
        );

    \I__2713\ : Span4Mux_v
    port map (
            O => \N__25849\,
            I => \N__25846\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__25846\,
            I => \N__25843\
        );

    \I__2711\ : Odrv4
    port map (
            O => \N__25843\,
            I => \c0.n26_adj_4517\
        );

    \I__2710\ : InMux
    port map (
            O => \N__25840\,
            I => \quad_counter0.n19493\
        );

    \I__2709\ : InMux
    port map (
            O => \N__25837\,
            I => \quad_counter0.n19494\
        );

    \I__2708\ : InMux
    port map (
            O => \N__25834\,
            I => \bfn_10_25_0_\
        );

    \I__2707\ : InMux
    port map (
            O => \N__25831\,
            I => \quad_counter0.n19496\
        );

    \I__2706\ : InMux
    port map (
            O => \N__25828\,
            I => \quad_counter0.n19497\
        );

    \I__2705\ : InMux
    port map (
            O => \N__25825\,
            I => \quad_counter0.n19498\
        );

    \I__2704\ : InMux
    port map (
            O => \N__25822\,
            I => \quad_counter0.n19499\
        );

    \I__2703\ : InMux
    port map (
            O => \N__25819\,
            I => \quad_counter0.n19500\
        );

    \I__2702\ : InMux
    port map (
            O => \N__25816\,
            I => \quad_counter0.n19501\
        );

    \I__2701\ : InMux
    port map (
            O => \N__25813\,
            I => \quad_counter0.n19485\
        );

    \I__2700\ : InMux
    port map (
            O => \N__25810\,
            I => \quad_counter0.n19486\
        );

    \I__2699\ : InMux
    port map (
            O => \N__25807\,
            I => \quad_counter0.n19487\
        );

    \I__2698\ : CEMux
    port map (
            O => \N__25804\,
            I => \N__25800\
        );

    \I__2697\ : CEMux
    port map (
            O => \N__25803\,
            I => \N__25797\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__25800\,
            I => \N__25793\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__25797\,
            I => \N__25790\
        );

    \I__2694\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25787\
        );

    \I__2693\ : Odrv4
    port map (
            O => \N__25793\,
            I => n14198
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__25790\,
            I => n14198
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__25787\,
            I => n14198
        );

    \I__2690\ : SRMux
    port map (
            O => \N__25780\,
            I => \N__25777\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__25777\,
            I => \N__25773\
        );

    \I__2688\ : SRMux
    port map (
            O => \N__25776\,
            I => \N__25770\
        );

    \I__2687\ : Span4Mux_h
    port map (
            O => \N__25773\,
            I => \N__25766\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__25770\,
            I => \N__25763\
        );

    \I__2685\ : InMux
    port map (
            O => \N__25769\,
            I => \N__25760\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__25766\,
            I => \b_delay_counter_15__N_4141\
        );

    \I__2683\ : Odrv4
    port map (
            O => \N__25763\,
            I => \b_delay_counter_15__N_4141\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__25760\,
            I => \b_delay_counter_15__N_4141\
        );

    \I__2681\ : InMux
    port map (
            O => \N__25753\,
            I => \bfn_10_24_0_\
        );

    \I__2680\ : InMux
    port map (
            O => \N__25750\,
            I => \quad_counter0.n19488\
        );

    \I__2679\ : InMux
    port map (
            O => \N__25747\,
            I => \quad_counter0.n19489\
        );

    \I__2678\ : InMux
    port map (
            O => \N__25744\,
            I => \quad_counter0.n19490\
        );

    \I__2677\ : InMux
    port map (
            O => \N__25741\,
            I => \quad_counter0.n19491\
        );

    \I__2676\ : InMux
    port map (
            O => \N__25738\,
            I => \quad_counter0.n19492\
        );

    \I__2675\ : InMux
    port map (
            O => \N__25735\,
            I => \quad_counter0.n19476\
        );

    \I__2674\ : InMux
    port map (
            O => \N__25732\,
            I => \quad_counter0.n19477\
        );

    \I__2673\ : InMux
    port map (
            O => \N__25729\,
            I => \quad_counter0.n19478\
        );

    \I__2672\ : InMux
    port map (
            O => \N__25726\,
            I => \quad_counter0.n19479\
        );

    \I__2671\ : InMux
    port map (
            O => \N__25723\,
            I => \bfn_10_23_0_\
        );

    \I__2670\ : InMux
    port map (
            O => \N__25720\,
            I => \quad_counter0.n19481\
        );

    \I__2669\ : InMux
    port map (
            O => \N__25717\,
            I => \quad_counter0.n19482\
        );

    \I__2668\ : InMux
    port map (
            O => \N__25714\,
            I => \quad_counter0.n19483\
        );

    \I__2667\ : InMux
    port map (
            O => \N__25711\,
            I => \quad_counter0.n19484\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__25708\,
            I => \n24100_cascade_\
        );

    \I__2665\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25702\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__25702\,
            I => n16706
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__25699\,
            I => \c0.tx.n23985_cascade_\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__25696\,
            I => \c0.tx.n31_adj_4216_cascade_\
        );

    \I__2661\ : InMux
    port map (
            O => \N__25693\,
            I => \N__25690\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__25690\,
            I => n187
        );

    \I__2659\ : InMux
    port map (
            O => \N__25687\,
            I => \bfn_10_22_0_\
        );

    \I__2658\ : InMux
    port map (
            O => \N__25684\,
            I => \quad_counter0.n19473\
        );

    \I__2657\ : InMux
    port map (
            O => \N__25681\,
            I => \quad_counter0.n19474\
        );

    \I__2656\ : InMux
    port map (
            O => \N__25678\,
            I => \quad_counter0.n19475\
        );

    \I__2655\ : InMux
    port map (
            O => \N__25675\,
            I => \N__25672\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__25672\,
            I => \N__25669\
        );

    \I__2653\ : Span4Mux_h
    port map (
            O => \N__25669\,
            I => \N__25666\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__25666\,
            I => \N__25663\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__25663\,
            I => n10_adj_4536
        );

    \I__2650\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25657\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__25657\,
            I => \c0.n5_adj_4422\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__25654\,
            I => \N__25651\
        );

    \I__2647\ : InMux
    port map (
            O => \N__25651\,
            I => \N__25648\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__25648\,
            I => \c0.n24059\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__25645\,
            I => \c0.n23850_cascade_\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__25642\,
            I => \n23852_cascade_\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__25639\,
            I => \N__25630\
        );

    \I__2642\ : InMux
    port map (
            O => \N__25638\,
            I => \N__25627\
        );

    \I__2641\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25623\
        );

    \I__2640\ : InMux
    port map (
            O => \N__25636\,
            I => \N__25620\
        );

    \I__2639\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25617\
        );

    \I__2638\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25614\
        );

    \I__2637\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25611\
        );

    \I__2636\ : InMux
    port map (
            O => \N__25630\,
            I => \N__25608\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__25627\,
            I => \N__25604\
        );

    \I__2634\ : InMux
    port map (
            O => \N__25626\,
            I => \N__25601\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__25623\,
            I => \N__25596\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__25620\,
            I => \N__25596\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__25617\,
            I => \N__25591\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__25614\,
            I => \N__25591\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__25611\,
            I => \N__25586\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__25608\,
            I => \N__25583\
        );

    \I__2627\ : InMux
    port map (
            O => \N__25607\,
            I => \N__25580\
        );

    \I__2626\ : Span4Mux_h
    port map (
            O => \N__25604\,
            I => \N__25577\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__25601\,
            I => \N__25570\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__25596\,
            I => \N__25570\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__25591\,
            I => \N__25570\
        );

    \I__2622\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25565\
        );

    \I__2621\ : InMux
    port map (
            O => \N__25589\,
            I => \N__25565\
        );

    \I__2620\ : Span4Mux_v
    port map (
            O => \N__25586\,
            I => \N__25558\
        );

    \I__2619\ : Span4Mux_v
    port map (
            O => \N__25583\,
            I => \N__25558\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__25580\,
            I => \N__25558\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__25577\,
            I => byte_transmit_counter_3
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__25570\,
            I => byte_transmit_counter_3
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__25565\,
            I => byte_transmit_counter_3
        );

    \I__2614\ : Odrv4
    port map (
            O => \N__25558\,
            I => byte_transmit_counter_3
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__25549\,
            I => \n10_adj_4537_cascade_\
        );

    \I__2612\ : InMux
    port map (
            O => \N__25546\,
            I => \N__25543\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__25543\,
            I => n24110
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__25540\,
            I => \N__25536\
        );

    \I__2609\ : InMux
    port map (
            O => \N__25539\,
            I => \N__25531\
        );

    \I__2608\ : InMux
    port map (
            O => \N__25536\,
            I => \N__25531\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__25531\,
            I => \r_Tx_Data_0\
        );

    \I__2606\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25525\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__25525\,
            I => n24195
        );

    \I__2604\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25518\
        );

    \I__2603\ : InMux
    port map (
            O => \N__25521\,
            I => \N__25515\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__25518\,
            I => \N__25512\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__25515\,
            I => \r_Tx_Data_5\
        );

    \I__2600\ : Odrv12
    port map (
            O => \N__25512\,
            I => \r_Tx_Data_5\
        );

    \I__2599\ : InMux
    port map (
            O => \N__25507\,
            I => \N__25504\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__25504\,
            I => \N__25500\
        );

    \I__2597\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25497\
        );

    \I__2596\ : Span4Mux_v
    port map (
            O => \N__25500\,
            I => \N__25494\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__25497\,
            I => \r_Tx_Data_4\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__25494\,
            I => \r_Tx_Data_4\
        );

    \I__2593\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25486\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__25486\,
            I => n10_adj_4533
        );

    \I__2591\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25479\
        );

    \I__2590\ : InMux
    port map (
            O => \N__25482\,
            I => \N__25476\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__25479\,
            I => data_out_frame_9_2
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__25476\,
            I => data_out_frame_9_2
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__25471\,
            I => \c0.n24180_cascade_\
        );

    \I__2586\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25465\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__25465\,
            I => n24106
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__25462\,
            I => \N__25459\
        );

    \I__2583\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25453\
        );

    \I__2582\ : InMux
    port map (
            O => \N__25458\,
            I => \N__25453\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__25453\,
            I => data_out_frame_7_0
        );

    \I__2580\ : InMux
    port map (
            O => \N__25450\,
            I => \N__25444\
        );

    \I__2579\ : InMux
    port map (
            O => \N__25449\,
            I => \N__25444\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__25444\,
            I => data_out_frame_6_0
        );

    \I__2577\ : InMux
    port map (
            O => \N__25441\,
            I => \bfn_10_17_0_\
        );

    \I__2576\ : InMux
    port map (
            O => \N__25438\,
            I => \N__25435\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__25435\,
            I => \N__25432\
        );

    \I__2574\ : Odrv4
    port map (
            O => \N__25432\,
            I => n2174
        );

    \I__2573\ : InMux
    port map (
            O => \N__25429\,
            I => \N__25426\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__25426\,
            I => \N__25422\
        );

    \I__2571\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25419\
        );

    \I__2570\ : Span4Mux_h
    port map (
            O => \N__25422\,
            I => \N__25416\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__25419\,
            I => data_out_frame_0_4
        );

    \I__2568\ : Odrv4
    port map (
            O => \N__25416\,
            I => data_out_frame_0_4
        );

    \I__2567\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25407\
        );

    \I__2566\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25404\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__25407\,
            I => data_out_frame_13_5
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__25404\,
            I => data_out_frame_13_5
        );

    \I__2563\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25393\
        );

    \I__2562\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25393\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__25393\,
            I => data_out_frame_9_3
        );

    \I__2560\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25387\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__25387\,
            I => \c0.n24171\
        );

    \I__2558\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25381\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__25381\,
            I => \c0.n24174\
        );

    \I__2556\ : InMux
    port map (
            O => \N__25378\,
            I => \N__25375\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__25375\,
            I => \c0.n23856\
        );

    \I__2554\ : InMux
    port map (
            O => \N__25372\,
            I => \N__25369\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__25369\,
            I => \N__25366\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__25366\,
            I => n24108
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__25363\,
            I => \n23858_cascade_\
        );

    \I__2550\ : InMux
    port map (
            O => \N__25360\,
            I => \bfn_10_16_0_\
        );

    \I__2549\ : InMux
    port map (
            O => \N__25357\,
            I => \quad_counter1.n19572\
        );

    \I__2548\ : InMux
    port map (
            O => \N__25354\,
            I => \quad_counter1.n19573\
        );

    \I__2547\ : InMux
    port map (
            O => \N__25351\,
            I => \N__25348\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__25348\,
            I => \N__25345\
        );

    \I__2545\ : Odrv12
    port map (
            O => \N__25345\,
            I => n2179
        );

    \I__2544\ : InMux
    port map (
            O => \N__25342\,
            I => \quad_counter1.n19574\
        );

    \I__2543\ : InMux
    port map (
            O => \N__25339\,
            I => \quad_counter1.n19575\
        );

    \I__2542\ : InMux
    port map (
            O => \N__25336\,
            I => \N__25333\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__25333\,
            I => n2177
        );

    \I__2540\ : InMux
    port map (
            O => \N__25330\,
            I => \quad_counter1.n19576\
        );

    \I__2539\ : InMux
    port map (
            O => \N__25327\,
            I => \quad_counter1.n19577\
        );

    \I__2538\ : InMux
    port map (
            O => \N__25324\,
            I => \quad_counter1.n19578\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__25321\,
            I => \N__25303\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__25320\,
            I => \N__25299\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__25319\,
            I => \N__25295\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__25318\,
            I => \N__25290\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__25317\,
            I => \N__25286\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__25316\,
            I => \N__25282\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__25315\,
            I => \N__25278\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__25314\,
            I => \N__25275\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__25313\,
            I => \N__25271\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__25312\,
            I => \N__25267\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__25311\,
            I => \N__25263\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__25310\,
            I => \N__25258\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__25309\,
            I => \N__25255\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__25308\,
            I => \N__25252\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__25307\,
            I => \N__25247\
        );

    \I__2522\ : InMux
    port map (
            O => \N__25306\,
            I => \N__25243\
        );

    \I__2521\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25230\
        );

    \I__2520\ : InMux
    port map (
            O => \N__25302\,
            I => \N__25230\
        );

    \I__2519\ : InMux
    port map (
            O => \N__25299\,
            I => \N__25230\
        );

    \I__2518\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25230\
        );

    \I__2517\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25230\
        );

    \I__2516\ : InMux
    port map (
            O => \N__25294\,
            I => \N__25230\
        );

    \I__2515\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25213\
        );

    \I__2514\ : InMux
    port map (
            O => \N__25290\,
            I => \N__25213\
        );

    \I__2513\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25213\
        );

    \I__2512\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25213\
        );

    \I__2511\ : InMux
    port map (
            O => \N__25285\,
            I => \N__25213\
        );

    \I__2510\ : InMux
    port map (
            O => \N__25282\,
            I => \N__25213\
        );

    \I__2509\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25213\
        );

    \I__2508\ : InMux
    port map (
            O => \N__25278\,
            I => \N__25213\
        );

    \I__2507\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25196\
        );

    \I__2506\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25196\
        );

    \I__2505\ : InMux
    port map (
            O => \N__25271\,
            I => \N__25196\
        );

    \I__2504\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25196\
        );

    \I__2503\ : InMux
    port map (
            O => \N__25267\,
            I => \N__25196\
        );

    \I__2502\ : InMux
    port map (
            O => \N__25266\,
            I => \N__25196\
        );

    \I__2501\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25196\
        );

    \I__2500\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25196\
        );

    \I__2499\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25187\
        );

    \I__2498\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25187\
        );

    \I__2497\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25187\
        );

    \I__2496\ : InMux
    port map (
            O => \N__25252\,
            I => \N__25187\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__25251\,
            I => \N__25183\
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__25250\,
            I => \N__25180\
        );

    \I__2493\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25174\
        );

    \I__2492\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25174\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__25243\,
            I => \N__25165\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__25230\,
            I => \N__25165\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__25213\,
            I => \N__25165\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__25196\,
            I => \N__25165\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__25187\,
            I => \N__25162\
        );

    \I__2486\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25153\
        );

    \I__2485\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25153\
        );

    \I__2484\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25153\
        );

    \I__2483\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25153\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__25174\,
            I => \N__25150\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__25165\,
            I => \N__25143\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__25162\,
            I => \N__25143\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__25153\,
            I => \N__25143\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__25150\,
            I => \N__25140\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__25143\,
            I => \N__25137\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__25140\,
            I => \quad_counter1.n2140\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__25137\,
            I => \quad_counter1.n2140\
        );

    \I__2474\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25129\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__25129\,
            I => \N__25126\
        );

    \I__2472\ : Odrv12
    port map (
            O => \N__25126\,
            I => n2191
        );

    \I__2471\ : InMux
    port map (
            O => \N__25123\,
            I => \quad_counter1.n19562\
        );

    \I__2470\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25117\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__25117\,
            I => n2190
        );

    \I__2468\ : InMux
    port map (
            O => \N__25114\,
            I => \bfn_10_15_0_\
        );

    \I__2467\ : InMux
    port map (
            O => \N__25111\,
            I => \quad_counter1.n19564\
        );

    \I__2466\ : InMux
    port map (
            O => \N__25108\,
            I => \quad_counter1.n19565\
        );

    \I__2465\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25102\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__25102\,
            I => \N__25099\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__25099\,
            I => n2187
        );

    \I__2462\ : InMux
    port map (
            O => \N__25096\,
            I => \quad_counter1.n19566\
        );

    \I__2461\ : InMux
    port map (
            O => \N__25093\,
            I => \quad_counter1.n19567\
        );

    \I__2460\ : InMux
    port map (
            O => \N__25090\,
            I => \quad_counter1.n19568\
        );

    \I__2459\ : InMux
    port map (
            O => \N__25087\,
            I => \quad_counter1.n19569\
        );

    \I__2458\ : InMux
    port map (
            O => \N__25084\,
            I => \N__25081\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__25081\,
            I => \N__25078\
        );

    \I__2456\ : Odrv12
    port map (
            O => \N__25078\,
            I => n2183
        );

    \I__2455\ : InMux
    port map (
            O => \N__25075\,
            I => \quad_counter1.n19570\
        );

    \I__2454\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25069\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__25069\,
            I => \N__25066\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__25066\,
            I => n2200
        );

    \I__2451\ : InMux
    port map (
            O => \N__25063\,
            I => \quad_counter1.n19553\
        );

    \I__2450\ : InMux
    port map (
            O => \N__25060\,
            I => \N__25057\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__25057\,
            I => n2199
        );

    \I__2448\ : InMux
    port map (
            O => \N__25054\,
            I => \quad_counter1.n19554\
        );

    \I__2447\ : InMux
    port map (
            O => \N__25051\,
            I => \bfn_10_14_0_\
        );

    \I__2446\ : InMux
    port map (
            O => \N__25048\,
            I => \quad_counter1.n19556\
        );

    \I__2445\ : InMux
    port map (
            O => \N__25045\,
            I => \quad_counter1.n19557\
        );

    \I__2444\ : InMux
    port map (
            O => \N__25042\,
            I => \quad_counter1.n19558\
        );

    \I__2443\ : InMux
    port map (
            O => \N__25039\,
            I => \quad_counter1.n19559\
        );

    \I__2442\ : InMux
    port map (
            O => \N__25036\,
            I => \quad_counter1.n19560\
        );

    \I__2441\ : InMux
    port map (
            O => \N__25033\,
            I => \quad_counter1.n19561\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__25030\,
            I => \c0.n22048_cascade_\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__25027\,
            I => \N__25022\
        );

    \I__2438\ : InMux
    port map (
            O => \N__25026\,
            I => \N__25018\
        );

    \I__2437\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25011\
        );

    \I__2436\ : InMux
    port map (
            O => \N__25022\,
            I => \N__25011\
        );

    \I__2435\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25011\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__25018\,
            I => encoder1_position_0
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__25011\,
            I => encoder1_position_0
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__25006\,
            I => \N__25003\
        );

    \I__2431\ : InMux
    port map (
            O => \N__25003\,
            I => \N__25000\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__25000\,
            I => \N__24997\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__24997\,
            I => \quad_counter1.count_direction\
        );

    \I__2428\ : InMux
    port map (
            O => \N__24994\,
            I => \N__24991\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__24991\,
            I => n2205
        );

    \I__2426\ : InMux
    port map (
            O => \N__24988\,
            I => \quad_counter1.n19548\
        );

    \I__2425\ : InMux
    port map (
            O => \N__24985\,
            I => \quad_counter1.n19549\
        );

    \I__2424\ : InMux
    port map (
            O => \N__24982\,
            I => \N__24979\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__24979\,
            I => \N__24976\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__24976\,
            I => n2203
        );

    \I__2421\ : InMux
    port map (
            O => \N__24973\,
            I => \quad_counter1.n19550\
        );

    \I__2420\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24967\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__24967\,
            I => \N__24964\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__24964\,
            I => n2202
        );

    \I__2417\ : InMux
    port map (
            O => \N__24961\,
            I => \quad_counter1.n19551\
        );

    \I__2416\ : InMux
    port map (
            O => \N__24958\,
            I => \quad_counter1.n19552\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__24955\,
            I => \N__24950\
        );

    \I__2414\ : InMux
    port map (
            O => \N__24954\,
            I => \N__24947\
        );

    \I__2413\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24942\
        );

    \I__2412\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24942\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__24947\,
            I => \N__24939\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__24942\,
            I => \N__24934\
        );

    \I__2409\ : Span4Mux_h
    port map (
            O => \N__24939\,
            I => \N__24931\
        );

    \I__2408\ : InMux
    port map (
            O => \N__24938\,
            I => \N__24926\
        );

    \I__2407\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24926\
        );

    \I__2406\ : Odrv12
    port map (
            O => \N__24934\,
            I => \A_filtered_adj_4538\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__24931\,
            I => \A_filtered_adj_4538\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__24926\,
            I => \A_filtered_adj_4538\
        );

    \I__2403\ : InMux
    port map (
            O => \N__24919\,
            I => \N__24915\
        );

    \I__2402\ : InMux
    port map (
            O => \N__24918\,
            I => \N__24912\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__24915\,
            I => \N__24906\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__24912\,
            I => \N__24906\
        );

    \I__2399\ : InMux
    port map (
            O => \N__24911\,
            I => \N__24903\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__24906\,
            I => \quad_counter1.B_delayed\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__24903\,
            I => \quad_counter1.B_delayed\
        );

    \I__2396\ : InMux
    port map (
            O => \N__24898\,
            I => \N__24895\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__24895\,
            I => \N__24892\
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__24892\,
            I => n39_adj_4545
        );

    \I__2393\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24884\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__24888\,
            I => \N__24881\
        );

    \I__2391\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24878\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__24884\,
            I => \N__24875\
        );

    \I__2389\ : InMux
    port map (
            O => \N__24881\,
            I => \N__24872\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__24878\,
            I => \N__24869\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__24875\,
            I => \N__24866\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__24872\,
            I => a_delay_counter_0_adj_4540
        );

    \I__2385\ : Odrv12
    port map (
            O => \N__24869\,
            I => a_delay_counter_0_adj_4540
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__24866\,
            I => a_delay_counter_0_adj_4540
        );

    \I__2383\ : CascadeMux
    port map (
            O => \N__24859\,
            I => \N__24855\
        );

    \I__2382\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24852\
        );

    \I__2381\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24849\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__24852\,
            I => \quad_counter1.a_delay_counter_10\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__24849\,
            I => \quad_counter1.a_delay_counter_10\
        );

    \I__2378\ : InMux
    port map (
            O => \N__24844\,
            I => \quad_counter1.n19527\
        );

    \I__2377\ : InMux
    port map (
            O => \N__24841\,
            I => \N__24837\
        );

    \I__2376\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24834\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__24837\,
            I => \quad_counter1.a_delay_counter_11\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__24834\,
            I => \quad_counter1.a_delay_counter_11\
        );

    \I__2373\ : InMux
    port map (
            O => \N__24829\,
            I => \quad_counter1.n19528\
        );

    \I__2372\ : InMux
    port map (
            O => \N__24826\,
            I => \quad_counter1.n19529\
        );

    \I__2371\ : InMux
    port map (
            O => \N__24823\,
            I => \quad_counter1.n19530\
        );

    \I__2370\ : InMux
    port map (
            O => \N__24820\,
            I => \N__24816\
        );

    \I__2369\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24813\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__24816\,
            I => \quad_counter1.a_delay_counter_14\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__24813\,
            I => \quad_counter1.a_delay_counter_14\
        );

    \I__2366\ : InMux
    port map (
            O => \N__24808\,
            I => \quad_counter1.n19531\
        );

    \I__2365\ : InMux
    port map (
            O => \N__24805\,
            I => \quad_counter1.n19532\
        );

    \I__2364\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24798\
        );

    \I__2363\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24795\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__24798\,
            I => \quad_counter1.a_delay_counter_15\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__24795\,
            I => \quad_counter1.a_delay_counter_15\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__24790\,
            I => \N__24786\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__24789\,
            I => \N__24783\
        );

    \I__2358\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24780\
        );

    \I__2357\ : InMux
    port map (
            O => \N__24783\,
            I => \N__24777\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__24780\,
            I => \N__24774\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__24777\,
            I => data_out_frame_11_6
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__24774\,
            I => data_out_frame_11_6
        );

    \I__2353\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24765\
        );

    \I__2352\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24762\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__24765\,
            I => \N__24757\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24757\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__24757\,
            I => \quad_counter1.a_delay_counter_1\
        );

    \I__2348\ : InMux
    port map (
            O => \N__24754\,
            I => \quad_counter1.n19518\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__24751\,
            I => \N__24747\
        );

    \I__2346\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24744\
        );

    \I__2345\ : InMux
    port map (
            O => \N__24747\,
            I => \N__24741\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__24744\,
            I => \quad_counter1.a_delay_counter_2\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__24741\,
            I => \quad_counter1.a_delay_counter_2\
        );

    \I__2342\ : InMux
    port map (
            O => \N__24736\,
            I => \quad_counter1.n19519\
        );

    \I__2341\ : InMux
    port map (
            O => \N__24733\,
            I => \N__24729\
        );

    \I__2340\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24726\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__24729\,
            I => \quad_counter1.a_delay_counter_3\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__24726\,
            I => \quad_counter1.a_delay_counter_3\
        );

    \I__2337\ : InMux
    port map (
            O => \N__24721\,
            I => \quad_counter1.n19520\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__24718\,
            I => \N__24714\
        );

    \I__2335\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24711\
        );

    \I__2334\ : InMux
    port map (
            O => \N__24714\,
            I => \N__24708\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__24711\,
            I => \quad_counter1.a_delay_counter_4\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__24708\,
            I => \quad_counter1.a_delay_counter_4\
        );

    \I__2331\ : InMux
    port map (
            O => \N__24703\,
            I => \quad_counter1.n19521\
        );

    \I__2330\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24696\
        );

    \I__2329\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24693\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__24696\,
            I => \quad_counter1.a_delay_counter_5\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__24693\,
            I => \quad_counter1.a_delay_counter_5\
        );

    \I__2326\ : InMux
    port map (
            O => \N__24688\,
            I => \quad_counter1.n19522\
        );

    \I__2325\ : InMux
    port map (
            O => \N__24685\,
            I => \quad_counter1.n19523\
        );

    \I__2324\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24678\
        );

    \I__2323\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24675\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__24678\,
            I => \N__24672\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__24675\,
            I => \quad_counter1.a_delay_counter_7\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__24672\,
            I => \quad_counter1.a_delay_counter_7\
        );

    \I__2319\ : InMux
    port map (
            O => \N__24667\,
            I => \quad_counter1.n19524\
        );

    \I__2318\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24660\
        );

    \I__2317\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24657\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__24660\,
            I => \N__24654\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__24657\,
            I => \quad_counter1.a_delay_counter_8\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__24654\,
            I => \quad_counter1.a_delay_counter_8\
        );

    \I__2313\ : InMux
    port map (
            O => \N__24649\,
            I => \bfn_10_10_0_\
        );

    \I__2312\ : InMux
    port map (
            O => \N__24646\,
            I => \quad_counter1.n19526\
        );

    \I__2311\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24640\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24636\
        );

    \I__2309\ : InMux
    port map (
            O => \N__24639\,
            I => \N__24633\
        );

    \I__2308\ : Span4Mux_h
    port map (
            O => \N__24636\,
            I => \N__24630\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__24633\,
            I => \r_Tx_Data_6\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__24630\,
            I => \r_Tx_Data_6\
        );

    \I__2305\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24622\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__24622\,
            I => \N__24618\
        );

    \I__2303\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24615\
        );

    \I__2302\ : Span4Mux_h
    port map (
            O => \N__24618\,
            I => \N__24612\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__24615\,
            I => \r_Tx_Data_2\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__24612\,
            I => \r_Tx_Data_2\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__24607\,
            I => \b_delay_counter_15__N_4141_cascade_\
        );

    \I__2298\ : InMux
    port map (
            O => \N__24604\,
            I => \bfn_10_9_0_\
        );

    \I__2297\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24597\
        );

    \I__2296\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24594\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__24597\,
            I => data_out_frame_0_2
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__24594\,
            I => data_out_frame_0_2
        );

    \I__2293\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24586\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__24586\,
            I => \c0.n6_adj_4521\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__24583\,
            I => \c0.n23859_cascade_\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__24580\,
            I => \n23861_cascade_\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__24577\,
            I => \N__24574\
        );

    \I__2288\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24571\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__24571\,
            I => \N__24568\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__24568\,
            I => n10_adj_4534
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__24565\,
            I => \N__24562\
        );

    \I__2284\ : InMux
    port map (
            O => \N__24562\,
            I => \N__24559\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__24559\,
            I => \c0.n5_adj_4522\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__24556\,
            I => \N__24553\
        );

    \I__2281\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24547\
        );

    \I__2280\ : InMux
    port map (
            O => \N__24552\,
            I => \N__24547\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__24547\,
            I => data_out_frame_6_2
        );

    \I__2278\ : InMux
    port map (
            O => \N__24544\,
            I => \N__24541\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__24541\,
            I => \c0.n24007\
        );

    \I__2276\ : InMux
    port map (
            O => \N__24538\,
            I => \N__24535\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__24535\,
            I => \c0.n6\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__24532\,
            I => \N__24529\
        );

    \I__2273\ : InMux
    port map (
            O => \N__24529\,
            I => \N__24526\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__24526\,
            I => \c0.n11_adj_4348\
        );

    \I__2271\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24520\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__24520\,
            I => \N__24517\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__24517\,
            I => n24102
        );

    \I__2268\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24511\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__24511\,
            I => \c0.n24047\
        );

    \I__2266\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24505\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__24505\,
            I => \c0.n5_adj_4358\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__24502\,
            I => \N__24499\
        );

    \I__2263\ : InMux
    port map (
            O => \N__24499\,
            I => \N__24493\
        );

    \I__2262\ : InMux
    port map (
            O => \N__24498\,
            I => \N__24493\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__24493\,
            I => data_out_frame_6_7
        );

    \I__2260\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24486\
        );

    \I__2259\ : InMux
    port map (
            O => \N__24489\,
            I => \N__24483\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__24486\,
            I => data_out_frame_0_3
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__24483\,
            I => data_out_frame_0_3
        );

    \I__2256\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24475\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__24475\,
            I => \N__24472\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__24472\,
            I => \c0.n24011\
        );

    \I__2253\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24466\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__24466\,
            I => \c0.n11_adj_4355\
        );

    \I__2251\ : InMux
    port map (
            O => \N__24463\,
            I => \N__24460\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__24460\,
            I => n23846
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__24457\,
            I => \n24114_cascade_\
        );

    \I__2248\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24451\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__24451\,
            I => \N__24448\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__24448\,
            I => \N__24445\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__24445\,
            I => n10
        );

    \I__2244\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24439\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__24439\,
            I => \N__24436\
        );

    \I__2242\ : Span4Mux_h
    port map (
            O => \N__24436\,
            I => \N__24433\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__24433\,
            I => \c0.n23895\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__24430\,
            I => \c0.n24051_cascade_\
        );

    \I__2239\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24424\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__24424\,
            I => \c0.n23844\
        );

    \I__2237\ : InMux
    port map (
            O => \N__24421\,
            I => \N__24418\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__24418\,
            I => \N__24415\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__24415\,
            I => \c0.n23847\
        );

    \I__2234\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24409\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__24409\,
            I => n24112
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__24406\,
            I => \n23849_cascade_\
        );

    \I__2231\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24399\
        );

    \I__2230\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24396\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__24399\,
            I => \N__24393\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__24396\,
            I => data_out_frame_10_3
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__24393\,
            I => data_out_frame_10_3
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__24388\,
            I => \c0.n24159_cascade_\
        );

    \I__2225\ : InMux
    port map (
            O => \N__24385\,
            I => \N__24382\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__24382\,
            I => \N__24379\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__24379\,
            I => \c0.n24162\
        );

    \I__2222\ : InMux
    port map (
            O => \N__24376\,
            I => \N__24373\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__24373\,
            I => \N__24370\
        );

    \I__2220\ : Odrv12
    port map (
            O => \N__24370\,
            I => n26
        );

    \I__2219\ : CascadeMux
    port map (
            O => \N__24367\,
            I => \n24118_cascade_\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__24364\,
            I => \c0.n23950_cascade_\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__24361\,
            I => \c0.n24147_cascade_\
        );

    \I__2216\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24355\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__24355\,
            I => \N__24352\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__24352\,
            I => \c0.n23882\
        );

    \I__2213\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24346\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__24346\,
            I => n24150
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__24343\,
            I => \n24097_cascade_\
        );

    \I__2210\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24337\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__24337\,
            I => n24117
        );

    \I__2208\ : InMux
    port map (
            O => \N__24334\,
            I => \quad_counter1.n19517\
        );

    \I__2207\ : InMux
    port map (
            O => \N__24331\,
            I => \N__24327\
        );

    \I__2206\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24324\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__24327\,
            I => \N__24321\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__24324\,
            I => \quad_counter1.b_delay_counter_15\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__24321\,
            I => \quad_counter1.b_delay_counter_15\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__24316\,
            I => \N__24312\
        );

    \I__2201\ : CEMux
    port map (
            O => \N__24315\,
            I => \N__24308\
        );

    \I__2200\ : InMux
    port map (
            O => \N__24312\,
            I => \N__24305\
        );

    \I__2199\ : CEMux
    port map (
            O => \N__24311\,
            I => \N__24302\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__24308\,
            I => \N__24299\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24294\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24294\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__24299\,
            I => \N__24291\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__24294\,
            I => \N__24288\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__24291\,
            I => n14377
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__24288\,
            I => n14377
        );

    \I__2191\ : SRMux
    port map (
            O => \N__24283\,
            I => \N__24279\
        );

    \I__2190\ : SRMux
    port map (
            O => \N__24282\,
            I => \N__24275\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__24279\,
            I => \N__24272\
        );

    \I__2188\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24268\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__24275\,
            I => \N__24265\
        );

    \I__2186\ : Span4Mux_v
    port map (
            O => \N__24272\,
            I => \N__24262\
        );

    \I__2185\ : InMux
    port map (
            O => \N__24271\,
            I => \N__24259\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__24268\,
            I => \b_delay_counter_15__N_4141_adj_4548\
        );

    \I__2183\ : Odrv12
    port map (
            O => \N__24265\,
            I => \b_delay_counter_15__N_4141_adj_4548\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__24262\,
            I => \b_delay_counter_15__N_4141_adj_4548\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__24259\,
            I => \b_delay_counter_15__N_4141_adj_4548\
        );

    \I__2180\ : InMux
    port map (
            O => \N__24250\,
            I => \N__24247\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__24247\,
            I => \quad_counter1.A_delayed\
        );

    \I__2178\ : InMux
    port map (
            O => \N__24244\,
            I => \N__24240\
        );

    \I__2177\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24237\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24233\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__24237\,
            I => \N__24230\
        );

    \I__2174\ : InMux
    port map (
            O => \N__24236\,
            I => \N__24227\
        );

    \I__2173\ : Span4Mux_h
    port map (
            O => \N__24233\,
            I => \N__24224\
        );

    \I__2172\ : Odrv12
    port map (
            O => \N__24230\,
            I => \B_filtered_adj_4539\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__24227\,
            I => \B_filtered_adj_4539\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__24224\,
            I => \B_filtered_adj_4539\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__24217\,
            I => \count_enable_adj_4544_cascade_\
        );

    \I__2168\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24208\
        );

    \I__2167\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24208\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__24208\,
            I => data_out_frame_10_6
        );

    \I__2165\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24202\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__24202\,
            I => \N__24198\
        );

    \I__2163\ : InMux
    port map (
            O => \N__24201\,
            I => \N__24195\
        );

    \I__2162\ : Span4Mux_h
    port map (
            O => \N__24198\,
            I => \N__24192\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__24195\,
            I => \quad_counter1.b_delay_counter_7\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__24192\,
            I => \quad_counter1.b_delay_counter_7\
        );

    \I__2159\ : InMux
    port map (
            O => \N__24187\,
            I => \quad_counter1.n19509\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__24184\,
            I => \N__24181\
        );

    \I__2157\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24177\
        );

    \I__2156\ : InMux
    port map (
            O => \N__24180\,
            I => \N__24174\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__24177\,
            I => \N__24171\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__24174\,
            I => \quad_counter1.b_delay_counter_8\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__24171\,
            I => \quad_counter1.b_delay_counter_8\
        );

    \I__2152\ : InMux
    port map (
            O => \N__24166\,
            I => \bfn_9_11_0_\
        );

    \I__2151\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24160\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__24160\,
            I => \N__24156\
        );

    \I__2149\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24153\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__24156\,
            I => \N__24150\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__24153\,
            I => \quad_counter1.b_delay_counter_9\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__24150\,
            I => \quad_counter1.b_delay_counter_9\
        );

    \I__2145\ : InMux
    port map (
            O => \N__24145\,
            I => \quad_counter1.n19511\
        );

    \I__2144\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24138\
        );

    \I__2143\ : InMux
    port map (
            O => \N__24141\,
            I => \N__24135\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__24138\,
            I => \N__24132\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__24135\,
            I => \quad_counter1.b_delay_counter_10\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__24132\,
            I => \quad_counter1.b_delay_counter_10\
        );

    \I__2139\ : InMux
    port map (
            O => \N__24127\,
            I => \quad_counter1.n19512\
        );

    \I__2138\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24120\
        );

    \I__2137\ : InMux
    port map (
            O => \N__24123\,
            I => \N__24117\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__24120\,
            I => \N__24114\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__24117\,
            I => \quad_counter1.b_delay_counter_11\
        );

    \I__2134\ : Odrv12
    port map (
            O => \N__24114\,
            I => \quad_counter1.b_delay_counter_11\
        );

    \I__2133\ : InMux
    port map (
            O => \N__24109\,
            I => \quad_counter1.n19513\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__24106\,
            I => \N__24103\
        );

    \I__2131\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24099\
        );

    \I__2130\ : InMux
    port map (
            O => \N__24102\,
            I => \N__24096\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__24099\,
            I => \N__24093\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__24096\,
            I => \quad_counter1.b_delay_counter_12\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__24093\,
            I => \quad_counter1.b_delay_counter_12\
        );

    \I__2126\ : InMux
    port map (
            O => \N__24088\,
            I => \quad_counter1.n19514\
        );

    \I__2125\ : InMux
    port map (
            O => \N__24085\,
            I => \N__24082\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__24082\,
            I => \N__24078\
        );

    \I__2123\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24075\
        );

    \I__2122\ : Span4Mux_h
    port map (
            O => \N__24078\,
            I => \N__24072\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__24075\,
            I => \quad_counter1.b_delay_counter_13\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__24072\,
            I => \quad_counter1.b_delay_counter_13\
        );

    \I__2119\ : InMux
    port map (
            O => \N__24067\,
            I => \quad_counter1.n19515\
        );

    \I__2118\ : InMux
    port map (
            O => \N__24064\,
            I => \N__24060\
        );

    \I__2117\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24057\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__24060\,
            I => \N__24054\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__24057\,
            I => \quad_counter1.b_delay_counter_14\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__24054\,
            I => \quad_counter1.b_delay_counter_14\
        );

    \I__2113\ : InMux
    port map (
            O => \N__24049\,
            I => \quad_counter1.n19516\
        );

    \I__2112\ : InMux
    port map (
            O => \N__24046\,
            I => \N__24043\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__24043\,
            I => \N__24038\
        );

    \I__2110\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24033\
        );

    \I__2109\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24033\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__24038\,
            I => b_delay_counter_0_adj_4541
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__24033\,
            I => b_delay_counter_0_adj_4541
        );

    \I__2106\ : InMux
    port map (
            O => \N__24028\,
            I => \N__24025\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__24025\,
            I => \N__24022\
        );

    \I__2104\ : Odrv12
    port map (
            O => \N__24022\,
            I => n187_adj_4546
        );

    \I__2103\ : InMux
    port map (
            O => \N__24019\,
            I => \bfn_9_10_0_\
        );

    \I__2102\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24013\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__24013\,
            I => \N__24009\
        );

    \I__2100\ : InMux
    port map (
            O => \N__24012\,
            I => \N__24006\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__24009\,
            I => \N__24003\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__24006\,
            I => \quad_counter1.b_delay_counter_1\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__24003\,
            I => \quad_counter1.b_delay_counter_1\
        );

    \I__2096\ : InMux
    port map (
            O => \N__23998\,
            I => \quad_counter1.n19503\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__23995\,
            I => \N__23992\
        );

    \I__2094\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23989\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__23989\,
            I => \N__23985\
        );

    \I__2092\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23982\
        );

    \I__2091\ : Span4Mux_h
    port map (
            O => \N__23985\,
            I => \N__23979\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__23982\,
            I => \quad_counter1.b_delay_counter_2\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__23979\,
            I => \quad_counter1.b_delay_counter_2\
        );

    \I__2088\ : InMux
    port map (
            O => \N__23974\,
            I => \quad_counter1.n19504\
        );

    \I__2087\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23967\
        );

    \I__2086\ : InMux
    port map (
            O => \N__23970\,
            I => \N__23964\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__23967\,
            I => \N__23961\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__23964\,
            I => \quad_counter1.b_delay_counter_3\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__23961\,
            I => \quad_counter1.b_delay_counter_3\
        );

    \I__2082\ : InMux
    port map (
            O => \N__23956\,
            I => \quad_counter1.n19505\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__23953\,
            I => \N__23950\
        );

    \I__2080\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23946\
        );

    \I__2079\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23943\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__23946\,
            I => \N__23940\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__23943\,
            I => \quad_counter1.b_delay_counter_4\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__23940\,
            I => \quad_counter1.b_delay_counter_4\
        );

    \I__2075\ : InMux
    port map (
            O => \N__23935\,
            I => \quad_counter1.n19506\
        );

    \I__2074\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23929\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__23929\,
            I => \N__23925\
        );

    \I__2072\ : InMux
    port map (
            O => \N__23928\,
            I => \N__23922\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__23925\,
            I => \N__23919\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__23922\,
            I => \quad_counter1.b_delay_counter_5\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__23919\,
            I => \quad_counter1.b_delay_counter_5\
        );

    \I__2068\ : InMux
    port map (
            O => \N__23914\,
            I => \quad_counter1.n19507\
        );

    \I__2067\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23908\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__23908\,
            I => \N__23904\
        );

    \I__2065\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23901\
        );

    \I__2064\ : Span4Mux_h
    port map (
            O => \N__23904\,
            I => \N__23898\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__23901\,
            I => \quad_counter1.b_delay_counter_6\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__23898\,
            I => \quad_counter1.b_delay_counter_6\
        );

    \I__2061\ : InMux
    port map (
            O => \N__23893\,
            I => \quad_counter1.n19508\
        );

    \I__2060\ : SRMux
    port map (
            O => \N__23890\,
            I => \N__23887\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__23887\,
            I => \N__23884\
        );

    \I__2058\ : Sp12to4
    port map (
            O => \N__23884\,
            I => \N__23881\
        );

    \I__2057\ : Odrv12
    port map (
            O => \N__23881\,
            I => \c0.n21322\
        );

    \I__2056\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23875\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__23875\,
            I => \N__23872\
        );

    \I__2054\ : Span4Mux_v
    port map (
            O => \N__23872\,
            I => \N__23868\
        );

    \I__2053\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23865\
        );

    \I__2052\ : Sp12to4
    port map (
            O => \N__23868\,
            I => \N__23860\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__23865\,
            I => \N__23860\
        );

    \I__2050\ : Span12Mux_h
    port map (
            O => \N__23860\,
            I => \N__23857\
        );

    \I__2049\ : Odrv12
    port map (
            O => \N__23857\,
            I => rx_i
        );

    \I__2048\ : InMux
    port map (
            O => \N__23854\,
            I => \N__23851\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__23851\,
            I => \quad_counter1.n27\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__23848\,
            I => \quad_counter1.n28_cascade_\
        );

    \I__2045\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23842\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__23842\,
            I => \quad_counter1.n25\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__23839\,
            I => \n9818_cascade_\
        );

    \I__2042\ : InMux
    port map (
            O => \N__23836\,
            I => \c0.n19616\
        );

    \I__2041\ : InMux
    port map (
            O => \N__23833\,
            I => \c0.n19617\
        );

    \I__2040\ : InMux
    port map (
            O => \N__23830\,
            I => \c0.n19618\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__23827\,
            I => \n23768_cascade_\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__23824\,
            I => \n23897_cascade_\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__23821\,
            I => \n10_adj_4532_cascade_\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__23818\,
            I => \quad_counter1.n26_adj_4207_cascade_\
        );

    \I__2035\ : InMux
    port map (
            O => \N__23815\,
            I => \N__23812\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__23812\,
            I => \quad_counter1.n25_adj_4209\
        );

    \I__2033\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23806\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__23806\,
            I => \N__23803\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__23803\,
            I => n12907
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__23800\,
            I => \N__23795\
        );

    \I__2029\ : InMux
    port map (
            O => \N__23799\,
            I => \N__23790\
        );

    \I__2028\ : InMux
    port map (
            O => \N__23798\,
            I => \N__23790\
        );

    \I__2027\ : InMux
    port map (
            O => \N__23795\,
            I => \N__23787\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__23790\,
            I => \N__23784\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__23787\,
            I => \quadB_delayed_adj_4543\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__23784\,
            I => \quadB_delayed_adj_4543\
        );

    \I__2023\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23773\
        );

    \I__2022\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23773\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__23773\,
            I => \N__23768\
        );

    \I__2020\ : InMux
    port map (
            O => \N__23772\,
            I => \N__23763\
        );

    \I__2019\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23763\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__23768\,
            I => \N__23760\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__23763\,
            I => \N__23757\
        );

    \I__2016\ : Sp12to4
    port map (
            O => \N__23760\,
            I => \N__23752\
        );

    \I__2015\ : Sp12to4
    port map (
            O => \N__23757\,
            I => \N__23752\
        );

    \I__2014\ : Span12Mux_v
    port map (
            O => \N__23752\,
            I => \N__23749\
        );

    \I__2013\ : Odrv12
    port map (
            O => \N__23749\,
            I => \PIN_13_c\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__23746\,
            I => \n12907_cascade_\
        );

    \I__2011\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23740\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__23740\,
            I => \quad_counter1.n27_adj_4208\
        );

    \I__2009\ : InMux
    port map (
            O => \N__23737\,
            I => \N__23734\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__23734\,
            I => \quad_counter1.n28_adj_4206\
        );

    \I__2007\ : InMux
    port map (
            O => \N__23731\,
            I => \c0.n19612\
        );

    \I__2006\ : InMux
    port map (
            O => \N__23728\,
            I => \c0.n19613\
        );

    \I__2005\ : InMux
    port map (
            O => \N__23725\,
            I => \c0.n19614\
        );

    \I__2004\ : InMux
    port map (
            O => \N__23722\,
            I => \c0.n19615\
        );

    \I__2003\ : IoInMux
    port map (
            O => \N__23719\,
            I => \N__23716\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__23716\,
            I => \N__23713\
        );

    \I__2001\ : IoSpan4Mux
    port map (
            O => \N__23713\,
            I => \N__23710\
        );

    \I__2000\ : Span4Mux_s3_v
    port map (
            O => \N__23710\,
            I => \N__23707\
        );

    \I__1999\ : Sp12to4
    port map (
            O => \N__23707\,
            I => \N__23704\
        );

    \I__1998\ : Span12Mux_v
    port map (
            O => \N__23704\,
            I => \N__23701\
        );

    \I__1997\ : Span12Mux_v
    port map (
            O => \N__23701\,
            I => \N__23698\
        );

    \I__1996\ : Odrv12
    port map (
            O => \N__23698\,
            I => \CLK_c\
        );

    \I__1995\ : IoInMux
    port map (
            O => \N__23695\,
            I => \N__23692\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__23692\,
            I => tx_enable
        );

    \I__1993\ : IoInMux
    port map (
            O => \N__23689\,
            I => \N__23686\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__23686\,
            I => \GB_BUFFER_PIN_9_c_THRU_CO\
        );

    \I__1991\ : IoInMux
    port map (
            O => \N__23683\,
            I => \N__23680\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__23680\,
            I => \N__23677\
        );

    \I__1989\ : Span12Mux_s2_v
    port map (
            O => \N__23677\,
            I => \N__23674\
        );

    \I__1988\ : Span12Mux_v
    port map (
            O => \N__23674\,
            I => \N__23671\
        );

    \I__1987\ : Odrv12
    port map (
            O => \N__23671\,
            I => \LED_c\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19555\,
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19563\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19571\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19579\,
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19587\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19595\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19603\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19611\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19510\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter1.n19525\,
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19480\,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_10_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n19495\,
            carryinitout => \bfn_10_25_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.tx.n19547\,
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_20_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_24_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_19_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_1_0_\
        );

    \IN_MUX_bfv_19_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19442_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_2_0_\
        );

    \IN_MUX_bfv_19_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19443_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_3_0_\
        );

    \IN_MUX_bfv_19_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19444_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_4_0_\
        );

    \IN_MUX_bfv_19_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19445_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_5_0_\
        );

    \IN_MUX_bfv_19_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19446_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_6_0_\
        );

    \IN_MUX_bfv_19_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19447_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_7_0_\
        );

    \IN_MUX_bfv_19_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19448_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_8_0_\
        );

    \IN_MUX_bfv_19_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19449_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_9_0_\
        );

    \IN_MUX_bfv_19_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19450_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_10_0_\
        );

    \IN_MUX_bfv_19_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19451_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_11_0_\
        );

    \IN_MUX_bfv_19_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19452_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_12_0_\
        );

    \IN_MUX_bfv_19_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19453_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_13_0_\
        );

    \IN_MUX_bfv_19_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19454_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_14_0_\
        );

    \IN_MUX_bfv_19_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19455_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_15_0_\
        );

    \IN_MUX_bfv_19_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19456_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_16_0_\
        );

    \IN_MUX_bfv_19_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19457_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_17_0_\
        );

    \IN_MUX_bfv_19_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19458_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_18_0_\
        );

    \IN_MUX_bfv_19_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19459_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_19_0_\
        );

    \IN_MUX_bfv_19_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19460_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_20_0_\
        );

    \IN_MUX_bfv_19_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19461_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_21_0_\
        );

    \IN_MUX_bfv_19_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19462_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_22_0_\
        );

    \IN_MUX_bfv_19_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19463_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_23_0_\
        );

    \IN_MUX_bfv_19_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19464_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_24_0_\
        );

    \IN_MUX_bfv_19_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19465_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_25_0_\
        );

    \IN_MUX_bfv_19_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19466_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_26_0_\
        );

    \IN_MUX_bfv_19_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19467_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_27_0_\
        );

    \IN_MUX_bfv_19_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19468_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_28_0_\
        );

    \IN_MUX_bfv_19_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19469_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_29_0_\
        );

    \IN_MUX_bfv_19_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19470_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_30_0_\
        );

    \IN_MUX_bfv_19_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19471_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_31_0_\
        );

    \IN_MUX_bfv_19_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \c0.n19472_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_19_32_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \c0.tx.i8_1_lut_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26517\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => tx_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_PIN_9_c_THRU_LUT4_0_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66880\,
            lcout => \GB_BUFFER_PIN_9_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rx_i_I_0_1_lut_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23871\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.quadB_delayed_62_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27574\,
            lcout => \quadB_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i23_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37641\,
            in2 => \_gnd_net_\,
            in3 => \N__52868\,
            lcout => \c0.FRAME_MATCHER_state_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66867\,
            ce => 'H',
            sr => \N__23890\
        );

    \c0.FRAME_MATCHER_state_i26_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37318\,
            in2 => \_gnd_net_\,
            in3 => \N__52891\,
            lcout => \c0.FRAME_MATCHER_state_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66870\,
            ce => 'H',
            sr => \N__29245\
        );

    \quad_counter1.quadA_delayed_61_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25946\,
            lcout => \quadA_delayed_adj_4542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66695\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.B_65_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101000"
        )
    port map (
            in0 => \N__24236\,
            in1 => \N__23771\,
            in2 => \N__23800\,
            in3 => \N__23809\,
            lcout => \B_filtered_adj_4539\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66723\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.quadB_delayed_62_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23772\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quadB_delayed_adj_4543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66723\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i9_4_lut_adj_1169_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__24163\,
            in1 => \N__23971\,
            in2 => \N__23953\,
            in3 => \N__24041\,
            lcout => \quad_counter1.n25_adj_4209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.b_delay_counter__i0_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__24028\,
            in1 => \N__24042\,
            in2 => \N__24316\,
            in3 => \N__24278\,
            lcout => b_delay_counter_0_adj_4541,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.quadB_I_0_79_2_lut_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23779\,
            lcout => \b_delay_counter_15__N_4141_adj_4548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i10_4_lut_adj_1167_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24142\,
            in1 => \N__24124\,
            in2 => \N__24184\,
            in3 => \N__23911\,
            lcout => OPEN,
            ltout => \quad_counter1.n26_adj_4207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i15_4_lut_adj_1170_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23737\,
            in1 => \N__23743\,
            in2 => \N__23818\,
            in3 => \N__23815\,
            lcout => n12907,
            ltout => \n12907_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_1918_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010000"
        )
    port map (
            in0 => \N__23799\,
            in1 => \N__23778\,
            in2 => \N__23746\,
            in3 => \N__24271\,
            lcout => n14377,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i11_4_lut_adj_1168_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24064\,
            in1 => \N__24205\,
            in2 => \N__24106\,
            in3 => \N__24331\,
            lcout => \quad_counter1.n27_adj_4208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i12_4_lut_adj_1166_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__24016\,
            in1 => \N__24085\,
            in2 => \N__23995\,
            in3 => \N__23932\,
            lcout => \quad_counter1.n28_adj_4206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1411__i0_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39189\,
            in2 => \N__39720\,
            in3 => \_gnd_net_\,
            lcout => \c0.byte_transmit_counter_0\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \c0.n19612\,
            clk => \N__66822\,
            ce => \N__39220\,
            sr => \N__39202\
        );

    \c0.byte_transmit_counter_1411__i1_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36742\,
            in2 => \_gnd_net_\,
            in3 => \N__23731\,
            lcout => \c0.byte_transmit_counter_1\,
            ltout => OPEN,
            carryin => \c0.n19612\,
            carryout => \c0.n19613\,
            clk => \N__66822\,
            ce => \N__39220\,
            sr => \N__39202\
        );

    \c0.byte_transmit_counter_1411__i2_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33863\,
            in2 => \_gnd_net_\,
            in3 => \N__23728\,
            lcout => \c0.byte_transmit_counter_2\,
            ltout => OPEN,
            carryin => \c0.n19613\,
            carryout => \c0.n19614\,
            clk => \N__66822\,
            ce => \N__39220\,
            sr => \N__39202\
        );

    \c0.byte_transmit_counter_1411__i3_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25626\,
            in2 => \_gnd_net_\,
            in3 => \N__23725\,
            lcout => byte_transmit_counter_3,
            ltout => OPEN,
            carryin => \c0.n19614\,
            carryout => \c0.n19615\,
            clk => \N__66822\,
            ce => \N__39220\,
            sr => \N__39202\
        );

    \c0.byte_transmit_counter_1411__i4_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26742\,
            in2 => \_gnd_net_\,
            in3 => \N__23722\,
            lcout => byte_transmit_counter_4,
            ltout => OPEN,
            carryin => \c0.n19615\,
            carryout => \c0.n19616\,
            clk => \N__66822\,
            ce => \N__39220\,
            sr => \N__39202\
        );

    \c0.byte_transmit_counter_1411__i5_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27308\,
            in2 => \_gnd_net_\,
            in3 => \N__23836\,
            lcout => byte_transmit_counter_5,
            ltout => OPEN,
            carryin => \c0.n19616\,
            carryout => \c0.n19617\,
            clk => \N__66822\,
            ce => \N__39220\,
            sr => \N__39202\
        );

    \c0.byte_transmit_counter_1411__i6_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26931\,
            in2 => \_gnd_net_\,
            in3 => \N__23833\,
            lcout => \c0.byte_transmit_counter_6\,
            ltout => OPEN,
            carryin => \c0.n19617\,
            carryout => \c0.n19618\,
            clk => \N__66822\,
            ce => \N__39220\,
            sr => \N__39202\
        );

    \c0.byte_transmit_counter_1411__i7_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26910\,
            in2 => \_gnd_net_\,
            in3 => \N__23830\,
            lcout => \c0.byte_transmit_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66822\,
            ce => \N__39220\,
            sr => \N__39202\
        );

    \c0.i2_3_lut_adj_1673_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__36741\,
            in1 => \N__33854\,
            in2 => \_gnd_net_\,
            in3 => \N__25589\,
            lcout => n23768,
            ltout => \n23768_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20202_4_lut_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__29443\,
            in1 => \N__24442\,
            in2 => \N__23827\,
            in3 => \N__26743\,
            lcout => OPEN,
            ltout => \n23897_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_1913_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__26744\,
            in1 => \N__24523\,
            in2 => \N__23824\,
            in3 => \N__25590\,
            lcout => OPEN,
            ltout => \n10_adj_4532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i5_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__29154\,
            in1 => \N__25521\,
            in2 => \N__23821\,
            in3 => \N__27309\,
            lcout => \r_Tx_Data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66834\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i2_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__24621\,
            in1 => \N__27322\,
            in2 => \N__24577\,
            in3 => \N__29144\,
            lcout => \r_Tx_Data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i6_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__29145\,
            in1 => \N__24639\,
            in2 => \N__27334\,
            in3 => \N__24454\,
            lcout => \r_Tx_Data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1517_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37640\,
            in2 => \_gnd_net_\,
            in3 => \N__40657\,
            lcout => \c0.n21322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Data_R_49_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.rx.r_Rx_Data_R\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_4_i26_3_lut_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39838\,
            in1 => \N__26098\,
            in2 => \_gnd_net_\,
            in3 => \N__29254\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__1__5428_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__34710\,
            in1 => \N__49179\,
            in2 => \N__32311\,
            in3 => \N__49040\,
            lcout => data_out_frame_12_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i9_4_lut_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__24699\,
            in1 => \N__24840\,
            in2 => \N__24718\,
            in3 => \N__24889\,
            lcout => \quad_counter1.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i11_4_lut_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24819\,
            in1 => \N__24682\,
            in2 => \N__24859\,
            in3 => \N__24801\,
            lcout => \quad_counter1.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i12_4_lut_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__24732\,
            in1 => \N__24664\,
            in2 => \N__24751\,
            in3 => \N__24768\,
            lcout => OPEN,
            ltout => \quad_counter1.n28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i15_4_lut_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26032\,
            in1 => \N__23854\,
            in2 => \N__23848\,
            in3 => \N__23845\,
            lcout => n9818,
            ltout => \n9818_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.A_63_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001000"
        )
    port map (
            in0 => \N__25959\,
            in1 => \N__25993\,
            in2 => \N__23839\,
            in3 => \N__24938\,
            lcout => \A_filtered_adj_4538\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i1073_1_lut_2_lut_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24911\,
            in2 => \_gnd_net_\,
            in3 => \N__24937\,
            lcout => \quad_counter1.n2140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.B_delayed_68_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24243\,
            lcout => \quad_counter1.B_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_86_2_lut_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24046\,
            in2 => \_gnd_net_\,
            in3 => \N__24019\,
            lcout => n187_adj_4546,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \quad_counter1.n19503\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.b_delay_counter__i1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24012\,
            in2 => \_gnd_net_\,
            in3 => \N__23998\,
            lcout => \quad_counter1.b_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter1.n19503\,
            carryout => \quad_counter1.n19504\,
            clk => \N__66709\,
            ce => \N__24311\,
            sr => \N__24283\
        );

    \quad_counter1.b_delay_counter__i2_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23988\,
            in2 => \_gnd_net_\,
            in3 => \N__23974\,
            lcout => \quad_counter1.b_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter1.n19504\,
            carryout => \quad_counter1.n19505\,
            clk => \N__66709\,
            ce => \N__24311\,
            sr => \N__24283\
        );

    \quad_counter1.b_delay_counter__i3_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23970\,
            in2 => \_gnd_net_\,
            in3 => \N__23956\,
            lcout => \quad_counter1.b_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter1.n19505\,
            carryout => \quad_counter1.n19506\,
            clk => \N__66709\,
            ce => \N__24311\,
            sr => \N__24283\
        );

    \quad_counter1.b_delay_counter__i4_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23949\,
            in2 => \_gnd_net_\,
            in3 => \N__23935\,
            lcout => \quad_counter1.b_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter1.n19506\,
            carryout => \quad_counter1.n19507\,
            clk => \N__66709\,
            ce => \N__24311\,
            sr => \N__24283\
        );

    \quad_counter1.b_delay_counter__i5_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23928\,
            in2 => \_gnd_net_\,
            in3 => \N__23914\,
            lcout => \quad_counter1.b_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter1.n19507\,
            carryout => \quad_counter1.n19508\,
            clk => \N__66709\,
            ce => \N__24311\,
            sr => \N__24283\
        );

    \quad_counter1.b_delay_counter__i6_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23907\,
            in2 => \_gnd_net_\,
            in3 => \N__23893\,
            lcout => \quad_counter1.b_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter1.n19508\,
            carryout => \quad_counter1.n19509\,
            clk => \N__66709\,
            ce => \N__24311\,
            sr => \N__24283\
        );

    \quad_counter1.b_delay_counter__i7_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24201\,
            in2 => \_gnd_net_\,
            in3 => \N__24187\,
            lcout => \quad_counter1.b_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter1.n19509\,
            carryout => \quad_counter1.n19510\,
            clk => \N__66709\,
            ce => \N__24311\,
            sr => \N__24283\
        );

    \quad_counter1.b_delay_counter__i8_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24180\,
            in2 => \_gnd_net_\,
            in3 => \N__24166\,
            lcout => \quad_counter1.b_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \quad_counter1.n19511\,
            clk => \N__66724\,
            ce => \N__24315\,
            sr => \N__24282\
        );

    \quad_counter1.b_delay_counter__i9_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24159\,
            in2 => \_gnd_net_\,
            in3 => \N__24145\,
            lcout => \quad_counter1.b_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter1.n19511\,
            carryout => \quad_counter1.n19512\,
            clk => \N__66724\,
            ce => \N__24315\,
            sr => \N__24282\
        );

    \quad_counter1.b_delay_counter__i10_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24141\,
            in2 => \_gnd_net_\,
            in3 => \N__24127\,
            lcout => \quad_counter1.b_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter1.n19512\,
            carryout => \quad_counter1.n19513\,
            clk => \N__66724\,
            ce => \N__24315\,
            sr => \N__24282\
        );

    \quad_counter1.b_delay_counter__i11_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24123\,
            in2 => \_gnd_net_\,
            in3 => \N__24109\,
            lcout => \quad_counter1.b_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter1.n19513\,
            carryout => \quad_counter1.n19514\,
            clk => \N__66724\,
            ce => \N__24315\,
            sr => \N__24282\
        );

    \quad_counter1.b_delay_counter__i12_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24102\,
            in2 => \_gnd_net_\,
            in3 => \N__24088\,
            lcout => \quad_counter1.b_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter1.n19514\,
            carryout => \quad_counter1.n19515\,
            clk => \N__66724\,
            ce => \N__24315\,
            sr => \N__24282\
        );

    \quad_counter1.b_delay_counter__i13_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24081\,
            in2 => \_gnd_net_\,
            in3 => \N__24067\,
            lcout => \quad_counter1.b_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter1.n19515\,
            carryout => \quad_counter1.n19516\,
            clk => \N__66724\,
            ce => \N__24315\,
            sr => \N__24282\
        );

    \quad_counter1.b_delay_counter__i14_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24063\,
            in2 => \_gnd_net_\,
            in3 => \N__24049\,
            lcout => \quad_counter1.b_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter1.n19516\,
            carryout => \quad_counter1.n19517\,
            clk => \N__66724\,
            ce => \N__24315\,
            sr => \N__24282\
        );

    \quad_counter1.b_delay_counter__i15_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24330\,
            in2 => \_gnd_net_\,
            in3 => \N__24334\,
            lcout => \quad_counter1.b_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66724\,
            ce => \N__24315\,
            sr => \N__24282\
        );

    \quad_counter1.A_delayed_67_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quad_counter1.A_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20187_4_lut_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__26446\,
            in1 => \N__36902\,
            in2 => \N__34654\,
            in3 => \N__33976\,
            lcout => \c0.n23882\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__0__5421_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__26212\,
            in1 => \N__49565\,
            in2 => \N__25027\,
            in3 => \N__49020\,
            lcout => data_out_frame_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1406_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25021\,
            in2 => \_gnd_net_\,
            in3 => \N__26320\,
            lcout => \c0.n6_adj_4308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.i3_4_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__24919\,
            in1 => \N__24250\,
            in2 => \N__24955\,
            in3 => \N__24244\,
            lcout => count_enable_adj_4544,
            ltout => \count_enable_adj_4544_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24994\,
            in2 => \N__24217\,
            in3 => \N__25025\,
            lcout => encoder1_position_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i6_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25060\,
            in1 => \N__38356\,
            in2 => \_gnd_net_\,
            in3 => \N__34957\,
            lcout => encoder1_position_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__6__5439_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49273\,
            in1 => \N__49022\,
            in2 => \N__35530\,
            in3 => \N__24214\,
            lcout => data_out_frame_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_20461_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__24213\,
            in1 => \N__36834\,
            in2 => \N__24790\,
            in3 => \N__39781\,
            lcout => \c0.n24153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__5__5464_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49274\,
            in1 => \N__49023\,
            in2 => \N__36004\,
            in3 => \N__26571\,
            lcout => data_out_frame_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20420_4_lut_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__26875\,
            in1 => \N__24340\,
            in2 => \N__26797\,
            in3 => \N__24376\,
            lcout => OPEN,
            ltout => \n24118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i4_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__29155\,
            in1 => \N__25503\,
            in2 => \N__24367\,
            in3 => \N__27338\,
            lcout => \r_Tx_Data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20414_4_lut_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__26266\,
            in1 => \N__33969\,
            in2 => \N__36910\,
            in3 => \N__24385\,
            lcout => n24112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20399_2_lut_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__39758\,
            in1 => \N__30115\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n23950_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_1__bdd_4_lut_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__26248\,
            in1 => \N__36906\,
            in2 => \N__24364\,
            in3 => \N__33970\,
            lcout => OPEN,
            ltout => \c0.n24147_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n24147_bdd_4_lut_4_lut_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100100"
        )
    port map (
            in0 => \N__39759\,
            in1 => \N__25429\,
            in2 => \N__24361\,
            in3 => \N__33938\,
            lcout => n24150,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20400_4_lut_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__24358\,
            in1 => \N__36907\,
            in2 => \N__30214\,
            in3 => \N__33971\,
            lcout => OPEN,
            ltout => \n24097_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20419_3_lut_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24349\,
            in2 => \N__24343\,
            in3 => \N__25638\,
            lcout => n24117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__3__5442_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49379\,
            in1 => \N__49013\,
            in2 => \N__30175\,
            in3 => \N__24402\,
            lcout => data_out_frame_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66766\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i15_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38411\,
            in1 => \N__25120\,
            in2 => \_gnd_net_\,
            in3 => \N__26311\,
            lcout => encoder1_position_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20154_4_lut_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__34753\,
            in1 => \N__24421\,
            in2 => \N__26874\,
            in3 => \N__26789\,
            lcout => OPEN,
            ltout => \n23849_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_1915_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__26790\,
            in1 => \N__24412\,
            in2 => \N__24406\,
            in3 => \N__25634\,
            lcout => n10_adj_4536,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_6_i11_3_lut_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29887\,
            in1 => \N__28543\,
            in2 => \_gnd_net_\,
            in3 => \N__39773\,
            lcout => \c0.n11_adj_4355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i28_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36495\,
            in1 => \N__25336\,
            in2 => \_gnd_net_\,
            in3 => \N__38412\,
            lcout => encoder1_position_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20151_4_lut_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__26865\,
            in1 => \N__24427\,
            in2 => \N__26796\,
            in3 => \N__29311\,
            lcout => n23846,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_20476_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__24403\,
            in1 => \N__36862\,
            in2 => \N__28525\,
            in3 => \N__39772\,
            lcout => \c0.n24171\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_20466_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__39771\,
            in1 => \N__28708\,
            in2 => \N__36900\,
            in3 => \N__28740\,
            lcout => OPEN,
            ltout => \c0.n24159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n24159_bdd_4_lut_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__26542\,
            in1 => \N__36863\,
            in2 => \N__24388\,
            in3 => \N__28723\,
            lcout => \c0.n24162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20416_4_lut_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__24469\,
            in1 => \N__33942\,
            in2 => \N__36901\,
            in3 => \N__28555\,
            lcout => OPEN,
            ltout => \n24114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_1916_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__26788\,
            in1 => \N__24463\,
            in2 => \N__24457\,
            in3 => \N__25635\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20200_4_lut_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__33889\,
            in1 => \N__36761\,
            in2 => \N__26557\,
            in3 => \N__24514\,
            lcout => \c0.n23895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_5_i11_3_lut_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25410\,
            in1 => \N__38020\,
            in2 => \_gnd_net_\,
            in3 => \N__39701\,
            lcout => \c0.n11_adj_4348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i31_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25438\,
            in1 => \N__38458\,
            in2 => \_gnd_net_\,
            in3 => \N__28771\,
            lcout => encoder1_position_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i18_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25105\,
            in1 => \N__38457\,
            in2 => \_gnd_net_\,
            in3 => \N__29032\,
            lcout => encoder1_position_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20355_3_lut_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__26677\,
            in1 => \N__33886\,
            in2 => \_gnd_net_\,
            in3 => \N__39700\,
            lcout => OPEN,
            ltout => \c0.n24051_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20149_4_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33888\,
            in1 => \N__39514\,
            in2 => \N__24430\,
            in3 => \N__36760\,
            lcout => \c0.n23844\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20152_4_lut_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__36759\,
            in1 => \N__33887\,
            in2 => \N__33790\,
            in3 => \N__24508\,
            lcout => \c0.n23847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20404_4_lut_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__36848\,
            in1 => \N__27079\,
            in2 => \N__24532\,
            in3 => \N__33948\,
            lcout => n24102,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_0__3__5522_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__24490\,
            in1 => \N__37193\,
            in2 => \_gnd_net_\,
            in3 => \N__40170\,
            lcout => data_out_frame_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20351_4_lut_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000100000000"
        )
    port map (
            in0 => \N__33946\,
            in1 => \N__36847\,
            in2 => \N__27181\,
            in3 => \N__39775\,
            lcout => \c0.n24047\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i6_4_lut_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001000100"
        )
    port map (
            in0 => \N__39776\,
            in1 => \N__24478\,
            in2 => \N__26893\,
            in3 => \N__33947\,
            lcout => \c0.n6_adj_4521\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_7_i5_3_lut_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33436\,
            in1 => \N__24498\,
            in2 => \_gnd_net_\,
            in3 => \N__39774\,
            lcout => \c0.n5_adj_4358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__7__5470_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__48844\,
            in1 => \N__49447\,
            in2 => \N__24502\,
            in3 => \N__41646\,
            lcout => data_out_frame_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__3__5418_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49446\,
            in1 => \N__48845\,
            in2 => \N__28357\,
            in3 => \N__26658\,
            lcout => data_out_frame_13_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66810\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20385_2_lut_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24489\,
            in2 => \_gnd_net_\,
            in3 => \N__36870\,
            lcout => \c0.n24007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20389_2_lut_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__36871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24600\,
            lcout => \c0.n24011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20161_4_lut_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__24538\,
            in1 => \N__36872\,
            in2 => \N__27196\,
            in3 => \N__33964\,
            lcout => \c0.n23856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_0__2__5523_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__24601\,
            in1 => \N__37204\,
            in2 => \_gnd_net_\,
            in3 => \N__40169\,
            lcout => data_out_frame_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20164_4_lut_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__24589\,
            in1 => \N__36873\,
            in2 => \N__24565\,
            in3 => \N__33965\,
            lcout => OPEN,
            ltout => \c0.n23859_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20166_4_lut_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26866\,
            in1 => \N__25858\,
            in2 => \N__24583\,
            in3 => \N__26791\,
            lcout => OPEN,
            ltout => \n23861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_1911_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__26792\,
            in1 => \N__25468\,
            in2 => \N__24580\,
            in3 => \N__25636\,
            lcout => n10_adj_4534,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i5_3_lut_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26371\,
            in1 => \N__24552\,
            in2 => \_gnd_net_\,
            in3 => \N__39779\,
            lcout => \c0.n5_adj_4522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__2__5475_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__49548\,
            in1 => \N__49021\,
            in2 => \N__24556\,
            in3 => \N__40063\,
            lcout => data_out_frame_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20362_4_lut_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010001010"
        )
    port map (
            in0 => \N__39780\,
            in1 => \N__28984\,
            in2 => \N__33975\,
            in3 => \N__36882\,
            lcout => \c0.n24059\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i6_4_lut_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100100010"
        )
    port map (
            in0 => \N__24544\,
            in1 => \N__33959\,
            in2 => \N__27229\,
            in3 => \N__39778\,
            lcout => \c0.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Bit_Index_2__bdd_4_lut_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__24643\,
            in1 => \N__24625\,
            in2 => \N__26989\,
            in3 => \N__27036\,
            lcout => n24195,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i0_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__25769\,
            in1 => \N__25796\,
            in2 => \N__27607\,
            in3 => \N__25693\,
            lcout => b_delay_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.quadA_delayed_61_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27824\,
            lcout => \quadA_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.quadB_I_0_79_2_lut_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27579\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27530\,
            lcout => \b_delay_counter_15__N_4141\,
            ltout => \b_delay_counter_15__N_4141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_1917_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110000"
        )
    port map (
            in0 => \N__27531\,
            in1 => \N__27578\,
            in2 => \N__24607\,
            in3 => \N__27376\,
            lcout => n14198,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i4_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37789\,
            in2 => \_gnd_net_\,
            in3 => \N__52890\,
            lcout => \c0.FRAME_MATCHER_state_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66864\,
            ce => 'H',
            sr => \N__34210\
        );

    \quad_counter0.quadA_I_0_73_2_lut_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27825\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27789\,
            lcout => \a_delay_counter_15__N_4124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1708_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28338\,
            in1 => \N__29710\,
            in2 => \_gnd_net_\,
            in3 => \N__53368\,
            lcout => \c0.n13360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1803_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29425\,
            in1 => \N__32592\,
            in2 => \N__32566\,
            in3 => \N__31636\,
            lcout => \c0.n24_adj_4502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_85_2_lut_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24887\,
            in2 => \_gnd_net_\,
            in3 => \N__24604\,
            lcout => n39_adj_4545,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \quad_counter1.n19518\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.a_delay_counter__i1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24769\,
            in2 => \_gnd_net_\,
            in3 => \N__24754\,
            lcout => \quad_counter1.a_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter1.n19518\,
            carryout => \quad_counter1.n19519\,
            clk => \N__66672\,
            ce => \N__25906\,
            sr => \N__26020\
        );

    \quad_counter1.a_delay_counter__i2_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24750\,
            in2 => \_gnd_net_\,
            in3 => \N__24736\,
            lcout => \quad_counter1.a_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter1.n19519\,
            carryout => \quad_counter1.n19520\,
            clk => \N__66672\,
            ce => \N__25906\,
            sr => \N__26020\
        );

    \quad_counter1.a_delay_counter__i3_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24733\,
            in2 => \_gnd_net_\,
            in3 => \N__24721\,
            lcout => \quad_counter1.a_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter1.n19520\,
            carryout => \quad_counter1.n19521\,
            clk => \N__66672\,
            ce => \N__25906\,
            sr => \N__26020\
        );

    \quad_counter1.a_delay_counter__i4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24717\,
            in2 => \_gnd_net_\,
            in3 => \N__24703\,
            lcout => \quad_counter1.a_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter1.n19521\,
            carryout => \quad_counter1.n19522\,
            clk => \N__66672\,
            ce => \N__25906\,
            sr => \N__26020\
        );

    \quad_counter1.a_delay_counter__i5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24700\,
            in2 => \_gnd_net_\,
            in3 => \N__24688\,
            lcout => \quad_counter1.a_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter1.n19522\,
            carryout => \quad_counter1.n19523\,
            clk => \N__66672\,
            ce => \N__25906\,
            sr => \N__26020\
        );

    \quad_counter1.a_delay_counter__i6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26044\,
            in2 => \_gnd_net_\,
            in3 => \N__24685\,
            lcout => \quad_counter1.a_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter1.n19523\,
            carryout => \quad_counter1.n19524\,
            clk => \N__66672\,
            ce => \N__25906\,
            sr => \N__26020\
        );

    \quad_counter1.a_delay_counter__i7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24681\,
            in2 => \_gnd_net_\,
            in3 => \N__24667\,
            lcout => \quad_counter1.a_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter1.n19524\,
            carryout => \quad_counter1.n19525\,
            clk => \N__66672\,
            ce => \N__25906\,
            sr => \N__26020\
        );

    \quad_counter1.a_delay_counter__i8_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24663\,
            in2 => \_gnd_net_\,
            in3 => \N__24649\,
            lcout => \quad_counter1.a_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \quad_counter1.n19526\,
            clk => \N__66683\,
            ce => \N__25905\,
            sr => \N__26016\
        );

    \quad_counter1.a_delay_counter__i9_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26058\,
            in2 => \_gnd_net_\,
            in3 => \N__24646\,
            lcout => \quad_counter1.a_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter1.n19526\,
            carryout => \quad_counter1.n19527\,
            clk => \N__66683\,
            ce => \N__25905\,
            sr => \N__26016\
        );

    \quad_counter1.a_delay_counter__i10_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24858\,
            in2 => \_gnd_net_\,
            in3 => \N__24844\,
            lcout => \quad_counter1.a_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter1.n19527\,
            carryout => \quad_counter1.n19528\,
            clk => \N__66683\,
            ce => \N__25905\,
            sr => \N__26016\
        );

    \quad_counter1.a_delay_counter__i11_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24841\,
            in2 => \_gnd_net_\,
            in3 => \N__24829\,
            lcout => \quad_counter1.a_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter1.n19528\,
            carryout => \quad_counter1.n19529\,
            clk => \N__66683\,
            ce => \N__25905\,
            sr => \N__26016\
        );

    \quad_counter1.a_delay_counter__i12_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26085\,
            in2 => \_gnd_net_\,
            in3 => \N__24826\,
            lcout => \quad_counter1.a_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter1.n19529\,
            carryout => \quad_counter1.n19530\,
            clk => \N__66683\,
            ce => \N__25905\,
            sr => \N__26016\
        );

    \quad_counter1.a_delay_counter__i13_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26071\,
            in2 => \_gnd_net_\,
            in3 => \N__24823\,
            lcout => \quad_counter1.a_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter1.n19530\,
            carryout => \quad_counter1.n19531\,
            clk => \N__66683\,
            ce => \N__25905\,
            sr => \N__26016\
        );

    \quad_counter1.a_delay_counter__i14_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24820\,
            in2 => \_gnd_net_\,
            in3 => \N__24808\,
            lcout => \quad_counter1.a_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter1.n19531\,
            carryout => \quad_counter1.n19532\,
            clk => \N__66683\,
            ce => \N__25905\,
            sr => \N__26016\
        );

    \quad_counter1.a_delay_counter__i15_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24802\,
            in2 => \_gnd_net_\,
            in3 => \N__24805\,
            lcout => \quad_counter1.a_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66683\,
            ce => \N__25905\,
            sr => \N__26016\
        );

    \c0.i3_4_lut_adj_1403_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35390\,
            in1 => \N__33085\,
            in2 => \N__28219\,
            in3 => \N__28426\,
            lcout => \c0.n10434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__6__5431_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__49017\,
            in1 => \N__49358\,
            in2 => \N__24789\,
            in3 => \N__28481\,
            lcout => data_out_frame_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i3_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24970\,
            in1 => \_gnd_net_\,
            in2 => \N__38410\,
            in3 => \N__28325\,
            lcout => encoder1_position_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__4__5433_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49357\,
            in1 => \N__49018\,
            in2 => \N__38941\,
            in3 => \N__26460\,
            lcout => data_out_frame_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.A_filtered_I_0_2_lut_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24954\,
            in2 => \_gnd_net_\,
            in3 => \N__24918\,
            lcout => \quad_counter1.count_direction\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.a_delay_counter__i0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__26004\,
            in1 => \N__24898\,
            in2 => \N__24888\,
            in3 => \N__25904\,
            lcout => a_delay_counter_0_adj_4540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i5_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38377\,
            in1 => \N__25072\,
            in2 => \_gnd_net_\,
            in3 => \N__32700\,
            lcout => encoder1_position_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1628_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31190\,
            in1 => \N__34348\,
            in2 => \N__32448\,
            in3 => \N__32552\,
            lcout => \c0.n20257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i14_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29640\,
            in1 => \N__38357\,
            in2 => \_gnd_net_\,
            in3 => \N__25132\,
            lcout => encoder1_position_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i2_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__38360\,
            in1 => \_gnd_net_\,
            in2 => \N__35042\,
            in3 => \N__24982\,
            lcout => encoder1_position_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i26_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35644\,
            in1 => \N__25351\,
            in2 => \_gnd_net_\,
            in3 => \N__38359\,
            lcout => encoder1_position_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1405_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36459\,
            in2 => \_gnd_net_\,
            in3 => \N__29639\,
            lcout => \c0.n22116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1807_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32784\,
            in2 => \_gnd_net_\,
            in3 => \N__35031\,
            lcout => OPEN,
            ltout => \c0.n22048_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1810_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31813\,
            in1 => \N__32498\,
            in2 => \N__25030\,
            in3 => \N__28321\,
            lcout => \c0.n20819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i22_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28470\,
            in1 => \N__25084\,
            in2 => \_gnd_net_\,
            in3 => \N__38358\,
            lcout => encoder1_position_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25179\,
            in2 => \N__25308\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \quad_counter1.n19548\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_2_lut_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25026\,
            in2 => \N__25006\,
            in3 => \N__24988\,
            lcout => n2205,
            ltout => OPEN,
            carryin => \quad_counter1.n19548\,
            carryout => \quad_counter1.n19549\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_3_lut_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32785\,
            in2 => \N__25309\,
            in3 => \N__24985\,
            lcout => n2204,
            ltout => OPEN,
            carryin => \quad_counter1.n19549\,
            carryout => \quad_counter1.n19550\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_4_lut_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35035\,
            in2 => \N__25250\,
            in3 => \N__24973\,
            lcout => n2203,
            ltout => OPEN,
            carryin => \quad_counter1.n19550\,
            carryout => \quad_counter1.n19551\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_5_lut_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28334\,
            in2 => \N__25310\,
            in3 => \N__24961\,
            lcout => n2202,
            ltout => OPEN,
            carryin => \quad_counter1.n19551\,
            carryout => \quad_counter1.n19552\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_6_lut_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35139\,
            in2 => \N__25251\,
            in3 => \N__24958\,
            lcout => n2201,
            ltout => OPEN,
            carryin => \quad_counter1.n19552\,
            carryout => \quad_counter1.n19553\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_7_lut_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25186\,
            in2 => \N__32734\,
            in3 => \N__25063\,
            lcout => n2200,
            ltout => OPEN,
            carryin => \quad_counter1.n19553\,
            carryout => \quad_counter1.n19554\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_8_lut_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25261\,
            in2 => \N__34966\,
            in3 => \N__25054\,
            lcout => n2199,
            ltout => OPEN,
            carryin => \quad_counter1.n19554\,
            carryout => \quad_counter1.n19555\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_9_lut_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25262\,
            in2 => \N__34929\,
            in3 => \N__25051\,
            lcout => n2198,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \quad_counter1.n19556\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_10_lut_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35381\,
            in2 => \N__25311\,
            in3 => \N__25048\,
            lcout => n2197,
            ltout => OPEN,
            carryin => \quad_counter1.n19556\,
            carryout => \quad_counter1.n19557\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_11_lut_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25266\,
            in2 => \N__32310\,
            in3 => \N__25045\,
            lcout => n2196,
            ltout => OPEN,
            carryin => \quad_counter1.n19557\,
            carryout => \quad_counter1.n19558\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_12_lut_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35220\,
            in2 => \N__25312\,
            in3 => \N__25042\,
            lcout => n2195,
            ltout => OPEN,
            carryin => \quad_counter1.n19558\,
            carryout => \quad_counter1.n19559\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_13_lut_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25270\,
            in2 => \N__32980\,
            in3 => \N__25039\,
            lcout => n2194,
            ltout => OPEN,
            carryin => \quad_counter1.n19559\,
            carryout => \quad_counter1.n19560\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_14_lut_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34635\,
            in2 => \N__25313\,
            in3 => \N__25036\,
            lcout => n2193,
            ltout => OPEN,
            carryin => \quad_counter1.n19560\,
            carryout => \quad_counter1.n19561\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_15_lut_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25274\,
            in2 => \N__38070\,
            in3 => \N__25033\,
            lcout => n2192,
            ltout => OPEN,
            carryin => \quad_counter1.n19561\,
            carryout => \quad_counter1.n19562\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_16_lut_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29655\,
            in2 => \N__25314\,
            in3 => \N__25123\,
            lcout => n2191,
            ltout => OPEN,
            carryin => \quad_counter1.n19562\,
            carryout => \quad_counter1.n19563\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_17_lut_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26310\,
            in2 => \N__25315\,
            in3 => \N__25114\,
            lcout => n2190,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \quad_counter1.n19564\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_18_lut_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25281\,
            in2 => \N__26427\,
            in3 => \N__25111\,
            lcout => n2189,
            ltout => OPEN,
            carryin => \quad_counter1.n19564\,
            carryout => \quad_counter1.n19565\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_19_lut_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37246\,
            in2 => \N__25316\,
            in3 => \N__25108\,
            lcout => n2188,
            ltout => OPEN,
            carryin => \quad_counter1.n19565\,
            carryout => \quad_counter1.n19566\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_20_lut_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25285\,
            in2 => \N__29049\,
            in3 => \N__25096\,
            lcout => n2187,
            ltout => OPEN,
            carryin => \quad_counter1.n19566\,
            carryout => \quad_counter1.n19567\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_21_lut_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30034\,
            in2 => \N__25317\,
            in3 => \N__25093\,
            lcout => n2186,
            ltout => OPEN,
            carryin => \quad_counter1.n19567\,
            carryout => \quad_counter1.n19568\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_22_lut_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25289\,
            in2 => \N__38934\,
            in3 => \N__25090\,
            lcout => n2185,
            ltout => OPEN,
            carryin => \quad_counter1.n19568\,
            carryout => \quad_counter1.n19569\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_23_lut_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28606\,
            in2 => \N__25318\,
            in3 => \N__25087\,
            lcout => n2184,
            ltout => OPEN,
            carryin => \quad_counter1.n19569\,
            carryout => \quad_counter1.n19570\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_24_lut_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25293\,
            in2 => \N__28487\,
            in3 => \N__25075\,
            lcout => n2183,
            ltout => OPEN,
            carryin => \quad_counter1.n19570\,
            carryout => \quad_counter1.n19571\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_25_lut_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25294\,
            in2 => \N__32900\,
            in3 => \N__25360\,
            lcout => n2182,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \quad_counter1.n19572\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_26_lut_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29958\,
            in2 => \N__25319\,
            in3 => \N__25357\,
            lcout => n2181,
            ltout => OPEN,
            carryin => \quad_counter1.n19572\,
            carryout => \quad_counter1.n19573\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_27_lut_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25298\,
            in2 => \N__33022\,
            in3 => \N__25354\,
            lcout => n2180,
            ltout => OPEN,
            carryin => \quad_counter1.n19573\,
            carryout => \quad_counter1.n19574\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_28_lut_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35645\,
            in2 => \N__25320\,
            in3 => \N__25342\,
            lcout => n2179,
            ltout => OPEN,
            carryin => \quad_counter1.n19574\,
            carryout => \quad_counter1.n19575\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_29_lut_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25302\,
            in2 => \N__30171\,
            in3 => \N__25339\,
            lcout => n2178,
            ltout => OPEN,
            carryin => \quad_counter1.n19575\,
            carryout => \quad_counter1.n19576\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_30_lut_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25246\,
            in2 => \N__36503\,
            in3 => \N__25330\,
            lcout => n2177,
            ltout => OPEN,
            carryin => \quad_counter1.n19576\,
            carryout => \quad_counter1.n19577\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_31_lut_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28954\,
            in2 => \N__25307\,
            in3 => \N__25327\,
            lcout => n2176,
            ltout => OPEN,
            carryin => \quad_counter1.n19577\,
            carryout => \quad_counter1.n19578\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_32_lut_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35517\,
            in2 => \N__25321\,
            in3 => \N__25324\,
            lcout => n2175,
            ltout => OPEN,
            carryin => \quad_counter1.n19578\,
            carryout => \quad_counter1.n19579\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.add_611_33_lut_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25306\,
            in1 => \N__28770\,
            in2 => \_gnd_net_\,
            in3 => \N__25441\,
            lcout => n2174,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20410_4_lut_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__25384\,
            in1 => \N__36765\,
            in2 => \N__27133\,
            in3 => \N__33937\,
            lcout => n24108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__3__5450_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49412\,
            in1 => \N__49007\,
            in2 => \N__41704\,
            in3 => \N__25399\,
            lcout => data_out_frame_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_0__4__5521_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__25425\,
            in1 => \N__37203\,
            in2 => \_gnd_net_\,
            in3 => \N__40171\,
            lcout => data_out_frame_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1600_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26745\,
            in2 => \_gnd_net_\,
            in3 => \N__25607\,
            lcout => \c0.n6_adj_4392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__5__5416_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__49411\,
            in1 => \N__25411\,
            in2 => \N__32740\,
            in3 => \N__49008\,
            lcout => data_out_frame_13_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66780\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n24171_bdd_4_lut_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101111001000"
        )
    port map (
            in0 => \N__25398\,
            in1 => \N__25390\,
            in2 => \N__36833\,
            in3 => \N__34675\,
            lcout => \c0.n24174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__0__5437_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__27156\,
            in1 => \N__49448\,
            in2 => \N__26428\,
            in3 => \N__48847\,
            lcout => data_out_frame_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20163_4_lut_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__26780\,
            in1 => \N__26590\,
            in2 => \N__26864\,
            in3 => \N__25378\,
            lcout => OPEN,
            ltout => \n23858_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_1912_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__25372\,
            in1 => \N__26782\,
            in2 => \N__25363\,
            in3 => \N__25637\,
            lcout => n10_adj_4533,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__2__5451_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49445\,
            in1 => \N__48846\,
            in2 => \N__53476\,
            in3 => \N__25483\,
            lcout => data_out_frame_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__26683\,
            in1 => \N__26781\,
            in2 => \N__25639\,
            in3 => \N__28651\,
            lcout => n10_adj_4535,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_2__I_0_i4_3_lut_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30432\,
            in1 => \N__25522\,
            in2 => \_gnd_net_\,
            in3 => \N__25507\,
            lcout => n4_adj_4554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i3_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__27055\,
            in1 => \N__25489\,
            in2 => \N__27342\,
            in3 => \N__29135\,
            lcout => \r_Tx_Data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_0_i5_3_lut_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25458\,
            in1 => \N__25449\,
            in2 => \_gnd_net_\,
            in3 => \N__39777\,
            lcout => \c0.n5_adj_4422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n24177_bdd_4_lut_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__28996\,
            in1 => \N__25482\,
            in2 => \N__39943\,
            in3 => \N__36896\,
            lcout => OPEN,
            ltout => \c0.n24180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20408_4_lut_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__36897\,
            in1 => \N__30097\,
            in2 => \N__25471\,
            in3 => \N__33963\,
            lcout => n24106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__0__5469_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__49415\,
            in1 => \N__48970\,
            in2 => \N__25462\,
            in3 => \N__39115\,
            lcout => data_out_frame_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__0__5477_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49414\,
            in1 => \N__48969\,
            in2 => \N__39334\,
            in3 => \N__25450\,
            lcout => data_out_frame_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i7_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__27330\,
            in1 => \N__29153\,
            in2 => \N__27070\,
            in3 => \N__25675\,
            lcout => \r_Tx_Data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20155_4_lut_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__25660\,
            in1 => \N__36899\,
            in2 => \N__25654\,
            in3 => \N__33967\,
            lcout => OPEN,
            ltout => \c0.n23850_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20157_4_lut_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__26783\,
            in1 => \N__26873\,
            in2 => \N__25645\,
            in3 => \N__28243\,
            lcout => OPEN,
            ltout => \n23852_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_4_lut_adj_1914_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__25546\,
            in1 => \N__26784\,
            in2 => \N__25642\,
            in3 => \N__25633\,
            lcout => OPEN,
            ltout => \n10_adj_4537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i0_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__27329\,
            in1 => \N__29152\,
            in2 => \N__25549\,
            in3 => \N__25539\,
            lcout => \r_Tx_Data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20412_4_lut_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__27139\,
            in1 => \N__36898\,
            in2 => \N__26197\,
            in3 => \N__33966\,
            lcout => n24110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n24195_bdd_4_lut_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__26966\,
            in1 => \N__27009\,
            in2 => \N__25540\,
            in3 => \N__25528\,
            lcout => n24198,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i0_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30929\,
            in1 => \N__41485\,
            in2 => \_gnd_net_\,
            in3 => \N__30910\,
            lcout => \c0.tx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13175_3_lut_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__27041\,
            in1 => \N__26987\,
            in2 => \_gnd_net_\,
            in3 => \N__29199\,
            lcout => n16706,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20402_4_lut_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__29200\,
            in1 => \N__30451\,
            in2 => \N__30736\,
            in3 => \N__27042\,
            lcout => OPEN,
            ltout => \n24100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i2_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__30452\,
            in1 => \N__30735\,
            in2 => \N__25708\,
            in3 => \N__25705\,
            lcout => \r_Bit_Index_2_adj_4551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i20364_4_lut_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26988\,
            in1 => \N__27040\,
            in2 => \N__30661\,
            in3 => \N__30450\,
            lcout => OPEN,
            ltout => \c0.tx.n23985_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i28_3_lut_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39274\,
            in2 => \N__25699\,
            in3 => \N__30731\,
            lcout => OPEN,
            ltout => \c0.tx.n31_adj_4216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i0_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000001010100"
        )
    port map (
            in0 => \N__41484\,
            in1 => \N__33734\,
            in2 => \N__25696\,
            in3 => \N__30660\,
            lcout => \c0.tx.r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66824\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_86_2_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27602\,
            in2 => \_gnd_net_\,
            in3 => \N__25687\,
            lcout => n187,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \quad_counter0.n19473\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_delay_counter__i1_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27481\,
            in2 => \_gnd_net_\,
            in3 => \N__25684\,
            lcout => \quad_counter0.b_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter0.n19473\,
            carryout => \quad_counter0.n19474\,
            clk => \N__66836\,
            ce => \N__25803\,
            sr => \N__25776\
        );

    \quad_counter0.b_delay_counter__i2_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27468\,
            in2 => \_gnd_net_\,
            in3 => \N__25681\,
            lcout => \quad_counter0.b_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter0.n19474\,
            carryout => \quad_counter0.n19475\,
            clk => \N__66836\,
            ce => \N__25803\,
            sr => \N__25776\
        );

    \quad_counter0.b_delay_counter__i3_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27646\,
            in2 => \_gnd_net_\,
            in3 => \N__25678\,
            lcout => \quad_counter0.b_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter0.n19475\,
            carryout => \quad_counter0.n19476\,
            clk => \N__66836\,
            ce => \N__25803\,
            sr => \N__25776\
        );

    \quad_counter0.b_delay_counter__i4_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27621\,
            in2 => \_gnd_net_\,
            in3 => \N__25735\,
            lcout => \quad_counter0.b_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter0.n19476\,
            carryout => \quad_counter0.n19477\,
            clk => \N__66836\,
            ce => \N__25803\,
            sr => \N__25776\
        );

    \quad_counter0.b_delay_counter__i5_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27454\,
            in2 => \_gnd_net_\,
            in3 => \N__25732\,
            lcout => \quad_counter0.b_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter0.n19477\,
            carryout => \quad_counter0.n19478\,
            clk => \N__66836\,
            ce => \N__25803\,
            sr => \N__25776\
        );

    \quad_counter0.b_delay_counter__i6_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27403\,
            in2 => \_gnd_net_\,
            in3 => \N__25729\,
            lcout => \quad_counter0.b_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter0.n19478\,
            carryout => \quad_counter0.n19479\,
            clk => \N__66836\,
            ce => \N__25803\,
            sr => \N__25776\
        );

    \quad_counter0.b_delay_counter__i7_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34101\,
            in2 => \_gnd_net_\,
            in3 => \N__25726\,
            lcout => \quad_counter0.b_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter0.n19479\,
            carryout => \quad_counter0.n19480\,
            clk => \N__66836\,
            ce => \N__25803\,
            sr => \N__25776\
        );

    \quad_counter0.b_delay_counter__i8_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27417\,
            in2 => \_gnd_net_\,
            in3 => \N__25723\,
            lcout => \quad_counter0.b_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \quad_counter0.n19481\,
            clk => \N__66847\,
            ce => \N__25804\,
            sr => \N__25780\
        );

    \quad_counter0.b_delay_counter__i9_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27634\,
            in2 => \_gnd_net_\,
            in3 => \N__25720\,
            lcout => \quad_counter0.b_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter0.n19481\,
            carryout => \quad_counter0.n19482\,
            clk => \N__66847\,
            ce => \N__25804\,
            sr => \N__25780\
        );

    \quad_counter0.b_delay_counter__i10_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27430\,
            in2 => \_gnd_net_\,
            in3 => \N__25717\,
            lcout => \quad_counter0.b_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter0.n19482\,
            carryout => \quad_counter0.n19483\,
            clk => \N__66847\,
            ce => \N__25804\,
            sr => \N__25780\
        );

    \quad_counter0.b_delay_counter__i11_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27442\,
            in2 => \_gnd_net_\,
            in3 => \N__25714\,
            lcout => \quad_counter0.b_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter0.n19483\,
            carryout => \quad_counter0.n19484\,
            clk => \N__66847\,
            ce => \N__25804\,
            sr => \N__25780\
        );

    \quad_counter0.b_delay_counter__i12_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34080\,
            in2 => \_gnd_net_\,
            in3 => \N__25711\,
            lcout => \quad_counter0.b_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter0.n19484\,
            carryout => \quad_counter0.n19485\,
            clk => \N__66847\,
            ce => \N__25804\,
            sr => \N__25780\
        );

    \quad_counter0.b_delay_counter__i13_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27493\,
            in2 => \_gnd_net_\,
            in3 => \N__25813\,
            lcout => \quad_counter0.b_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter0.n19485\,
            carryout => \quad_counter0.n19486\,
            clk => \N__66847\,
            ce => \N__25804\,
            sr => \N__25780\
        );

    \quad_counter0.b_delay_counter__i14_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34119\,
            in2 => \_gnd_net_\,
            in3 => \N__25810\,
            lcout => \quad_counter0.b_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter0.n19486\,
            carryout => \quad_counter0.n19487\,
            clk => \N__66847\,
            ce => \N__25804\,
            sr => \N__25780\
        );

    \quad_counter0.b_delay_counter__i15_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34062\,
            in2 => \_gnd_net_\,
            in3 => \N__25807\,
            lcout => \quad_counter0.b_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66847\,
            ce => \N__25804\,
            sr => \N__25780\
        );

    \quad_counter0.add_85_2_lut_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27714\,
            in2 => \_gnd_net_\,
            in3 => \N__25753\,
            lcout => n39,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \quad_counter0.n19488\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_delay_counter__i1_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27919\,
            in2 => \_gnd_net_\,
            in3 => \N__25750\,
            lcout => \quad_counter0.a_delay_counter_1\,
            ltout => OPEN,
            carryin => \quad_counter0.n19488\,
            carryout => \quad_counter0.n19489\,
            clk => \N__66857\,
            ce => \N__27772\,
            sr => \N__27747\
        );

    \quad_counter0.a_delay_counter__i2_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27933\,
            in2 => \_gnd_net_\,
            in3 => \N__25747\,
            lcout => \quad_counter0.a_delay_counter_2\,
            ltout => OPEN,
            carryin => \quad_counter0.n19489\,
            carryout => \quad_counter0.n19490\,
            clk => \N__66857\,
            ce => \N__27772\,
            sr => \N__27747\
        );

    \quad_counter0.a_delay_counter__i3_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27958\,
            in2 => \_gnd_net_\,
            in3 => \N__25744\,
            lcout => \quad_counter0.a_delay_counter_3\,
            ltout => OPEN,
            carryin => \quad_counter0.n19490\,
            carryout => \quad_counter0.n19491\,
            clk => \N__66857\,
            ce => \N__27772\,
            sr => \N__27747\
        );

    \quad_counter0.a_delay_counter__i4_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27882\,
            in2 => \_gnd_net_\,
            in3 => \N__25741\,
            lcout => \quad_counter0.a_delay_counter_4\,
            ltout => OPEN,
            carryin => \quad_counter0.n19491\,
            carryout => \quad_counter0.n19492\,
            clk => \N__66857\,
            ce => \N__27772\,
            sr => \N__27747\
        );

    \quad_counter0.a_delay_counter__i5_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27907\,
            in2 => \_gnd_net_\,
            in3 => \N__25738\,
            lcout => \quad_counter0.a_delay_counter_5\,
            ltout => OPEN,
            carryin => \quad_counter0.n19492\,
            carryout => \quad_counter0.n19493\,
            clk => \N__66857\,
            ce => \N__27772\,
            sr => \N__27747\
        );

    \quad_counter0.a_delay_counter__i6_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28098\,
            in2 => \_gnd_net_\,
            in3 => \N__25840\,
            lcout => \quad_counter0.a_delay_counter_6\,
            ltout => OPEN,
            carryin => \quad_counter0.n19493\,
            carryout => \quad_counter0.n19494\,
            clk => \N__66857\,
            ce => \N__27772\,
            sr => \N__27747\
        );

    \quad_counter0.a_delay_counter__i7_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27672\,
            in2 => \_gnd_net_\,
            in3 => \N__25837\,
            lcout => \quad_counter0.a_delay_counter_7\,
            ltout => OPEN,
            carryin => \quad_counter0.n19494\,
            carryout => \quad_counter0.n19495\,
            clk => \N__66857\,
            ce => \N__27772\,
            sr => \N__27747\
        );

    \quad_counter0.a_delay_counter__i8_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27946\,
            in2 => \_gnd_net_\,
            in3 => \N__25834\,
            lcout => \quad_counter0.a_delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_10_25_0_\,
            carryout => \quad_counter0.n19496\,
            clk => \N__66865\,
            ce => \N__27768\,
            sr => \N__27748\
        );

    \quad_counter0.a_delay_counter__i9_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28084\,
            in2 => \_gnd_net_\,
            in3 => \N__25831\,
            lcout => \quad_counter0.a_delay_counter_9\,
            ltout => OPEN,
            carryin => \quad_counter0.n19496\,
            carryout => \quad_counter0.n19497\,
            clk => \N__66865\,
            ce => \N__27768\,
            sr => \N__27748\
        );

    \quad_counter0.a_delay_counter__i10_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27658\,
            in2 => \_gnd_net_\,
            in3 => \N__25828\,
            lcout => \quad_counter0.a_delay_counter_10\,
            ltout => OPEN,
            carryin => \quad_counter0.n19497\,
            carryout => \quad_counter0.n19498\,
            clk => \N__66865\,
            ce => \N__27768\,
            sr => \N__27748\
        );

    \quad_counter0.a_delay_counter__i11_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27895\,
            in2 => \_gnd_net_\,
            in3 => \N__25825\,
            lcout => \quad_counter0.a_delay_counter_11\,
            ltout => OPEN,
            carryin => \quad_counter0.n19498\,
            carryout => \quad_counter0.n19499\,
            clk => \N__66865\,
            ce => \N__27768\,
            sr => \N__27748\
        );

    \quad_counter0.a_delay_counter__i12_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28123\,
            in2 => \_gnd_net_\,
            in3 => \N__25822\,
            lcout => \quad_counter0.a_delay_counter_12\,
            ltout => OPEN,
            carryin => \quad_counter0.n19499\,
            carryout => \quad_counter0.n19500\,
            clk => \N__66865\,
            ce => \N__27768\,
            sr => \N__27748\
        );

    \quad_counter0.a_delay_counter__i13_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28111\,
            in2 => \_gnd_net_\,
            in3 => \N__25819\,
            lcout => \quad_counter0.a_delay_counter_13\,
            ltout => OPEN,
            carryin => \quad_counter0.n19500\,
            carryout => \quad_counter0.n19501\,
            clk => \N__66865\,
            ce => \N__27768\,
            sr => \N__27748\
        );

    \quad_counter0.a_delay_counter__i14_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27697\,
            in2 => \_gnd_net_\,
            in3 => \N__25816\,
            lcout => \quad_counter0.a_delay_counter_14\,
            ltout => OPEN,
            carryin => \quad_counter0.n19501\,
            carryout => \quad_counter0.n19502\,
            clk => \N__66865\,
            ce => \N__27768\,
            sr => \N__27748\
        );

    \quad_counter0.a_delay_counter__i15_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27685\,
            in2 => \_gnd_net_\,
            in3 => \N__25888\,
            lcout => \quad_counter0.a_delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66865\,
            ce => \N__27768\,
            sr => \N__27748\
        );

    \c0.i1_2_lut_3_lut_adj_1876_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__31485\,
            in1 => \N__29564\,
            in2 => \_gnd_net_\,
            in3 => \N__34426\,
            lcout => \c0.n22317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32792\,
            in1 => \N__35057\,
            in2 => \_gnd_net_\,
            in3 => \N__29788\,
            lcout => OPEN,
            ltout => \c0.n18_adj_4414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1805_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31489\,
            in1 => \N__25885\,
            in2 => \N__25879\,
            in3 => \N__28189\,
            lcout => \c0.n26_adj_4504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1396_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__32565\,
            in1 => \N__32516\,
            in2 => \_gnd_net_\,
            in3 => \N__34828\,
            lcout => OPEN,
            ltout => \c0.n23550_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1804_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25876\,
            in1 => \N__34476\,
            in2 => \N__25870\,
            in3 => \N__31798\,
            lcout => OPEN,
            ltout => \c0.n22_adj_4503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__1__5292_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28012\,
            in1 => \N__29292\,
            in2 => \N__25867\,
            in3 => \N__25864\,
            lcout => \c0.data_out_frame_29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66659\,
            ce => \N__40953\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i26_3_lut_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26148\,
            in1 => \N__26119\,
            in2 => \_gnd_net_\,
            in3 => \N__39835\,
            lcout => \c0.n26_adj_4517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1408_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__32039\,
            in1 => \N__32790\,
            in2 => \_gnd_net_\,
            in3 => \N__31964\,
            lcout => \c0.n10462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1400_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31927\,
            in2 => \_gnd_net_\,
            in3 => \N__32115\,
            lcout => OPEN,
            ltout => \c0.n21305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__2__5299_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26113\,
            in1 => \N__28035\,
            in2 => \N__26122\,
            in3 => \N__29562\,
            lcout => \c0.data_out_frame_28_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66664\,
            ce => \N__40951\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1889_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__32149\,
            in1 => \N__29353\,
            in2 => \_gnd_net_\,
            in3 => \N__32206\,
            lcout => \c0.n6_adj_4515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1870_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28171\,
            in1 => \N__32791\,
            in2 => \N__32046\,
            in3 => \N__32517\,
            lcout => \c0.n12532\,
            ltout => \c0.n12532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1641_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__29423\,
            in1 => \_gnd_net_\,
            in2 => \N__26104\,
            in3 => \N__32205\,
            lcout => \c0.n22126\,
            ltout => \c0.n22126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__4__5297_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31840\,
            in2 => \N__26101\,
            in3 => \N__34850\,
            lcout => \c0.data_out_frame_28_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66664\,
            ce => \N__40951\,
            sr => \_gnd_net_\
        );

    \quad_counter1.i10_4_lut_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26086\,
            in1 => \N__26070\,
            in2 => \N__26059\,
            in3 => \N__26043\,
            lcout => \quad_counter1.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.quadA_I_0_73_2_lut_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25966\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25991\,
            lcout => \a_delay_counter_15__N_4124_adj_4547\,
            ltout => \a_delay_counter_15__N_4124_adj_4547_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110000"
        )
    port map (
            in0 => \N__25992\,
            in1 => \N__25965\,
            in2 => \N__25921\,
            in3 => \N__25918\,
            lcout => n14228,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_2_lut_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41913\,
            in2 => \_gnd_net_\,
            in3 => \N__43079\,
            lcout => \c0.n161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__2__5291_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__28269\,
            in1 => \N__49410\,
            in2 => \N__26152\,
            in3 => \N__49019\,
            lcout => data_out_frame_29_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1724_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31926\,
            in1 => \N__32116\,
            in2 => \N__29377\,
            in3 => \N__32148\,
            lcout => \data_out_frame_28__3__N_1881\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_rx_data_ready_prev_5283_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43110\,
            lcout => \c0.FRAME_MATCHER_rx_data_ready_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_DV_52_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__57028\,
            in1 => \N__43111\,
            in2 => \N__54343\,
            in3 => \N__56950\,
            lcout => rx_data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i9_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38505\,
            in1 => \N__26137\,
            in2 => \_gnd_net_\,
            in3 => \N__32286\,
            lcout => encoder1_position_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__3__5290_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__49569\,
            in1 => \N__26622\,
            in2 => \N__49047\,
            in3 => \N__29293\,
            lcout => data_out_frame_29_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1454_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26482\,
            in1 => \N__35149\,
            in2 => \N__28965\,
            in3 => \N__38870\,
            lcout => \c0.n13079\,
            ltout => \c0.n13079_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1413_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35911\,
            in1 => \N__26161\,
            in2 => \N__26125\,
            in3 => \N__35723\,
            lcout => \c0.n21056\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i3_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43109\,
            in1 => \N__30611\,
            in2 => \_gnd_net_\,
            in3 => \N__30338\,
            lcout => data_in_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1407_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26335\,
            in1 => \N__26230\,
            in2 => \N__26224\,
            in3 => \N__35839\,
            lcout => \c0.n20175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_0_i11_3_lut_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39822\,
            in1 => \N__26211\,
            in2 => \_gnd_net_\,
            in3 => \N__35341\,
            lcout => \c0.n11_adj_4424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1485_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26334\,
            in2 => \_gnd_net_\,
            in3 => \N__35449\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4335_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1486_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35030\,
            in1 => \N__28678\,
            in2 => \N__26179\,
            in3 => \N__26423\,
            lcout => \c0.n21229\,
            ltout => \c0.n21229_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1685_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__28311\,
            in1 => \_gnd_net_\,
            in2 => \N__26176\,
            in3 => \N__31256\,
            lcout => \c0.n21152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i12_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34631\,
            in1 => \N__26173\,
            in2 => \_gnd_net_\,
            in3 => \N__38395\,
            lcout => encoder1_position_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66699\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1705_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33163\,
            in1 => \N__26325\,
            in2 => \N__28786\,
            in3 => \N__26419\,
            lcout => \c0.n6_adj_4309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__5__5448_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49561\,
            in1 => \N__48968\,
            in2 => \N__36082\,
            in3 => \N__27108\,
            lcout => data_out_frame_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1429_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__33161\,
            in1 => \N__26418\,
            in2 => \_gnd_net_\,
            in3 => \N__26324\,
            lcout => \c0.n22293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1483_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28660\,
            in1 => \N__35445\,
            in2 => \N__37072\,
            in3 => \N__33160\,
            lcout => \c0.n20330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38497\,
            in1 => \N__26344\,
            in2 => \_gnd_net_\,
            in3 => \N__32789\,
            lcout => encoder1_position_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1414_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35519\,
            in2 => \_gnd_net_\,
            in3 => \N__33162\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4310_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1415_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__26481\,
            in1 => \N__38179\,
            in2 => \N__26338\,
            in3 => \N__38875\,
            lcout => \c0.n22037\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__7__5422_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__49002\,
            in1 => \N__49380\,
            in2 => \N__26278\,
            in3 => \N__26326\,
            lcout => data_out_frame_12_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_7_i11_3_lut_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32068\,
            in1 => \N__26274\,
            in2 => \_gnd_net_\,
            in3 => \N__39756\,
            lcout => \c0.n11_adj_4360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i8_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38498\,
            in1 => \N__26254\,
            in2 => \_gnd_net_\,
            in3 => \N__35391\,
            lcout => encoder1_position_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_4_i5_3_lut_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26238\,
            in1 => \N__30388\,
            in2 => \_gnd_net_\,
            in3 => \N__39757\,
            lcout => \c0.n5_adj_4227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__4__5465_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__49004\,
            in1 => \N__49382\,
            in2 => \N__36136\,
            in3 => \N__26239\,
            lcout => data_out_frame_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__3__5298_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__49003\,
            in1 => \N__49381\,
            in2 => \N__26608\,
            in3 => \N__28065\,
            lcout => data_out_frame_28_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1849_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39499\,
            in1 => \N__35418\,
            in2 => \N__35794\,
            in3 => \N__38586\,
            lcout => \c0.n10422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.encoder0_position_27__I_0_2_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33386\,
            in2 => \_gnd_net_\,
            in3 => \N__40056\,
            lcout => \c0.data_out_frame_29__7__N_850\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20186_3_lut_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26464\,
            in1 => \N__26379\,
            in2 => \_gnd_net_\,
            in3 => \N__39805\,
            lcout => \c0.n23881\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i16_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38491\,
            in1 => \N__26434\,
            in2 => \_gnd_net_\,
            in3 => \N__26417\,
            lcout => encoder1_position_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__4__5441_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__49553\,
            in1 => \N__26380\,
            in2 => \N__36505\,
            in3 => \N__48939\,
            lcout => data_out_frame_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i11_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43154\,
            in1 => \N__28846\,
            in2 => \_gnd_net_\,
            in3 => \N__30328\,
            lcout => data_in_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__2__5467_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49554\,
            in1 => \N__48938\,
            in2 => \N__41758\,
            in3 => \N__26364\,
            lcout => data_out_frame_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i17_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26350\,
            in1 => \N__37250\,
            in2 => \_gnd_net_\,
            in3 => \N__38492\,
            lcout => encoder1_position_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i19_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43193\,
            in1 => \N__28845\,
            in2 => \_gnd_net_\,
            in3 => \N__36595\,
            lcout => data_in_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i21_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28610\,
            in1 => \N__26644\,
            in2 => \_gnd_net_\,
            in3 => \N__38499\,
            lcout => encoder1_position_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i23_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38500\,
            in1 => \N__26638\,
            in2 => \_gnd_net_\,
            in3 => \N__32892\,
            lcout => encoder1_position_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i29_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28958\,
            in1 => \N__26632\,
            in2 => \_gnd_net_\,
            in3 => \N__38501\,
            lcout => encoder1_position_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i26_3_lut_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39807\,
            in1 => \N__26626\,
            in2 => \_gnd_net_\,
            in3 => \N__26607\,
            lcout => \c0.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i30_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38502\,
            in1 => \N__26581\,
            in2 => \_gnd_net_\,
            in3 => \N__35518\,
            lcout => encoder1_position_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66753\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_5_i5_3_lut_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26575\,
            in1 => \N__36286\,
            in2 => \_gnd_net_\,
            in3 => \N__39806\,
            lcout => \c0.n5_adj_4346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__3__5474_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49517\,
            in1 => \N__49006\,
            in2 => \N__33394\,
            in3 => \N__27210\,
            lcout => data_out_frame_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__7__5446_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__49005\,
            in1 => \N__49413\,
            in2 => \N__33253\,
            in3 => \N__26541\,
            lcout => data_out_frame_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.o_Tx_Serial_45_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__26493\,
            in1 => \N__30748\,
            in2 => \_gnd_net_\,
            in3 => \N__41491\,
            lcout => tx_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66767\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1604_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__33864\,
            in1 => \N__39626\,
            in2 => \N__36817\,
            in3 => \N__26938\,
            lcout => OPEN,
            ltout => \c0.n23574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1675_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27310\,
            in1 => \N__26932\,
            in2 => \N__26914\,
            in3 => \N__26911\,
            lcout => \c0.n38_adj_4387\,
            ltout => \c0.n38_adj_4387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20438_2_lut_3_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39273\,
            in2 => \N__26896\,
            in3 => \N__37147\,
            lcout => \c0.tx_transmit_N_3651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__5__5456_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__48978\,
            in1 => \N__49519\,
            in2 => \N__27091\,
            in3 => \N__35725\,
            lcout => data_out_frame_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__5__5432_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49518\,
            in1 => \N__48979\,
            in2 => \N__28615\,
            in3 => \N__27123\,
            lcout => data_out_frame_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__2__5483_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__48976\,
            in1 => \N__39487\,
            in2 => \N__49551\,
            in3 => \N__26889\,
            lcout => data_out_frame_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20169_4_lut_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__27991\,
            in1 => \N__33988\,
            in2 => \N__26863\,
            in3 => \N__26779\,
            lcout => n23864,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__6__5479_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__48977\,
            in1 => \N__42307\,
            in2 => \N__49552\,
            in3 => \N__26673\,
            lcout => data_out_frame_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i11_3_lut_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39749\,
            in1 => \N__26659\,
            in2 => \_gnd_net_\,
            in3 => \N__28911\,
            lcout => \c0.n11_adj_4218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_20456_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__36894\,
            in1 => \N__28929\,
            in2 => \N__27124\,
            in3 => \N__39750\,
            lcout => OPEN,
            ltout => \c0.n24141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n24141_bdd_4_lut_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__36895\,
            in1 => \N__27112\,
            in2 => \N__27094\,
            in3 => \N__27087\,
            lcout => \c0.n24144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_Bit_Index_2__bdd_4_lut_20490_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__27066\,
            in1 => \N__27054\,
            in2 => \N__26978\,
            in3 => \N__27043\,
            lcout => OPEN,
            ltout => \n24189_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n24189_bdd_4_lut_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__27016\,
            in1 => \N__27255\,
            in2 => \N__26992\,
            in3 => \N__26970\,
            lcout => n24192,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i8_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30502\,
            in1 => \N__43155\,
            in2 => \_gnd_net_\,
            in3 => \N__27245\,
            lcout => data_in_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i0_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011001100"
        )
    port map (
            in0 => \N__30729\,
            in1 => \N__30443\,
            in2 => \_gnd_net_\,
            in3 => \N__29193\,
            lcout => \r_Bit_Index_0_adj_4553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Bit_Index_i1_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101000100010"
        )
    port map (
            in0 => \N__26971\,
            in1 => \N__29192\,
            in2 => \N__30453\,
            in3 => \N__30730\,
            lcout => \r_Bit_Index_1_adj_4552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1694_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__43045\,
            in1 => \N__36994\,
            in2 => \N__27247\,
            in3 => \N__29069\,
            lcout => \c0.n16_adj_4476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Data_i1_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__27256\,
            in1 => \N__27352\,
            in2 => \N__27343\,
            in3 => \N__29117\,
            lcout => \r_Tx_Data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__43044\,
            in1 => \N__29068\,
            in2 => \N__27246\,
            in3 => \N__30618\,
            lcout => \c0.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1888_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43411\,
            in1 => \N__37799\,
            in2 => \N__41011\,
            in3 => \N__34247\,
            lcout => \c0.n20_adj_4482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__3__5482_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49549\,
            in1 => \N__48975\,
            in2 => \N__41815\,
            in3 => \N__27228\,
            lcout => data_out_frame_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_3_i5_3_lut_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39799\,
            in1 => \N__37102\,
            in2 => \_gnd_net_\,
            in3 => \N__27211\,
            lcout => \c0.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__5__5480_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__48974\,
            in1 => \N__49550\,
            in2 => \N__27180\,
            in3 => \N__40213\,
            lcout => data_out_frame_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_20471_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__39800\,
            in1 => \N__27157\,
            in2 => \N__29089\,
            in3 => \N__36887\,
            lcout => OPEN,
            ltout => \c0.n24165_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n24165_bdd_4_lut_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__36888\,
            in1 => \N__34030\,
            in2 => \N__27142\,
            in3 => \N__37018\,
            lcout => \c0.n24168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i22_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34302\,
            in2 => \_gnd_net_\,
            in3 => \N__52858\,
            lcout => \c0.FRAME_MATCHER_state_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66813\,
            ce => 'H',
            sr => \N__29173\
        );

    \quad_counter0.i3_4_lut_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27358\,
            in1 => \N__27973\,
            in2 => \N__27868\,
            in3 => \N__27503\,
            lcout => count_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i9_4_lut_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__27645\,
            in1 => \N__27633\,
            in2 => \N__27622\,
            in3 => \N__27606\,
            lcout => \quad_counter0.n25_adj_4201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i1072_1_lut_2_lut_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27972\,
            in2 => \_gnd_net_\,
            in3 => \N__27864\,
            lcout => \quad_counter0.n2227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.B_65_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101000"
        )
    port map (
            in0 => \N__27504\,
            in1 => \N__27583\,
            in2 => \N__27538\,
            in3 => \N__27372\,
            lcout => \B_filtered\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66825\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.B_delayed_68_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27505\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quad_counter0.B_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66825\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i12_4_lut_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__27492\,
            in1 => \N__27480\,
            in2 => \N__27469\,
            in3 => \N__27453\,
            lcout => \quad_counter0.n28_adj_4198\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i10_4_lut_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27441\,
            in1 => \N__27429\,
            in2 => \N__27418\,
            in3 => \N__27402\,
            lcout => OPEN,
            ltout => \quad_counter0.n26_adj_4199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i15_4_lut_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27391\,
            in1 => \N__34048\,
            in2 => \N__27385\,
            in3 => \N__27382\,
            lcout => n12909,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.A_delayed_67_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27859\,
            lcout => \quad_counter0.A_delayed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.A_filtered_I_0_2_lut_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27971\,
            in2 => \_gnd_net_\,
            in3 => \N__27858\,
            lcout => \quad_counter0.count_direction\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i12_4_lut_adj_1161_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__27957\,
            in1 => \N__27945\,
            in2 => \N__27934\,
            in3 => \N__27918\,
            lcout => \quad_counter0.n28_adj_4202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i9_4_lut_adj_1164_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__27906\,
            in1 => \N__27894\,
            in2 => \N__27883\,
            in3 => \N__27713\,
            lcout => \quad_counter0.n25_adj_4205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.A_63_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001000000"
        )
    port map (
            in0 => \N__28132\,
            in1 => \N__27832\,
            in2 => \N__27799\,
            in3 => \N__27863\,
            lcout => \A_filtered\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1764_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__53012\,
            in1 => \N__37846\,
            in2 => \_gnd_net_\,
            in3 => \N__53195\,
            lcout => \c0.n21362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__27831\,
            in1 => \N__27795\,
            in2 => \_gnd_net_\,
            in3 => \N__28131\,
            lcout => n14421,
            ltout => \n14421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_delay_counter__i0_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__27746\,
            in1 => \N__27724\,
            in2 => \N__27718\,
            in3 => \N__27715\,
            lcout => a_delay_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i11_4_lut_adj_1163_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27696\,
            in1 => \N__27684\,
            in2 => \N__27673\,
            in3 => \N__27657\,
            lcout => OPEN,
            ltout => \quad_counter0.n27_adj_4204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i15_4_lut_adj_1165_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28147\,
            in1 => \N__28072\,
            in2 => \N__28141\,
            in3 => \N__28138\,
            lcout => n9821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i10_4_lut_adj_1162_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28122\,
            in1 => \N__28110\,
            in2 => \N__28099\,
            in3 => \N__28083\,
            lcout => \quad_counter0.n26_adj_4203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__1__5300_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28066\,
            in1 => \N__30981\,
            in2 => \N__28042\,
            in3 => \N__29215\,
            lcout => \c0.data_out_frame_28_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66638\,
            ce => \N__40952\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1801_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31458\,
            in2 => \_gnd_net_\,
            in3 => \N__32212\,
            lcout => \c0.n21062\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1582_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31770\,
            in1 => \N__29563\,
            in2 => \N__32389\,
            in3 => \N__35614\,
            lcout => \c0.n20376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_1_i26_3_lut_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28006\,
            in1 => \N__27997\,
            in2 => \_gnd_net_\,
            in3 => \N__39833\,
            lcout => \c0.n26_adj_4519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1864_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31631\,
            in1 => \N__29805\,
            in2 => \N__31420\,
            in3 => \N__31132\,
            lcout => \c0.n12542\,
            ltout => \c0.n12542_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_3_lut_4_lut_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31683\,
            in1 => \N__29270\,
            in2 => \N__27976\,
            in3 => \N__31632\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1495_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31089\,
            in1 => \N__29209\,
            in2 => \N__28192\,
            in3 => \N__31569\,
            lcout => \data_out_frame_29__2__N_1749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1863_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__29602\,
            in1 => \N__29804\,
            in2 => \N__31419\,
            in3 => \N__31131\,
            lcout => \c0.n20320\,
            ltout => \c0.n20320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1880_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34399\,
            in1 => \N__31682\,
            in2 => \N__28183\,
            in3 => \N__31415\,
            lcout => \c0.n21219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1845_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29354\,
            in2 => \_gnd_net_\,
            in3 => \N__29416\,
            lcout => \c0.n21128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1707_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35122\,
            in1 => \N__29695\,
            in2 => \N__28356\,
            in3 => \N__53386\,
            lcout => \c0.n22180\,
            ltout => \c0.n22180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_4_lut_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28352\,
            in2 => \N__28180\,
            in3 => \N__28169\,
            lcout => \c0.n10498\,
            ltout => \c0.n10498_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1835_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28498\,
            in1 => \N__28153\,
            in2 => \N__28177\,
            in3 => \N__32931\,
            lcout => \c0.n21058\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1591_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31285\,
            in1 => \N__31630\,
            in2 => \N__31348\,
            in3 => \N__31130\,
            lcout => \c0.n22024\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1840_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31209\,
            in2 => \_gnd_net_\,
            in3 => \N__34344\,
            lcout => \c0.n20253\,
            ltout => \c0.n20253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1834_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28363\,
            in1 => \N__31839\,
            in2 => \N__28174\,
            in3 => \N__28170\,
            lcout => \c0.n15_adj_4513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1811_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__32505\,
            in1 => \N__29600\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \c0.n21998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1411_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__53387\,
            in1 => \_gnd_net_\,
            in2 => \N__29705\,
            in3 => \_gnd_net_\,
            lcout => \c0.n22066\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1610_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28344\,
            in1 => \N__32035\,
            in2 => \N__32799\,
            in3 => \N__31272\,
            lcout => \c0.n10496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1484_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__31273\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28345\,
            lcout => OPEN,
            ltout => \c0.n21071_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__0__5293_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28225\,
            in1 => \N__28255\,
            in2 => \N__28273\,
            in3 => \N__28270\,
            lcout => \c0.data_out_frame_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66665\,
            ce => \N__40944\,
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1799_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31438\,
            in1 => \N__29608\,
            in2 => \N__32449\,
            in3 => \N__31152\,
            lcout => \c0.n17_adj_4501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_0_i26_3_lut_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28249\,
            in1 => \N__29479\,
            in2 => \_gnd_net_\,
            in3 => \N__39834\,
            lcout => \c0.n26_adj_4423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1798_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32617\,
            in1 => \N__32210\,
            in2 => \N__31349\,
            in3 => \N__29767\,
            lcout => \c0.n16_adj_4500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1615_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28392\,
            in1 => \N__35386\,
            in2 => \N__28218\,
            in3 => \N__28489\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4313_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1420_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35310\,
            in1 => \N__34870\,
            in2 => \N__28375\,
            in3 => \N__38965\,
            lcout => \c0.n21156\,
            ltout => \c0.n21156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1713_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29854\,
            in2 => \N__28372\,
            in3 => \N__34793\,
            lcout => \c0.n21231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_adj_1613_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28393\,
            in1 => \N__28488\,
            in2 => \N__36078\,
            in3 => \N__35385\,
            lcout => \c0.n10_adj_4330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1464_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32857\,
            in1 => \N__32823\,
            in2 => \N__35283\,
            in3 => \N__28391\,
            lcout => \c0.n21175\,
            ltout => \c0.n21175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1712_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__29829\,
            in1 => \N__34794\,
            in2 => \N__28369\,
            in3 => \N__31151\,
            lcout => \c0.n21150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1423_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35309\,
            in1 => \N__39035\,
            in2 => \_gnd_net_\,
            in3 => \N__28624\,
            lcout => \c0.n22991\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1652_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29978\,
            in1 => \N__34622\,
            in2 => \N__31892\,
            in3 => \N__35609\,
            lcout => \c0.n20276\,
            ltout => \c0.n20276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1808_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28366\,
            in3 => \N__31257\,
            lcout => \c0.n21116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1674_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29980\,
            in1 => \N__34623\,
            in2 => \_gnd_net_\,
            in3 => \N__35610\,
            lcout => OPEN,
            ltout => \c0.n21110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1886_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35120\,
            in1 => \N__32371\,
            in2 => \N__28501\,
            in3 => \N__31886\,
            lcout => \c0.n14_adj_4514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1428_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32273\,
            in2 => \_gnd_net_\,
            in3 => \N__28474\,
            lcout => \c0.n22277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i4_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35121\,
            in1 => \N__38396\,
            in2 => \_gnd_net_\,
            in3 => \N__28438\,
            lcout => encoder1_position_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1394_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29977\,
            in1 => \N__36454\,
            in2 => \_gnd_net_\,
            in3 => \N__38063\,
            lcout => \c0.n21065\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1728_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34621\,
            in1 => \N__29979\,
            in2 => \N__32975\,
            in3 => \N__32856\,
            lcout => \c0.n21166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1449_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29664\,
            in1 => \N__31252\,
            in2 => \N__32901\,
            in3 => \N__29998\,
            lcout => \c0.n17_adj_4323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1839_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41872\,
            in1 => \N__39056\,
            in2 => \_gnd_net_\,
            in3 => \N__39495\,
            lcout => \c0.n22102\,
            ltout => \c0.n22102_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1451_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28422\,
            in1 => \N__38515\,
            in2 => \N__28405\,
            in3 => \N__28402\,
            lcout => OPEN,
            ltout => \c0.n15_adj_4325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1452_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41293\,
            in1 => \N__31757\,
            in2 => \N__28396\,
            in3 => \N__35461\,
            lcout => \c0.n21041\,
            ltout => \c0.n21041_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1453_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__35369\,
            in1 => \_gnd_net_\,
            in2 => \N__28378\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \c0.n22361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1422_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__28633\,
            in1 => \N__41682\,
            in2 => \N__28627\,
            in3 => \N__35932\,
            lcout => \c0.n10_adj_4314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__6__5455_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49335\,
            in1 => \N__49001\,
            in2 => \N__35899\,
            in3 => \N__28566\,
            lcout => data_out_frame_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__1__5460_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__48999\,
            in1 => \N__49336\,
            in2 => \N__38728\,
            in3 => \N__33474\,
            lcout => data_out_frame_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1689_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28611\,
            in1 => \N__36558\,
            in2 => \_gnd_net_\,
            in3 => \N__38648\,
            lcout => \c0.n22408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i3_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42202\,
            in1 => \N__33103\,
            in2 => \_gnd_net_\,
            in3 => \N__41673\,
            lcout => encoder0_position_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n24153_bdd_4_lut_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__29898\,
            in1 => \N__28582\,
            in2 => \N__28567\,
            in3 => \N__36908\,
            lcout => \c0.n24156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__6__5423_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49334\,
            in1 => \N__49000\,
            in2 => \N__29665\,
            in3 => \N__28539\,
            lcout => data_out_frame_12_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66713\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1445_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36504\,
            in1 => \N__29937\,
            in2 => \N__41683\,
            in3 => \N__38724\,
            lcout => \c0.n19_adj_4319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__3__5434_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__48945\,
            in1 => \N__49403\,
            in2 => \N__28521\,
            in3 => \N__30029\,
            lcout => data_out_frame_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i4_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43192\,
            in1 => \N__28811\,
            in2 => \_gnd_net_\,
            in3 => \N__36382\,
            lcout => data_in_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i24_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38503\,
            in1 => \N__28690\,
            in2 => \_gnd_net_\,
            in3 => \N__29947\,
            lcout => encoder1_position_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66727\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1469_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37060\,
            in2 => \_gnd_net_\,
            in3 => \N__35895\,
            lcout => \c0.n22224\,
            ltout => \c0.n22224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1471_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29042\,
            in1 => \N__28639\,
            in2 => \N__28666\,
            in3 => \N__36028\,
            lcout => \c0.n13349\,
            ltout => \c0.n13349_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1482_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28663\,
            in3 => \N__28781\,
            lcout => \c0.n6_adj_4334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1693_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44619\,
            in1 => \N__41871\,
            in2 => \_gnd_net_\,
            in3 => \N__41750\,
            lcout => \c0.n22412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i14_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__43219\,
            in1 => \_gnd_net_\,
            in2 => \N__28897\,
            in3 => \N__36426\,
            lcout => data_in_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66740\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20406_4_lut_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__33460\,
            in1 => \N__36889\,
            in2 => \N__34696\,
            in3 => \N__33968\,
            lcout => n24104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1470_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35772\,
            in2 => \_gnd_net_\,
            in3 => \N__38246\,
            lcout => \c0.n22405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__1__5444_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__49391\,
            in1 => \N__36924\,
            in2 => \N__33017\,
            in3 => \N__48891\,
            lcout => data_out_frame_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66740\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__7__5438_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__48889\,
            in1 => \N__49393\,
            in2 => \N__28741\,
            in3 => \N__28782\,
            lcout => data_out_frame_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66740\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__7__5454_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49392\,
            in1 => \N__48890\,
            in2 => \N__36265\,
            in3 => \N__28722\,
            lcout => data_out_frame_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66740\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1547_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__36427\,
            in1 => \N__30278\,
            in2 => \N__36961\,
            in3 => \N__30580\,
            lcout => \c0.n19_adj_4367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i15_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30279\,
            in1 => \N__36960\,
            in2 => \_gnd_net_\,
            in3 => \N__43260\,
            lcout => data_in_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i16_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43258\,
            in1 => \N__36625\,
            in2 => \_gnd_net_\,
            in3 => \N__30498\,
            lcout => data_in_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__7__5430_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__48933\,
            in1 => \N__32893\,
            in2 => \N__49451\,
            in3 => \N__28704\,
            lcout => data_out_frame_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i20_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43259\,
            in1 => \N__34192\,
            in2 => \_gnd_net_\,
            in3 => \N__29074\,
            lcout => data_in_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1771_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__30557\,
            in1 => \N__28888\,
            in2 => \N__41960\,
            in3 => \N__41994\,
            lcout => \c0.n15_adj_4496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i6_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28889\,
            in1 => \N__43261\,
            in2 => \_gnd_net_\,
            in3 => \N__30300\,
            lcout => data_in_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__3__5426_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__48934\,
            in1 => \N__32979\,
            in2 => \N__49452\,
            in3 => \N__28912\,
            lcout => data_out_frame_12_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1756_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__41998\,
            in1 => \N__28844\,
            in2 => \N__30256\,
            in3 => \N__28864\,
            lcout => OPEN,
            ltout => \c0.n7_adj_4492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1761_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__40242\,
            in1 => \N__28857\,
            in2 => \N__28900\,
            in3 => \N__28870\,
            lcout => \c0.n63_adj_4301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_2_lut_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28896\,
            in2 => \_gnd_net_\,
            in3 => \N__30366\,
            lcout => \c0.n9_adj_4493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i7_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28858\,
            in1 => \N__30283\,
            in2 => \_gnd_net_\,
            in3 => \N__43262\,
            lcout => data_in_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66768\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1706_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__30550\,
            in1 => \N__41967\,
            in2 => \N__28822\,
            in3 => \N__30591\,
            lcout => \c0.n23600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1769_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__28856\,
            in1 => \N__40241\,
            in2 => \_gnd_net_\,
            in3 => \N__30252\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4495_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1772_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__28843\,
            in1 => \N__28818\,
            in2 => \N__28795\,
            in3 => \N__28792\,
            lcout => \c0.n21767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1773_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35253\,
            in2 => \_gnd_net_\,
            in3 => \N__34193\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4231_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1241_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__34165\,
            in1 => \N__36993\,
            in2 => \N__29164\,
            in3 => \N__29161\,
            lcout => \c0.n13003\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_3_lut_4_lut_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__41445\,
            in1 => \N__39268\,
            in2 => \N__33771\,
            in3 => \N__30711\,
            lcout => n9539,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__0__5445_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49512\,
            in1 => \N__48944\,
            in2 => \N__29962\,
            in3 => \N__29088\,
            lcout => data_out_frame_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i28_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__64872\,
            in1 => \N__43267\,
            in2 => \_gnd_net_\,
            in3 => \N__29070\,
            lcout => data_in_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i9_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__43266\,
            in1 => \_gnd_net_\,
            in2 => \N__30558\,
            in3 => \N__36220\,
            lcout => data_in_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__2__5435_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__48943\,
            in1 => \N__49513\,
            in2 => \N__29050\,
            in3 => \N__29010\,
            lcout => data_out_frame_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_20481_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__30133\,
            in1 => \N__36883\,
            in2 => \N__29011\,
            in3 => \N__39804\,
            lcout => \c0.n24177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__0__5485_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49476\,
            in1 => \N__48896\,
            in2 => \N__44623\,
            in3 => \N__28983\,
            lcout => data_out_frame_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__5__5440_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__49475\,
            in1 => \N__28966\,
            in2 => \N__28930\,
            in3 => \N__48897\,
            lcout => data_out_frame_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_1181_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33768\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30643\,
            lcout => OPEN,
            ltout => \c0.tx.n16631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_adj_1187_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__30707\,
            in1 => \N__41443\,
            in2 => \N__29203\,
            in3 => \N__33706\,
            lcout => \c0.tx.n14296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i2_4_lut_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__33767\,
            in1 => \N__30706\,
            in2 => \N__41467\,
            in3 => \N__30642\,
            lcout => n14442,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i2_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30644\,
            in1 => \N__33769\,
            in2 => \N__30721\,
            in3 => \N__41444\,
            lcout => \r_SM_Main_2_adj_4549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i3_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30844\,
            in1 => \N__41456\,
            in2 => \_gnd_net_\,
            in3 => \N__30826\,
            lcout => \c0.tx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1770_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__34301\,
            in1 => \N__52981\,
            in2 => \_gnd_net_\,
            in3 => \N__53194\,
            lcout => \c0.n21370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1597_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46176\,
            in2 => \_gnd_net_\,
            in3 => \N__42985\,
            lcout => \c0.n38_adj_4390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i1_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30898\,
            in1 => \N__41455\,
            in2 => \_gnd_net_\,
            in3 => \N__30880\,
            lcout => \c0.tx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i2_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41454\,
            in1 => \N__30871\,
            in2 => \_gnd_net_\,
            in3 => \N__30853\,
            lcout => \c0.tx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1776_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__37334\,
            in1 => \N__53181\,
            in2 => \_gnd_net_\,
            in3 => \N__53011\,
            lcout => \c0.n21376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1598_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110001"
        )
    port map (
            in0 => \N__31009\,
            in1 => \N__42834\,
            in2 => \N__46177\,
            in3 => \N__40471\,
            lcout => \c0.n4_adj_4391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i8_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34246\,
            in2 => \_gnd_net_\,
            in3 => \N__52870\,
            lcout => \c0.FRAME_MATCHER_state_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66826\,
            ce => 'H',
            sr => \N__34222\
        );

    \c0.FRAME_MATCHER_state_i17_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37847\,
            in2 => \_gnd_net_\,
            in3 => \N__52873\,
            lcout => \c0.FRAME_MATCHER_state_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66838\,
            ce => 'H',
            sr => \N__29233\
        );

    \c0.FRAME_MATCHER_state_i18_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37903\,
            in2 => \_gnd_net_\,
            in3 => \N__52874\,
            lcout => \c0.FRAME_MATCHER_state_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66849\,
            ce => 'H',
            sr => \N__37570\
        );

    \c0.i1_2_lut_3_lut_adj_1762_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__37876\,
            in1 => \N__53175\,
            in2 => \_gnd_net_\,
            in3 => \N__53027\,
            lcout => \c0.n21360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1759_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__34564\,
            in1 => \N__53197\,
            in2 => \_gnd_net_\,
            in3 => \N__53028\,
            lcout => \c0.n21356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1846_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31993\,
            in1 => \N__31434\,
            in2 => \N__29227\,
            in3 => \N__31570\,
            lcout => \c0.n12_adj_4516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1874_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__34454\,
            in1 => \N__29578\,
            in2 => \_gnd_net_\,
            in3 => \N__31070\,
            lcout => \c0.n9_adj_4339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1885_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__31404\,
            in1 => \N__29411\,
            in2 => \_gnd_net_\,
            in3 => \N__34452\,
            lcout => \c0.n22018\,
            ltout => \c0.n22018_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1398_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32204\,
            in1 => \N__29577\,
            in2 => \N__29380\,
            in3 => \N__30967\,
            lcout => \c0.n21946\,
            ltout => \c0.n21946_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1627_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29358\,
            in2 => \N__29362\,
            in3 => \N__29412\,
            lcout => \c0.n6_adj_4402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_3_lut_4_lut_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31688\,
            in1 => \N__34453\,
            in2 => \N__31351\,
            in3 => \N__31295\,
            lcout => \c0.n22188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1599_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31634\,
            in1 => \N__31341\,
            in2 => \N__31418\,
            in3 => \N__31297\,
            lcout => OPEN,
            ltout => \c0.n12491_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__6__5295_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29466\,
            in1 => \N__29359\,
            in2 => \N__29320\,
            in3 => \N__34362\,
            lcout => \c0.data_out_frame_28_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66644\,
            ce => \N__40950\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_6_i26_3_lut_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31777\,
            in1 => \N__29317\,
            in2 => \_gnd_net_\,
            in3 => \N__39836\,
            lcout => \c0.n26_adj_4351\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_adj_1608_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31296\,
            in1 => \N__31337\,
            in2 => \N__31219\,
            in3 => \N__31633\,
            lcout => OPEN,
            ltout => \c0.n7_adj_4307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1401_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31088\,
            in1 => \N__29271\,
            in2 => \N__29296\,
            in3 => \N__29529\,
            lcout => \data_out_frame_29__3__N_1662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__4__5289_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29530\,
            in1 => \N__29491\,
            in2 => \N__31102\,
            in3 => \N__29272\,
            lcout => \c0.data_out_frame_29_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66644\,
            ce => \N__40950\,
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1832_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__31405\,
            in1 => \N__31217\,
            in2 => \_gnd_net_\,
            in3 => \N__31071\,
            lcout => \c0.n22151\,
            ltout => \c0.n22151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__5__5288_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29485\,
            in3 => \N__29742\,
            lcout => \c0.data_out_frame_29_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66644\,
            ce => \N__40950\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1618_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__32380\,
            in1 => \N__31988\,
            in2 => \_gnd_net_\,
            in3 => \N__32932\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4397_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__0__5301_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__29728\,
            in1 => \N__32114\,
            in2 => \N__29482\,
            in3 => \N__29806\,
            lcout => \c0.data_out_frame_28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66651\,
            ce => \N__40954\,
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1825_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32113\,
            in1 => \N__32245\,
            in2 => \N__31838\,
            in3 => \N__29727\,
            lcout => \c0.n21876\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__5__5296_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__32211\,
            in1 => \_gnd_net_\,
            in2 => \N__29473\,
            in3 => \N__31462\,
            lcout => \c0.data_out_frame_28_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66651\,
            ce => \N__40954\,
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_5_i26_3_lut_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39837\,
            in1 => \N__29455\,
            in2 => \_gnd_net_\,
            in3 => \N__29449\,
            lcout => \c0.n26_adj_4347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1714_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29853\,
            in1 => \N__31208\,
            in2 => \_gnd_net_\,
            in3 => \N__29766\,
            lcout => \c0.n21210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1819_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__31656\,
            in1 => \N__29424\,
            in2 => \_gnd_net_\,
            in3 => \N__32248\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1820_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34928\,
            in1 => \N__29575\,
            in2 => \N__29611\,
            in3 => \N__34817\,
            lcout => \c0.n22393\,
            ltout => \c0.n22393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1822_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__29601\,
            in1 => \N__31218\,
            in2 => \N__29584\,
            in3 => \N__32014\,
            lcout => OPEN,
            ltout => \c0.n14_adj_4510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1823_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38295\,
            in1 => \N__31922\,
            in2 => \N__29581\,
            in3 => \N__29509\,
            lcout => \c0.n22346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1875_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__29576\,
            in1 => \N__34445\,
            in2 => \_gnd_net_\,
            in3 => \N__29520\,
            lcout => \c0.n10_adj_4511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1818_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__32733\,
            in1 => \N__53392\,
            in2 => \_gnd_net_\,
            in3 => \N__29824\,
            lcout => \c0.n22177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1865_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__29851\,
            in1 => \N__38966\,
            in2 => \N__32738\,
            in3 => \N__29780\,
            lcout => \c0.n20274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1424_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29850\,
            in2 => \_gnd_net_\,
            in3 => \N__29764\,
            lcout => \c0.n21192\,
            ltout => \c0.n21192_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1463_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__30082\,
            in1 => \N__29503\,
            in2 => \N__29497\,
            in3 => \N__38590\,
            lcout => \c0.n20931\,
            ltout => \c0.n20931_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1867_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__38967\,
            in1 => \N__32726\,
            in2 => \N__29494\,
            in3 => \N__29825\,
            lcout => \c0.n21283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1421_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__29852\,
            in1 => \_gnd_net_\,
            in2 => \N__29830\,
            in3 => \_gnd_net_\,
            lcout => \c0.n12554\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1868_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__29781\,
            in1 => \N__32725\,
            in2 => \N__38971\,
            in3 => \N__29765\,
            lcout => \c0.n21189\,
            ltout => \c0.n21189_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1802_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31377\,
            in2 => \N__29746\,
            in3 => \N__29743\,
            lcout => \c0.n20151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1878_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35213\,
            in1 => \N__32824\,
            in2 => \N__32302\,
            in3 => \N__29721\,
            lcout => \c0.n10513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1697_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38294\,
            in1 => \N__35116\,
            in2 => \N__32739\,
            in3 => \N__29706\,
            lcout => \c0.n10467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1742_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__29659\,
            in1 => \_gnd_net_\,
            in2 => \N__36460\,
            in3 => \N__35316\,
            lcout => \c0.n13480\,
            ltout => \c0.n13480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1737_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31877\,
            in2 => \N__29671\,
            in3 => \N__31956\,
            lcout => \c0.n21122\,
            ltout => \c0.n21122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1589_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32367\,
            in1 => \N__31882\,
            in2 => \N__29668\,
            in3 => \N__32420\,
            lcout => \c0.data_out_frame_29__7__N_1144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20421_2_lut_3_lut_4_lut_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31881\,
            in1 => \N__36458\,
            in2 => \N__35320\,
            in3 => \N__29660\,
            lcout => \c0.n24119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1426_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__30164\,
            in1 => \N__39292\,
            in2 => \_gnd_net_\,
            in3 => \N__39430\,
            lcout => \c0.n20767\,
            ltout => \c0.n20767_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1427_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29965\,
            in3 => \N__34627\,
            lcout => \c0.n21848\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1882_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31957\,
            in1 => \N__32493\,
            in2 => \_gnd_net_\,
            in3 => \N__32421\,
            lcout => \c0.n21112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1409_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__36165\,
            in1 => \N__33244\,
            in2 => \N__29957\,
            in3 => \N__38563\,
            lcout => \c0.n21943\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i10_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29914\,
            in1 => \N__38459\,
            in2 => \_gnd_net_\,
            in3 => \N__35209\,
            lcout => encoder1_position_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__6__5447_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__49332\,
            in1 => \N__49026\,
            in2 => \N__29902\,
            in3 => \N__36166\,
            lcout => data_out_frame_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__6__5415_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__49024\,
            in1 => \N__49333\,
            in2 => \N__34984\,
            in3 => \N__29883\,
            lcout => data_out_frame_13_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__4__5457_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__49331\,
            in1 => \N__49025\,
            in2 => \N__30232\,
            in3 => \N__38874\,
            lcout => data_out_frame_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i11_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29866\,
            in1 => \N__38460\,
            in2 => \_gnd_net_\,
            in3 => \N__32965\,
            lcout => encoder1_position_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_2_i11_3_lut_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39818\,
            in1 => \N__35002\,
            in2 => \_gnd_net_\,
            in3 => \N__35170\,
            lcout => \c0.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1462_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53388\,
            in1 => \N__35284\,
            in2 => \N__41605\,
            in3 => \N__39060\,
            lcout => \c0.n14_adj_4329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i7_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34907\,
            in1 => \N__30073\,
            in2 => \_gnd_net_\,
            in3 => \N__38465\,
            lcout => encoder1_position_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i13_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38461\,
            in1 => \N__30061\,
            in2 => \_gnd_net_\,
            in3 => \N__38046\,
            lcout => encoder1_position_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1690_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38247\,
            in1 => \N__35762\,
            in2 => \N__30030\,
            in3 => \N__48533\,
            lcout => \c0.n21855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i19_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30049\,
            in1 => \_gnd_net_\,
            in2 => \N__38496\,
            in3 => \N__30025\,
            lcout => encoder1_position_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__30004\,
            in1 => \N__35668\,
            in2 => \_gnd_net_\,
            in3 => \N__30238\,
            lcout => \c0.n23557\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i2_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42222\,
            in1 => \N__33112\,
            in2 => \_gnd_net_\,
            in3 => \N__53448\,
            lcout => encoder0_position_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i30_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48553\,
            in1 => \N__33325\,
            in2 => \_gnd_net_\,
            in3 => \N__42223\,
            lcout => encoder0_position_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i25_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38466\,
            in1 => \N__29992\,
            in2 => \_gnd_net_\,
            in3 => \N__33010\,
            lcout => encoder1_position_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i7_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__33199\,
            in1 => \_gnd_net_\,
            in2 => \N__42231\,
            in3 => \N__33249\,
            lcout => encoder0_position_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1441_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33230\,
            in2 => \_gnd_net_\,
            in3 => \N__41811\,
            lcout => OPEN,
            ltout => \c0.n21914_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1446_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53436\,
            in1 => \N__38167\,
            in2 => \N__30241\,
            in3 => \N__37061\,
            lcout => \c0.n21_adj_4320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i19_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42180\,
            in1 => \N__33286\,
            in2 => \_gnd_net_\,
            in3 => \N__38652\,
            lcout => encoder0_position_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20185_3_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39817\,
            in1 => \N__30192\,
            in2 => \_gnd_net_\,
            in3 => \N__30231\,
            lcout => \c0.n23880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__4__5449_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__39040\,
            in1 => \N__48946\,
            in2 => \N__30196\,
            in3 => \N__49402\,
            lcout => data_out_frame_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i27_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38506\,
            in1 => \N__30184\,
            in2 => \_gnd_net_\,
            in3 => \N__30163\,
            lcout => encoder1_position_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66728\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_10__2__5443_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49472\,
            in1 => \N__48887\,
            in2 => \N__35659\,
            in3 => \N__30129\,
            lcout => data_out_frame_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66728\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__4__5481_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__48886\,
            in1 => \N__49474\,
            in2 => \N__42403\,
            in3 => \N__30111\,
            lcout => data_out_frame_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66728\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__4__5473_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__49473\,
            in1 => \N__30384\,
            in2 => \N__38785\,
            in3 => \N__48888\,
            lcout => data_out_frame_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66728\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20139_4_lut_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30340\,
            in1 => \N__36381\,
            in2 => \N__36310\,
            in3 => \N__36594\,
            lcout => \c0.n23834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1691_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35997\,
            in1 => \N__36122\,
            in2 => \N__33243\,
            in3 => \N__41810\,
            lcout => \c0.n22449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i4_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30809\,
            in1 => \N__41486\,
            in2 => \_gnd_net_\,
            in3 => \N__30793\,
            lcout => \c0.tx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1536_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__30370\,
            in1 => \N__30299\,
            in2 => \N__36216\,
            in3 => \N__36646\,
            lcout => OPEN,
            ltout => \c0.n20_adj_4362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_1596_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30355\,
            in2 => \N__30349\,
            in3 => \N__30346\,
            lcout => \c0.n63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1702_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__36948\,
            in1 => \N__30339\,
            in2 => \N__30301\,
            in3 => \N__36587\,
            lcout => OPEN,
            ltout => \c0.n17_adj_4479_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1703_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__30277\,
            in1 => \N__36645\,
            in2 => \N__30259\,
            in3 => \N__36343\,
            lcout => \c0.n13006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1765_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__41893\,
            in1 => \N__36624\,
            in2 => \_gnd_net_\,
            in3 => \N__30478\,
            lcout => \c0.n13023\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i5_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30513\,
            in1 => \N__43269\,
            in2 => \_gnd_net_\,
            in3 => \N__41968\,
            lcout => data_in_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66755\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1695_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__30619\,
            in1 => \N__30592\,
            in2 => \N__35260\,
            in3 => \N__30579\,
            lcout => \c0.n17_adj_4477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Tx_Active_47_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__30568\,
            in1 => \N__37142\,
            in2 => \_gnd_net_\,
            in3 => \N__30720\,
            lcout => \c0.tx_active\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66755\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i10_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34164\,
            in1 => \_gnd_net_\,
            in2 => \N__43273\,
            in3 => \N__36324\,
            lcout => data_in_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66755\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i1_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__30526\,
            in1 => \_gnd_net_\,
            in2 => \N__30559\,
            in3 => \N__43268\,
            lcout => data_in_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66755\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1763_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__36323\,
            in1 => \N__30525\,
            in2 => \N__30514\,
            in3 => \N__30494\,
            lcout => \c0.n10_adj_4494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1699_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__34156\,
            in1 => \N__34197\,
            in2 => \N__30472\,
            in3 => \N__30460\,
            lcout => \c0.n117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1744_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__39264\,
            in1 => \N__37135\,
            in2 => \_gnd_net_\,
            in3 => \N__37171\,
            lcout => \c0.n44_adj_4336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1448020_i1_3_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__30454\,
            in1 => \N__30409\,
            in2 => \_gnd_net_\,
            in3 => \N__30400\,
            lcout => OPEN,
            ltout => \o_Tx_Serial_N_3783_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i26_3_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001010"
        )
    port map (
            in0 => \N__30704\,
            in1 => \_gnd_net_\,
            in2 => \N__30751\,
            in3 => \N__33763\,
            lcout => \c0.tx.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_SM_Main_i1_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__30650\,
            in1 => \N__30705\,
            in2 => \N__33772\,
            in3 => \N__41490\,
            lcout => \r_SM_Main_1_adj_4550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_1184_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33756\,
            in2 => \_gnd_net_\,
            in3 => \N__30703\,
            lcout => \c0.tx.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i7_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__31024\,
            in1 => \N__31047\,
            in2 => \N__41496\,
            in3 => \N__41382\,
            lcout => \r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66769\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41547\,
            in2 => \_gnd_net_\,
            in3 => \N__30778\,
            lcout => OPEN,
            ltout => \c0.tx.n6_adj_4214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4_4_lut_adj_1180_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41342\,
            in1 => \N__31043\,
            in2 => \N__30664\,
            in3 => \N__30958\,
            lcout => \c0.tx.n16630\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_4_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__41457\,
            in1 => \N__41343\,
            in2 => \N__30943\,
            in3 => \N__41548\,
            lcout => n8,
            ltout => \n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i5_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__30760\,
            in1 => \N__30781\,
            in2 => \N__30622\,
            in3 => \N__41458\,
            lcout => \r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i1_2_lut_adj_1186_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30816\,
            in2 => \_gnd_net_\,
            in3 => \N__30842\,
            lcout => OPEN,
            ltout => \c0.tx.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4_4_lut_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30934\,
            in1 => \N__30896\,
            in2 => \N__30961\,
            in3 => \N__30869\,
            lcout => \c0.tx.n31\,
            ltout => \c0.tx.n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i4_4_lut_adj_1185_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__31042\,
            in1 => \N__30779\,
            in2 => \N__30952\,
            in3 => \N__30949\,
            lcout => \c0.tx.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_2_lut_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__41374\,
            in1 => \N__30933\,
            in2 => \_gnd_net_\,
            in3 => \N__30901\,
            lcout => \c0.tx.n23960\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \c0.tx.n19540\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_3_lut_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__41377\,
            in1 => \N__30897\,
            in2 => \_gnd_net_\,
            in3 => \N__30874\,
            lcout => \c0.tx.n23961\,
            ltout => OPEN,
            carryin => \c0.tx.n19540\,
            carryout => \c0.tx.n19541\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_4_lut_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__41376\,
            in1 => \N__30870\,
            in2 => \_gnd_net_\,
            in3 => \N__30847\,
            lcout => \c0.tx.n23958\,
            ltout => OPEN,
            carryin => \c0.tx.n19541\,
            carryout => \c0.tx.n19542\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_5_lut_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__41378\,
            in1 => \N__30843\,
            in2 => \_gnd_net_\,
            in3 => \N__30820\,
            lcout => \c0.tx.n23963\,
            ltout => OPEN,
            carryin => \c0.tx.n19542\,
            carryout => \c0.tx.n19543\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_6_lut_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__41375\,
            in1 => \N__30817\,
            in2 => \_gnd_net_\,
            in3 => \N__30784\,
            lcout => \c0.tx.n23953\,
            ltout => OPEN,
            carryin => \c0.tx.n19543\,
            carryout => \c0.tx.n19544\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_7_lut_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30780\,
            in2 => \_gnd_net_\,
            in3 => \N__30754\,
            lcout => n316,
            ltout => OPEN,
            carryin => \c0.tx.n19544\,
            carryout => \c0.tx.n19545\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_8_lut_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__41373\,
            in1 => \N__41546\,
            in2 => \_gnd_net_\,
            in3 => \N__31051\,
            lcout => \c0.tx.n23987\,
            ltout => OPEN,
            carryin => \c0.tx.n19545\,
            carryout => \c0.tx.n19546\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_9_lut_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31048\,
            in2 => \_gnd_net_\,
            in3 => \N__31015\,
            lcout => n314,
            ltout => OPEN,
            carryin => \c0.tx.n19546\,
            carryout => \c0.tx.n19547\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.add_59_10_lut_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__41344\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31012\,
            lcout => n313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1585_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__68638\,
            in2 => \_gnd_net_\,
            in3 => \N__42643\,
            lcout => \c0.n12878\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i27_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34279\,
            in2 => \_gnd_net_\,
            in3 => \N__52869\,
            lcout => \c0.FRAME_MATCHER_state_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66814\,
            ce => 'H',
            sr => \N__34264\
        );

    \c0.FRAME_MATCHER_state_i9_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37545\,
            in2 => \_gnd_net_\,
            in3 => \N__52871\,
            lcout => \c0.FRAME_MATCHER_state_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66827\,
            ce => 'H',
            sr => \N__37582\
        );

    \c0.FRAME_MATCHER_state_i16_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37881\,
            in2 => \_gnd_net_\,
            in3 => \N__52872\,
            lcout => \c0.FRAME_MATCHER_state_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66839\,
            ce => 'H',
            sr => \N__31003\
        );

    \c0.FRAME_MATCHER_state_i14_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34565\,
            in2 => \_gnd_net_\,
            in3 => \N__52889\,
            lcout => \c0.FRAME_MATCHER_state_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66858\,
            ce => 'H',
            sr => \N__30988\
        );

    \c0.i2_2_lut_4_lut_adj_1879_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34387\,
            in1 => \N__31687\,
            in2 => \N__31416\,
            in3 => \N__30982\,
            lcout => \c0.n6_adj_4305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i64_4_lut_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111010001011"
        )
    port map (
            in0 => \N__31852\,
            in1 => \N__34386\,
            in2 => \N__31504\,
            in3 => \N__31969\,
            lcout => \c0.n21050\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1842_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32518\,
            in1 => \N__31468\,
            in2 => \N__31693\,
            in3 => \N__31989\,
            lcout => \c0.n20658\,
            ltout => \c0.n20658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1844_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31457\,
            in2 => \N__31441\,
            in3 => \N__32109\,
            lcout => \c0.n22166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1709_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34388\,
            in1 => \N__31707\,
            in2 => \N__31417\,
            in3 => \N__31635\,
            lcout => \c0.n21811\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1412_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31350\,
            in2 => \_gnd_net_\,
            in3 => \N__31294\,
            lcout => \c0.n21168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1410_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__31159\,
            in1 => \_gnd_net_\,
            in2 => \N__33064\,
            in3 => \N__31128\,
            lcout => \c0.n20298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1404_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31213\,
            in1 => \N__33060\,
            in2 => \_gnd_net_\,
            in3 => \N__31158\,
            lcout => \c0.n22736\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1487_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__31129\,
            in1 => \N__34455\,
            in2 => \_gnd_net_\,
            in3 => \N__32641\,
            lcout => \c0.n21135\,
            ltout => \c0.n21135_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1794_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31093\,
            in1 => \N__31072\,
            in2 => \N__31054\,
            in3 => \N__31565\,
            lcout => \c0.n23260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1790_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__31729\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31527\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__6__5287_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31537\,
            in1 => \N__31720\,
            in2 => \N__31801\,
            in3 => \N__31797\,
            lcout => \c0.data_out_frame_29_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66645\,
            ce => \N__40946\,
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1588_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31771\,
            in1 => \N__35605\,
            in2 => \N__32385\,
            in3 => \N__31536\,
            lcout => \c0.n21852\,
            ltout => \c0.n21852_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1827_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32323\,
            in1 => \N__31741\,
            in2 => \N__31732\,
            in3 => \N__31728\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1828_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31719\,
            in1 => \N__31708\,
            in2 => \N__31696\,
            in3 => \N__31515\,
            lcout => \c0.n20201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1488_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31692\,
            in2 => \_gnd_net_\,
            in3 => \N__31623\,
            lcout => OPEN,
            ltout => \c0.n21162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1816_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31582\,
            in1 => \N__31561\,
            in2 => \N__31540\,
            in3 => \N__32626\,
            lcout => \c0.n12526\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_29__7__5286_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__31528\,
            in1 => \_gnd_net_\,
            in2 => \N__31519\,
            in3 => \N__32561\,
            lcout => \c0.data_out_frame_29_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66645\,
            ce => \N__40946\,
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__7__5414_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__49322\,
            in1 => \N__32064\,
            in2 => \N__34933\,
            in3 => \N__48980\,
            lcout => data_out_frame_13_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1812_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32246\,
            in1 => \N__32002\,
            in2 => \N__32050\,
            in3 => \N__32013\,
            lcout => \c0.n20_adj_4505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1620_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33057\,
            in1 => \N__32446\,
            in2 => \_gnd_net_\,
            in3 => \N__32141\,
            lcout => \c0.n22072\,
            ltout => \c0.n22072_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1619_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31912\,
            in2 => \N__31996\,
            in3 => \N__32100\,
            lcout => \c0.n22073\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1647_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__33058\,
            in1 => \N__31894\,
            in2 => \N__32384\,
            in3 => \N__31968\,
            lcout => \c0.n20249\,
            ltout => \c0.n20249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1726_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32247\,
            in1 => \N__32554\,
            in2 => \N__31930\,
            in3 => \N__32512\,
            lcout => \c0.n12528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1395_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32373\,
            in2 => \_gnd_net_\,
            in3 => \N__31893\,
            lcout => \c0.n21842\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1850_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__32447\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33059\,
            lcout => \c0.n20230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1611_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34978\,
            in1 => \N__35134\,
            in2 => \N__32724\,
            in3 => \N__34927\,
            lcout => \c0.n6_adj_4394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1869_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__35135\,
            in1 => \N__38296\,
            in2 => \_gnd_net_\,
            in3 => \N__32704\,
            lcout => OPEN,
            ltout => \c0.n22163_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1813_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__34979\,
            in1 => \N__34857\,
            in2 => \N__32653\,
            in3 => \N__34792\,
            lcout => OPEN,
            ltout => \c0.n19_adj_4506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1815_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32572\,
            in1 => \N__32650\,
            in2 => \N__32644\,
            in3 => \N__32637\,
            lcout => \c0.n6_adj_4508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1814_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32616\,
            in1 => \N__32593\,
            in2 => \N__35064\,
            in3 => \N__33050\,
            lcout => \c0.n21_adj_4507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1881_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32553\,
            in1 => \N__32494\,
            in2 => \_gnd_net_\,
            in3 => \N__32442\,
            lcout => \c0.n21253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1851_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32372\,
            in2 => \_gnd_net_\,
            in3 => \N__32919\,
            lcout => \c0.n22078\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1877_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35208\,
            in1 => \N__32816\,
            in2 => \N__32309\,
            in3 => \N__32233\,
            lcout => \c0.n20180\,
            ltout => \c0.n20180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1890_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32186\,
            in1 => \N__33056\,
            in2 => \N__32152\,
            in3 => \N__32135\,
            lcout => \c0.n20465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1710_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35201\,
            in1 => \N__32918\,
            in2 => \N__33084\,
            in3 => \N__32852\,
            lcout => \c0.n21196\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1437_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35568\,
            in1 => \N__39488\,
            in2 => \N__33018\,
            in3 => \N__35401\,
            lcout => \c0.n20232\,
            ltout => \c0.n20232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1439_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__32955\,
            in1 => \_gnd_net_\,
            in2 => \N__32935\,
            in3 => \N__35590\,
            lcout => \c0.n21146\,
            ltout => \c0.n21146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1440_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32905\,
            in3 => \N__35200\,
            lcout => \c0.n22483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1417_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__32902\,
            in1 => \N__36058\,
            in2 => \N__38149\,
            in3 => \N__32845\,
            lcout => \c0.n20744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i27_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33366\,
            in1 => \N__42248\,
            in2 => \_gnd_net_\,
            in3 => \N__33343\,
            lcout => encoder0_position_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i1_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__33121\,
            in1 => \_gnd_net_\,
            in2 => \N__42252\,
            in3 => \N__35765\,
            lcout => encoder0_position_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__1__5420_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__49272\,
            in1 => \N__34731\,
            in2 => \N__32800\,
            in3 => \N__48895\,
            lcout => data_out_frame_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i20_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__33277\,
            in1 => \_gnd_net_\,
            in2 => \N__42253\,
            in3 => \N__36121\,
            lcout => encoder0_position_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i13_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33175\,
            in1 => \N__42240\,
            in2 => \_gnd_net_\,
            in3 => \N__35713\,
            lcout => encoder0_position_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i14_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__42241\,
            in1 => \_gnd_net_\,
            in2 => \N__35890\,
            in3 => \N__33310\,
            lcout => encoder0_position_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1862_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38257\,
            in1 => \N__35877\,
            in2 => \N__33376\,
            in3 => \N__35812\,
            lcout => \c0.n20160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_1_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33606\,
            in2 => \N__33679\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \quad_counter0.n19580\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_2_lut_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37046\,
            in2 => \N__33145\,
            in3 => \N__33124\,
            lcout => n2271,
            ltout => OPEN,
            carryin => \quad_counter0.n19580\,
            carryout => \quad_counter0.n19581\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_3_lut_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35764\,
            in2 => \N__33680\,
            in3 => \N__33115\,
            lcout => n2270,
            ltout => OPEN,
            carryin => \quad_counter0.n19581\,
            carryout => \quad_counter0.n19582\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_4_lut_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53457\,
            in2 => \N__33676\,
            in3 => \N__33106\,
            lcout => n2269,
            ltout => OPEN,
            carryin => \quad_counter0.n19582\,
            carryout => \quad_counter0.n19583\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_5_lut_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41696\,
            in2 => \N__33681\,
            in3 => \N__33091\,
            lcout => n2268,
            ltout => OPEN,
            carryin => \quad_counter0.n19583\,
            carryout => \quad_counter0.n19584\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_6_lut_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39036\,
            in2 => \N__33677\,
            in3 => \N__33088\,
            lcout => n2267,
            ltout => OPEN,
            carryin => \quad_counter0.n19584\,
            carryout => \quad_counter0.n19585\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_7_lut_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36062\,
            in2 => \N__33682\,
            in3 => \N__33259\,
            lcout => n2266,
            ltout => OPEN,
            carryin => \quad_counter0.n19585\,
            carryout => \quad_counter0.n19586\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_8_lut_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36159\,
            in2 => \N__33678\,
            in3 => \N__33256\,
            lcout => n2265,
            ltout => OPEN,
            carryin => \quad_counter0.n19586\,
            carryout => \quad_counter0.n19587\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_9_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33628\,
            in2 => \N__33245\,
            in3 => \N__33193\,
            lcout => n2264,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \quad_counter0.n19588\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_10_lut_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40305\,
            in2 => \N__33683\,
            in3 => \N__33190\,
            lcout => n2263,
            ltout => OPEN,
            carryin => \quad_counter0.n19588\,
            carryout => \quad_counter0.n19589\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_11_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33632\,
            in2 => \N__38723\,
            in3 => \N__33187\,
            lcout => n2262,
            ltout => OPEN,
            carryin => \quad_counter0.n19589\,
            carryout => \quad_counter0.n19590\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_12_lut_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39975\,
            in2 => \N__33684\,
            in3 => \N__33184\,
            lcout => n2261,
            ltout => OPEN,
            carryin => \quad_counter0.n19590\,
            carryout => \quad_counter0.n19591\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_13_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33636\,
            in2 => \N__39394\,
            in3 => \N__33181\,
            lcout => n2260,
            ltout => OPEN,
            carryin => \quad_counter0.n19591\,
            carryout => \quad_counter0.n19592\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_14_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38869\,
            in2 => \N__33685\,
            in3 => \N__33178\,
            lcout => n2259,
            ltout => OPEN,
            carryin => \quad_counter0.n19592\,
            carryout => \quad_counter0.n19593\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_15_lut_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33640\,
            in2 => \N__35724\,
            in3 => \N__33166\,
            lcout => n2258,
            ltout => OPEN,
            carryin => \quad_counter0.n19593\,
            carryout => \quad_counter0.n19594\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_16_lut_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35891\,
            in2 => \N__33686\,
            in3 => \N__33301\,
            lcout => n2257,
            ltout => OPEN,
            carryin => \quad_counter0.n19594\,
            carryout => \quad_counter0.n19595\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_17_lut_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36252\,
            in2 => \N__33691\,
            in3 => \N__33298\,
            lcout => n2256,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \quad_counter0.n19596\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_18_lut_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33663\,
            in2 => \N__39114\,
            in3 => \N__33295\,
            lcout => n2255,
            ltout => OPEN,
            carryin => \quad_counter0.n19596\,
            carryout => \quad_counter0.n19597\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_19_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33664\,
            in2 => \N__36556\,
            in3 => \N__33292\,
            lcout => n2254,
            ltout => OPEN,
            carryin => \quad_counter0.n19597\,
            carryout => \quad_counter0.n19598\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_20_lut_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41754\,
            in2 => \N__33692\,
            in3 => \N__33289\,
            lcout => n2253,
            ltout => OPEN,
            carryin => \quad_counter0.n19598\,
            carryout => \quad_counter0.n19599\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_21_lut_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33668\,
            in2 => \N__38662\,
            in3 => \N__33280\,
            lcout => n2252,
            ltout => OPEN,
            carryin => \quad_counter0.n19599\,
            carryout => \quad_counter0.n19600\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_22_lut_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36123\,
            in2 => \N__33693\,
            in3 => \N__33268\,
            lcout => n2251,
            ltout => OPEN,
            carryin => \quad_counter0.n19600\,
            carryout => \quad_counter0.n19601\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_23_lut_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33672\,
            in2 => \N__35993\,
            in3 => \N__33265\,
            lcout => n2250,
            ltout => OPEN,
            carryin => \quad_counter0.n19601\,
            carryout => \quad_counter0.n19602\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_24_lut_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42045\,
            in2 => \N__33694\,
            in3 => \N__33262\,
            lcout => n2249,
            ltout => OPEN,
            carryin => \quad_counter0.n19602\,
            carryout => \quad_counter0.n19603\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_25_lut_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33644\,
            in2 => \N__40366\,
            in3 => \N__33406\,
            lcout => n2248,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \quad_counter0.n19604\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_26_lut_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39320\,
            in2 => \N__33687\,
            in3 => \N__33403\,
            lcout => n2247,
            ltout => OPEN,
            carryin => \quad_counter0.n19604\,
            carryout => \quad_counter0.n19605\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_27_lut_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33648\,
            in2 => \N__39907\,
            in3 => \N__33400\,
            lcout => n2246,
            ltout => OPEN,
            carryin => \quad_counter0.n19605\,
            carryout => \quad_counter0.n19606\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_28_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40059\,
            in2 => \N__33688\,
            in3 => \N__33397\,
            lcout => n2245,
            ltout => OPEN,
            carryin => \quad_counter0.n19606\,
            carryout => \quad_counter0.n19607\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_29_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33652\,
            in2 => \N__33387\,
            in3 => \N__33334\,
            lcout => n2244,
            ltout => OPEN,
            carryin => \quad_counter0.n19607\,
            carryout => \quad_counter0.n19608\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_30_lut_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38784\,
            in2 => \N__33689\,
            in3 => \N__33331\,
            lcout => n2243,
            ltout => OPEN,
            carryin => \quad_counter0.n19608\,
            carryout => \quad_counter0.n19609\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_31_lut_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33656\,
            in2 => \N__38248\,
            in3 => \N__33328\,
            lcout => n2242,
            ltout => OPEN,
            carryin => \quad_counter0.n19609\,
            carryout => \quad_counter0.n19610\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_32_lut_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48551\,
            in2 => \N__33690\,
            in3 => \N__33313\,
            lcout => n2241,
            ltout => OPEN,
            carryin => \quad_counter0.n19610\,
            carryout => \quad_counter0.n19611\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.add_645_33_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41628\,
            in1 => \N__33605\,
            in2 => \_gnd_net_\,
            in3 => \N__33496\,
            lcout => n2240,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1390_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__37945\,
            in1 => \N__37468\,
            in2 => \_gnd_net_\,
            in3 => \N__37501\,
            lcout => OPEN,
            ltout => \c0.n14474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18960_4_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__37502\,
            in1 => \N__42506\,
            in2 => \N__33493\,
            in3 => \N__37409\,
            lcout => \c0.n22651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__1__5452_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49450\,
            in1 => \N__48743\,
            in2 => \N__35776\,
            in3 => \N__33490\,
            lcout => data_out_frame_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.n24183_bdd_4_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__33489\,
            in1 => \N__36652\,
            in2 => \N__33481\,
            in3 => \N__36890\,
            lcout => \c0.n24186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i23_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42106\,
            in1 => \N__33448\,
            in2 => \_gnd_net_\,
            in3 => \N__40355\,
            lcout => encoder0_position_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i31_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__42107\,
            in1 => \N__33442\,
            in2 => \N__41645\,
            in3 => \_gnd_net_\,
            lcout => encoder0_position_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__7__5462_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49449\,
            in1 => \N__48742\,
            in2 => \N__40367\,
            in3 => \N__33432\,
            lcout => data_out_frame_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__1__5484_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__48737\,
            in1 => \N__49455\,
            in2 => \N__33418\,
            in3 => \N__41870\,
            lcout => data_out_frame_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20396_3_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__33944\,
            in1 => \N__33414\,
            in2 => \_gnd_net_\,
            in3 => \N__39815\,
            lcout => \c0.n24093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1204_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44929\,
            in2 => \_gnd_net_\,
            in3 => \N__59353\,
            lcout => \c0.n22358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__1__5468_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__49453\,
            in1 => \N__48739\,
            in2 => \N__34009\,
            in3 => \N__36559\,
            lcout => data_out_frame_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_5__7__5478_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__48738\,
            in1 => \N__49456\,
            in2 => \N__42352\,
            in3 => \N__33804\,
            lcout => data_out_frame_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__0__5461_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49454\,
            in1 => \N__48740\,
            in2 => \N__40312\,
            in3 => \N__34023\,
            lcout => data_out_frame_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66756\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_1_i5_3_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39816\,
            in1 => \N__34005\,
            in2 => \_gnd_net_\,
            in3 => \N__37083\,
            lcout => OPEN,
            ltout => \c0.n5_adj_4518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20167_4_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__33945\,
            in1 => \N__33997\,
            in2 => \N__33991\,
            in3 => \N__36909\,
            lcout => \c0.n23862\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1682_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__68570\,
            in1 => \N__46148\,
            in2 => \_gnd_net_\,
            in3 => \N__42639\,
            lcout => \c0.n20_adj_4327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20358_3_lut_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__39814\,
            in1 => \N__33943\,
            in2 => \_gnd_net_\,
            in3 => \N__33805\,
            lcout => \c0.n24054\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.i3737_2_lut_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33770\,
            in2 => \_gnd_net_\,
            in3 => \N__39269\,
            lcout => \c0.tx.n7086\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1389_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__37469\,
            in1 => \N__37424\,
            in2 => \_gnd_net_\,
            in3 => \N__37494\,
            lcout => \c0.n9668\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1900_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__37495\,
            in1 => \N__37389\,
            in2 => \N__37432\,
            in3 => \N__37470\,
            lcout => \data_out_frame_29_7_N_1483_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i12_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43263\,
            in1 => \N__34198\,
            in2 => \_gnd_net_\,
            in3 => \N__36367\,
            lcout => data_in_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66770\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i18_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43264\,
            in1 => \N__34157\,
            in2 => \_gnd_net_\,
            in3 => \N__43043\,
            lcout => data_in_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66770\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1872_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34542\,
            in1 => \N__34129\,
            in2 => \N__41155\,
            in3 => \N__34036\,
            lcout => \c0.n13_adj_4388\,
            ltout => \c0.n13_adj_4388_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1887_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__37819\,
            in1 => \_gnd_net_\,
            in2 => \N__34132\,
            in3 => \N__37620\,
            lcout => \c0.n21789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1393_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43539\,
            in1 => \N__34308\,
            in2 => \N__37335\,
            in3 => \N__37753\,
            lcout => \c0.n23135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i11_4_lut_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34123\,
            in1 => \N__34105\,
            in2 => \N__34087\,
            in3 => \N__34066\,
            lcout => \quad_counter0.n27_adj_4200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1358_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34277\,
            in2 => \_gnd_net_\,
            in3 => \N__34503\,
            lcout => \c0.n14457\,
            ltout => \c0.n14457_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_adj_1645_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34309\,
            in1 => \N__41053\,
            in2 => \N__34282\,
            in3 => \N__41007\,
            lcout => \c0.n49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1774_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__37609\,
            in1 => \N__53193\,
            in2 => \_gnd_net_\,
            in3 => \N__52947\,
            lcout => \c0.n21372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1522_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34278\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40652\,
            lcout => \c0.n21330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1526_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40653\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34504\,
            lcout => \c0.n21326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1635_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37914\,
            in2 => \_gnd_net_\,
            in3 => \N__43455\,
            lcout => OPEN,
            ltout => \c0.n30_adj_4411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i22_4_lut_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41151\,
            in1 => \N__34576\,
            in2 => \N__34252\,
            in3 => \N__34248\,
            lcout => \c0.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1751_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__52974\,
            in1 => \N__34249\,
            in2 => \_gnd_net_\,
            in3 => \N__53170\,
            lcout => \c0.n21344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1778_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__53169\,
            in1 => \N__42547\,
            in2 => \N__37803\,
            in3 => \N__42767\,
            lcout => \c0.n21336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1746_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__42766\,
            in1 => \N__42870\,
            in2 => \_gnd_net_\,
            in3 => \N__40633\,
            lcout => \c0.n4_adj_4345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i25_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37752\,
            in2 => \_gnd_net_\,
            in3 => \N__52860\,
            lcout => \c0.FRAME_MATCHER_state_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66815\,
            ce => 'H',
            sr => \N__37726\
        );

    \c0.i16_4_lut_adj_1636_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34567\,
            in1 => \N__37750\,
            in2 => \N__34543\,
            in3 => \N__37880\,
            lcout => \c0.n44_adj_4412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1768_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__53189\,
            in1 => \N__34540\,
            in2 => \_gnd_net_\,
            in3 => \N__53009\,
            lcout => \c0.n21368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1891_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37541\,
            in1 => \N__37716\,
            in2 => \N__42936\,
            in3 => \N__34566\,
            lcout => \c0.n19_adj_4481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i21_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34541\,
            in2 => \_gnd_net_\,
            in3 => \N__52885\,
            lcout => \c0.FRAME_MATCHER_state_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66840\,
            ce => 'H',
            sr => \N__34516\
        );

    \c0.FRAME_MATCHER_state_i29_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34502\,
            in2 => \_gnd_net_\,
            in3 => \N__52887\,
            lcout => \c0.FRAME_MATCHER_state_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66850\,
            ce => 'H',
            sr => \N__34486\
        );

    \c0.i6_4_lut_adj_1623_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52183\,
            in1 => \N__54685\,
            in2 => \N__61072\,
            in3 => \N__48241\,
            lcout => \c0.n14_adj_4400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1795_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34477\,
            in1 => \N__34456\,
            in2 => \N__34398\,
            in3 => \N__34366\,
            lcout => OPEN,
            ltout => \c0.n16_adj_4498_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_28__7__5294_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34343\,
            in1 => \N__34318\,
            in2 => \N__34312\,
            in3 => \N__34774\,
            lcout => \c0.data_out_frame_28_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66639\,
            ce => \N__40945\,
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1796_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__34861\,
            in1 => \N__34834\,
            in2 => \N__34827\,
            in3 => \N__34801\,
            lcout => \c0.n17_adj_4499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_7_i26_3_lut_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39734\,
            in1 => \N__34768\,
            in2 => \_gnd_net_\,
            in3 => \N__34759\,
            lcout => \c0.n26_adj_4359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_1_i11_3_lut_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34735\,
            in1 => \N__34717\,
            in2 => \_gnd_net_\,
            in3 => \N__39733\,
            lcout => \c0.n11_adj_4520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1543_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__50350\,
            in1 => \N__44165\,
            in2 => \N__47523\,
            in3 => \N__51712\,
            lcout => \c0.n14_adj_4364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i30_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__67214\,
            in1 => \N__43216\,
            in2 => \_gnd_net_\,
            in3 => \N__35245\,
            lcout => data_in_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__3__5458_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__49255\,
            in1 => \N__34668\,
            in2 => \N__39391\,
            in3 => \N__48949\,
            lcout => data_out_frame_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_4_i11_3_lut_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39732\,
            in1 => \N__35080\,
            in2 => \_gnd_net_\,
            in3 => \N__34584\,
            lcout => \c0.n11_adj_4303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__4__5425_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__49254\,
            in1 => \N__48947\,
            in2 => \N__34588\,
            in3 => \N__34636\,
            lcout => data_out_frame_12_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__0__5429_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__49253\,
            in1 => \N__35334\,
            in2 => \N__35395\,
            in3 => \N__48948\,
            lcout => data_out_frame_12_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1456_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__34925\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35308\,
            lcout => \c0.n22174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i22_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35252\,
            in1 => \N__43175\,
            in2 => \_gnd_net_\,
            in3 => \N__36406\,
            lcout => data_in_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__2__5427_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__49269\,
            in1 => \N__49045\,
            in2 => \N__35169\,
            in3 => \N__35221\,
            lcout => data_out_frame_12_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1657_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40057\,
            in1 => \N__39903\,
            in2 => \N__39390\,
            in3 => \N__42351\,
            lcout => \c0.n21918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1476_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40304\,
            in2 => \_gnd_net_\,
            in3 => \N__40369\,
            lcout => \c0.n22474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__4__5417_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__49044\,
            in1 => \N__49271\,
            in2 => \N__35140\,
            in3 => \N__35079\,
            lcout => data_out_frame_13_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_13__2__5419_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49270\,
            in1 => \N__49046\,
            in2 => \N__35065\,
            in3 => \N__34998\,
            lcout => data_out_frame_13_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1418_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34980\,
            in2 => \_gnd_net_\,
            in3 => \N__34926\,
            lcout => \c0.n21896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1438_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39426\,
            in1 => \N__40261\,
            in2 => \N__35655\,
            in3 => \N__42046\,
            lcout => \c0.n20236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1447_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35431\,
            in1 => \N__35572\,
            in2 => \N__35545\,
            in3 => \N__35536\,
            lcout => OPEN,
            ltout => \c0.n16_adj_4321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_adj_1448_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35529\,
            in2 => \N__35479\,
            in3 => \N__38059\,
            lcout => OPEN,
            ltout => \c0.n18_adj_4322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1450_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53502\,
            in1 => \N__38905\,
            in2 => \N__35476\,
            in3 => \N__35473\,
            lcout => \c0.n14_adj_4324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1826_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38677\,
            in1 => \N__37263\,
            in2 => \N__36557\,
            in3 => \N__35928\,
            lcout => \c0.n22376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1465_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35701\,
            in2 => \_gnd_net_\,
            in3 => \N__35872\,
            lcout => \c0.n13619\,
            ltout => \c0.n13619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1467_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38676\,
            in1 => \N__38242\,
            in2 => \N__35425\,
            in3 => \N__53409\,
            lcout => \c0.n10_adj_4331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1431_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36549\,
            in2 => \_gnd_net_\,
            in3 => \N__38667\,
            lcout => OPEN,
            ltout => \c0.n13524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1436_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35422\,
            in1 => \N__38821\,
            in2 => \N__35404\,
            in3 => \N__35824\,
            lcout => \c0.n10_adj_4317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1906_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38243\,
            in1 => \N__38783\,
            in2 => \N__48570\,
            in3 => \N__35810\,
            lcout => \c0.n20328\,
            ltout => \c0.n20328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1692_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__35873\,
            in1 => \_gnd_net_\,
            in2 => \N__35842\,
            in3 => \N__35702\,
            lcout => \c0.n22367\,
            ltout => \c0.n22367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1435_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38599\,
            in1 => \N__36027\,
            in2 => \N__35827\,
            in3 => \N__36258\,
            lcout => \c0.n23569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1443_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39014\,
            in2 => \_gnd_net_\,
            in3 => \N__36056\,
            lcout => \c0.n22230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1442_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__36154\,
            in1 => \N__35979\,
            in2 => \_gnd_net_\,
            in3 => \N__42396\,
            lcout => \c0.n22382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i0_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42249\,
            in1 => \N__35818\,
            in2 => \_gnd_net_\,
            in3 => \N__37047\,
            lcout => encoder0_position_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_3_lut_4_lut_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48552\,
            in2 => \_gnd_net_\,
            in3 => \N__35811\,
            lcout => OPEN,
            ltout => \c0.n22461_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1444_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__35787\,
            in1 => \N__35763\,
            in2 => \N__35728\,
            in3 => \N__35703\,
            lcout => \c0.n20_adj_4318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i6_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36155\,
            in1 => \N__42251\,
            in2 => \_gnd_net_\,
            in3 => \N__36172\,
            lcout => encoder0_position_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1472_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36111\,
            in2 => \_gnd_net_\,
            in3 => \N__41799\,
            lcout => \c0.n21970\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i5_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36057\,
            in1 => \N__42250\,
            in2 => \_gnd_net_\,
            in3 => \N__36088\,
            lcout => encoder0_position_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66675\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1688_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41648\,
            in1 => \N__38756\,
            in2 => \N__48566\,
            in3 => \N__39091\,
            lcout => \c0.n21808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i21_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35989\,
            in1 => \N__36010\,
            in2 => \_gnd_net_\,
            in3 => \N__42208\,
            lcout => encoder0_position_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i9_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42209\,
            in1 => \N__35953\,
            in2 => \_gnd_net_\,
            in3 => \N__38722\,
            lcout => encoder0_position_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i11_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__35947\,
            in1 => \N__42204\,
            in2 => \N__39393\,
            in3 => \_gnd_net_\,
            lcout => encoder0_position_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i17_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__35938\,
            in1 => \_gnd_net_\,
            in2 => \N__42239\,
            in3 => \N__36531\,
            lcout => encoder0_position_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1479_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41649\,
            lcout => \c0.n10394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1640_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41647\,
            in1 => \N__44607\,
            in2 => \N__36257\,
            in3 => \N__36530\,
            lcout => \c0.n22248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1711_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39288\,
            in1 => \N__36499\,
            in2 => \N__39392\,
            in3 => \N__39403\,
            lcout => \c0.n13338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i182_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__59168\,
            in1 => \N__67201\,
            in2 => \_gnd_net_\,
            in3 => \N__63455\,
            lcout => data_in_frame_22_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1701_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36196\,
            in1 => \N__36299\,
            in2 => \N__36425\,
            in3 => \N__36377\,
            lcout => \c0.n16_adj_4478\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i2_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36300\,
            in1 => \N__43217\,
            in2 => \_gnd_net_\,
            in3 => \N__36331\,
            lcout => data_in_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__5__5472_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49570\,
            in1 => \N__48833\,
            in2 => \N__38245\,
            in3 => \N__36285\,
            lcout => data_out_frame_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i15_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42168\,
            in1 => \N__36271\,
            in2 => \_gnd_net_\,
            in3 => \N__36256\,
            lcout => encoder0_position_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i17_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36197\,
            in1 => \N__43218\,
            in2 => \_gnd_net_\,
            in3 => \N__40243\,
            lcout => data_in_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i24_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__36178\,
            in1 => \_gnd_net_\,
            in2 => \N__42221\,
            in3 => \N__39324\,
            lcout => encoder0_position_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i31_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__43243\,
            in1 => \_gnd_net_\,
            in2 => \N__65591\,
            in3 => \N__36985\,
            lcout => data_in_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i226_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__64561\,
            in1 => \N__63853\,
            in2 => \N__49962\,
            in3 => \N__67672\,
            lcout => \c0.data_in_frame_28_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i29_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42167\,
            in1 => \N__37000\,
            in2 => \_gnd_net_\,
            in3 => \N__38221\,
            lcout => encoder0_position_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i32_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__68974\,
            in1 => \N__43245\,
            in2 => \_gnd_net_\,
            in3 => \N__36643\,
            lcout => data_in_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i23_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43239\,
            in1 => \N__36986\,
            in2 => \_gnd_net_\,
            in3 => \N__36947\,
            lcout => data_in_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_0__bdd_4_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__36928\,
            in1 => \N__36818\,
            in2 => \N__37222\,
            in3 => \N__39726\,
            lcout => \c0.n24183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i24_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__36644\,
            in1 => \_gnd_net_\,
            in2 => \N__43265\,
            in3 => \N__36623\,
            lcout => data_in_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i27_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36586\,
            in1 => \N__43244\,
            in2 => \_gnd_net_\,
            in3 => \N__68377\,
            lcout => data_in_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66715\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__56934\,
            in1 => \N__57027\,
            in2 => \_gnd_net_\,
            in3 => \N__56836\,
            lcout => \c0.rx.n21783\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_11__1__5436_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__37221\,
            in1 => \N__48741\,
            in2 => \N__37264\,
            in3 => \N__49427\,
            lcout => data_out_frame_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_3_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__49425\,
            in1 => \N__39138\,
            in2 => \_gnd_net_\,
            in3 => \N__40150\,
            lcout => OPEN,
            ltout => \c0.n9_adj_4415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1748_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40734\,
            in2 => \N__37207\,
            in3 => \N__40775\,
            lcout => n14252,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20381_3_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__37170\,
            in1 => \_gnd_net_\,
            in2 => \N__37146\,
            in3 => \N__39248\,
            lcout => \c0.n23965\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1494_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37111\,
            in1 => \N__40149\,
            in2 => \N__40744\,
            in3 => \N__37360\,
            lcout => n22661,
            ltout => \n22661_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__3__5466_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__37098\,
            in1 => \N__49426\,
            in2 => \N__37105\,
            in3 => \N__38666\,
            lcout => data_out_frame_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1263_2_lut_3_lut_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__40445\,
            in1 => \N__40595\,
            in2 => \_gnd_net_\,
            in3 => \N__42705\,
            lcout => \c0.n3239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__1__5476_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49443\,
            in1 => \N__48736\,
            in2 => \N__39902\,
            in3 => \N__37084\,
            lcout => data_out_frame_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66743\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_9__0__5453_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__48735\,
            in1 => \N__49444\,
            in2 => \N__37071\,
            in3 => \N__37014\,
            lcout => data_out_frame_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66743\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1234_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111111"
        )
    port map (
            in0 => \N__42704\,
            in1 => \N__40446\,
            in2 => \N__42507\,
            in3 => \N__40113\,
            lcout => \c0.n12967\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1698_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__37297\,
            in1 => \N__37940\,
            in2 => \_gnd_net_\,
            in3 => \N__42703\,
            lcout => \c0.n12996\,
            ltout => \c0.n12996_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__42706\,
            in1 => \N__42502\,
            in2 => \N__37288\,
            in3 => \N__40114\,
            lcout => \c0.n13020\,
            ltout => \c0.n13020_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1677_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110101"
        )
    port map (
            in0 => \N__40447\,
            in1 => \N__40596\,
            in2 => \N__37285\,
            in3 => \N__42707\,
            lcout => \c0.n13021\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i0_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__50107\,
            in1 => \N__69375\,
            in2 => \N__59690\,
            in3 => \N__59940\,
            lcout => rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66743\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100110011"
        )
    port map (
            in0 => \N__37473\,
            in1 => \N__37428\,
            in2 => \N__37519\,
            in3 => \N__40402\,
            lcout => \c0.data_out_frame_29_7_N_1483_1\,
            ltout => \c0.data_out_frame_29_7_N_1483_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1678_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001111"
        )
    port map (
            in0 => \N__37430\,
            in1 => \_gnd_net_\,
            in2 => \N__37282\,
            in3 => \N__37279\,
            lcout => \c0.n4_adj_4419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i157_4_lut_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101010101"
        )
    port map (
            in0 => \N__37472\,
            in1 => \N__42498\,
            in2 => \N__37390\,
            in3 => \N__37514\,
            lcout => \c0.n6650\,
            ltout => \c0.n6650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1331_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__37429\,
            in1 => \N__37270\,
            in2 => \N__37273\,
            in3 => \N__37356\,
            lcout => \c0.n31_adj_4271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_adj_1783_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__37471\,
            in1 => \N__40401\,
            in2 => \N__37944\,
            in3 => \N__37513\,
            lcout => \c0.n6_adj_4270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1696_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__37515\,
            in1 => \N__37388\,
            in2 => \_gnd_net_\,
            in3 => \N__37474\,
            lcout => OPEN,
            ltout => \c0.n16958_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1491_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37345\,
            in2 => \N__37435\,
            in3 => \N__37431\,
            lcout => OPEN,
            ltout => \c0.n22695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i2_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__42568\,
            in1 => \N__42589\,
            in2 => \N__37393\,
            in3 => \N__40090\,
            lcout => \c0.FRAME_MATCHER_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66757\,
            ce => 'H',
            sr => \N__40934\
        );

    \c0.i14419_2_lut_4_lut_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__37818\,
            in1 => \N__37621\,
            in2 => \N__37372\,
            in3 => \N__42708\,
            lcout => \c0.n9207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1658_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__40575\,
            in1 => \N__40527\,
            in2 => \_gnd_net_\,
            in3 => \N__42709\,
            lcout => \c0.n12990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1490_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__42954\,
            in1 => \N__40419\,
            in2 => \N__42433\,
            in3 => \N__43340\,
            lcout => \c0.n14_adj_4337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_adj_1671_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__40745\,
            in1 => \N__40702\,
            in2 => \_gnd_net_\,
            in3 => \N__42710\,
            lcout => OPEN,
            ltout => \c0.n7_adj_4352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1533_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__54093\,
            in1 => \N__43341\,
            in2 => \N__37339\,
            in3 => \N__43291\,
            lcout => \c0.n6_adj_4353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_adj_1637_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38109\,
            in1 => \N__42937\,
            in2 => \N__52663\,
            in3 => \N__37336\,
            lcout => OPEN,
            ltout => \c0.n48_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_4_lut_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37525\,
            in1 => \N__37762\,
            in2 => \N__37663\,
            in3 => \N__37660\,
            lcout => \c0.n54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_1639_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37604\,
            in1 => \N__37653\,
            in2 => \N__41104\,
            in3 => \N__43540\,
            lcout => \c0.n45_adj_4413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1434_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43503\,
            in1 => \N__52659\,
            in2 => \N__37654\,
            in3 => \N__37603\,
            lcout => \c0.n14_adj_4316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i24_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37605\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52815\,
            lcout => \c0.FRAME_MATCHER_state_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66784\,
            ce => 'H',
            sr => \N__37588\
        );

    \c0.i14273_2_lut_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40599\,
            in2 => \_gnd_net_\,
            in3 => \N__42768\,
            lcout => \c0.data_out_frame_29_7_N_1483_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1781_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__42769\,
            in1 => \N__37686\,
            in2 => \N__53168\,
            in3 => \N__42546\,
            lcout => \c0.n21342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1752_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__52970\,
            in1 => \_gnd_net_\,
            in2 => \N__37555\,
            in3 => \N__53116\,
            lcout => \c0.n21346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1766_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__53115\,
            in1 => \_gnd_net_\,
            in2 => \N__37918\,
            in3 => \N__52971\,
            lcout => \c0.n21364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18_4_lut_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43504\,
            in1 => \N__37852\,
            in2 => \N__42508\,
            in3 => \N__37551\,
            lcout => \c0.n46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1704_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37685\,
            in1 => \N__38108\,
            in2 => \N__43456\,
            in3 => \N__41100\,
            lcout => OPEN,
            ltout => \c0.n21_adj_4480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_3_lut_adj_1716_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37969\,
            in2 => \N__37957\,
            in3 => \N__37954\,
            lcout => \c0.n14789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1871_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37913\,
            in1 => \N__41041\,
            in2 => \N__37885\,
            in3 => \N__37848\,
            lcout => \c0.n21682\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_1638_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37714\,
            in1 => \N__37687\,
            in2 => \N__43410\,
            in3 => \N__37804\,
            lcout => \c0.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1775_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__37751\,
            in1 => \N__53136\,
            in2 => \_gnd_net_\,
            in3 => \N__52973\,
            lcout => \c0.n21374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1753_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__53137\,
            in1 => \N__37715\,
            in2 => \_gnd_net_\,
            in3 => \N__52972\,
            lcout => \c0.n21348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i10_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37717\,
            in2 => \_gnd_net_\,
            in3 => \N__52859\,
            lcout => \c0.FRAME_MATCHER_state_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66816\,
            ce => 'H',
            sr => \N__37693\
        );

    \c0.FRAME_MATCHER_state_i7_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37684\,
            in2 => \_gnd_net_\,
            in3 => \N__52884\,
            lcout => \c0.FRAME_MATCHER_state_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66828\,
            ce => 'H',
            sr => \N__38119\
        );

    \c0.i1_2_lut_3_lut_adj_1755_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__38110\,
            in1 => \N__53010\,
            in2 => \_gnd_net_\,
            in3 => \N__53176\,
            lcout => \c0.n21350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i11_LC_15_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38107\,
            in2 => \_gnd_net_\,
            in3 => \N__52888\,
            lcout => \c0.FRAME_MATCHER_state_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66859\,
            ce => 'H',
            sr => \N__38083\
        );

    \c0.i14074_2_lut_3_lut_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__56699\,
            in1 => \N__56573\,
            in2 => \_gnd_net_\,
            in3 => \N__56434\,
            lcout => \c0.n17596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_12__5__5424_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49144\,
            in1 => \N__49048\,
            in2 => \N__38071\,
            in3 => \N__38007\,
            lcout => data_out_frame_12_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66634\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1648_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__56589\,
            in1 => \N__56435\,
            in2 => \_gnd_net_\,
            in3 => \N__46030\,
            lcout => \c0.n4_adj_4373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1626_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47908\,
            in2 => \_gnd_net_\,
            in3 => \N__47956\,
            lcout => \c0.n20875\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1545_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51777\,
            in1 => \N__43870\,
            in2 => \N__48171\,
            in3 => \N__43919\,
            lcout => \c0.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1544_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50345\,
            in1 => \N__51778\,
            in2 => \N__47522\,
            in3 => \N__51711\,
            lcout => \c0.n14_adj_4365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1546_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43871\,
            in1 => \N__44167\,
            in2 => \N__48172\,
            in3 => \N__43920\,
            lcout => OPEN,
            ltout => \c0.n13_adj_4366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14078_4_lut_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110000"
        )
    port map (
            in0 => \N__37993\,
            in1 => \N__37984\,
            in2 => \N__37978\,
            in3 => \N__37975\,
            lcout => \c0.n17600\,
            ltout => \c0.n17600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1624_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47266\,
            in1 => \N__38137\,
            in2 => \N__38131\,
            in3 => \N__54832\,
            lcout => \c0.n23648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i6_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41083\,
            in2 => \_gnd_net_\,
            in3 => \N__52886\,
            lcout => \c0.FRAME_MATCHER_state_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66643\,
            ce => 'H',
            sr => \N__41065\
        );

    \c0.i8_4_lut_adj_1629_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111101"
        )
    port map (
            in0 => \N__54767\,
            in1 => \N__41215\,
            in2 => \N__44257\,
            in3 => \N__43990\,
            lcout => \c0.n18_adj_4403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1306_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52391\,
            in2 => \_gnd_net_\,
            in3 => \N__54766\,
            lcout => \c0.n21825\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1307_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38127\,
            in1 => \N__47930\,
            in2 => \N__48317\,
            in3 => \N__48255\,
            lcout => \c0.n13677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i85_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__62493\,
            in1 => \N__69211\,
            in2 => \N__63217\,
            in3 => \N__38128\,
            lcout => \c0.data_in_frame_10_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i67_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__65970\,
            in1 => \N__62494\,
            in2 => \N__47937\,
            in3 => \N__68416\,
            lcout => \c0.data_in_frame_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i68_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62491\,
            in1 => \N__65972\,
            in2 => \N__48321\,
            in3 => \N__64851\,
            lcout => \c0.data_in_frame_8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1665_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__56601\,
            in1 => \N__56456\,
            in2 => \N__56742\,
            in3 => \N__68097\,
            lcout => n21760,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i69_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__62492\,
            in1 => \N__65973\,
            in2 => \N__63216\,
            in3 => \N__47450\,
            lcout => \c0.data_in_frame_8_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i78_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__67215\,
            in1 => \N__62495\,
            in2 => \N__69876\,
            in3 => \N__47823\,
            lcout => \c0.data_in_frame_9_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i66_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62490\,
            in1 => \N__65971\,
            in2 => \N__52407\,
            in3 => \N__63865\,
            lcout => \c0.data_in_frame_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1475_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40058\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39898\,
            lcout => \c0.n21908\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter1.count_i0_i20_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38504\,
            in1 => \N__38311\,
            in2 => \_gnd_net_\,
            in3 => \N__38914\,
            lcout => encoder1_position_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1419_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41601\,
            in1 => \N__41869\,
            in2 => \N__38887\,
            in3 => \N__39101\,
            lcout => \c0.n13839\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1468_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48562\,
            in2 => \_gnd_net_\,
            in3 => \N__38772\,
            lcout => \c0.n22015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.encoder0_position_29__I_0_2_lut_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__38773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38244\,
            lcout => \c0.data_out_frame_29__7__N_856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1416_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__38163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38610\,
            lcout => \c0.n6_adj_4311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1481_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38986\,
            in1 => \N__38556\,
            in2 => \N__38611\,
            in3 => \N__38809\,
            lcout => \c0.n22427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1843_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39476\,
            in1 => \N__41862\,
            in2 => \N__38668\,
            in3 => \N__41800\,
            lcout => \c0.n21885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_1177_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59884\,
            in2 => \_gnd_net_\,
            in3 => \N__57109\,
            lcout => n18678,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1473_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42034\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42395\,
            lcout => \c0.n22200\,
            ltout => \c0.n22200_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1848_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40208\,
            in1 => \N__39477\,
            in2 => \N__38593\,
            in3 => \N__38579\,
            lcout => \c0.n13705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1908_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48450\,
            in1 => \N__47454\,
            in2 => \_gnd_net_\,
            in3 => \N__47254\,
            lcout => \c0.n13190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i12_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42235\,
            in1 => \N__38545\,
            in2 => \_gnd_net_\,
            in3 => \N__38859\,
            lcout => encoder0_position_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i4_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39016\,
            in1 => \N__42237\,
            in2 => \_gnd_net_\,
            in3 => \N__38536\,
            lcout => encoder0_position_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i10_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42234\,
            in1 => \N__38524\,
            in2 => \_gnd_net_\,
            in3 => \N__39974\,
            lcout => encoder0_position_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i16_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39090\,
            in1 => \N__42236\,
            in2 => \_gnd_net_\,
            in3 => \N__39127\,
            lcout => encoder0_position_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1474_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41722\,
            in1 => \N__39089\,
            in2 => \_gnd_net_\,
            in3 => \N__39475\,
            lcout => \c0.n22128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1460_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38916\,
            in1 => \N__53465\,
            in2 => \_gnd_net_\,
            in3 => \N__48558\,
            lcout => OPEN,
            ltout => \c0.n22227_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1461_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39064\,
            in1 => \N__39015\,
            in2 => \N__38989\,
            in3 => \N__38985\,
            lcout => \c0.n10444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1700_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__38915\,
            in1 => \N__48557\,
            in2 => \N__44618\,
            in3 => \N__53464\,
            lcout => \c0.n6_adj_4312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1478_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38714\,
            in1 => \N__38847\,
            in2 => \_gnd_net_\,
            in3 => \N__39340\,
            lcout => \c0.n22477\,
            ltout => \c0.n22477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1480_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38812\,
            in3 => \N__40257\,
            lcout => \c0.n6_adj_4333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i28_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38800\,
            in1 => \N__42233\,
            in2 => \_gnd_net_\,
            in3 => \N__38771\,
            lcout => encoder0_position_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1432_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38715\,
            in2 => \_gnd_net_\,
            in3 => \N__40368\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1433_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39318\,
            in1 => \N__40209\,
            in2 => \N__39433\,
            in3 => \N__42338\,
            lcout => \c0.n20171\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1687_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__42337\,
            in1 => \N__40040\,
            in2 => \_gnd_net_\,
            in3 => \N__39893\,
            lcout => \c0.data_out_frame_29__7__N_847\,
            ltout => \c0.data_out_frame_29__7__N_847_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1477_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39317\,
            in1 => \N__39966\,
            in2 => \N__39397\,
            in3 => \N__39360\,
            lcout => \c0.n10_adj_4332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1425_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__39967\,
            in1 => \N__39319\,
            in2 => \N__42306\,
            in3 => \N__39894\,
            lcout => \c0.n21931\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx_transmit_5282_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110110001000"
        )
    port map (
            in0 => \N__40158\,
            in1 => \N__39166\,
            in2 => \N__40750\,
            in3 => \N__49203\,
            lcout => \c0.r_SM_Main_2_N_3755_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66697\,
            ce => 'H',
            sr => \N__40777\
        );

    \c0.i2_3_lut_adj_1649_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__40776\,
            in1 => \N__40081\,
            in2 => \_gnd_net_\,
            in3 => \N__40455\,
            lcout => \c0.n14322\,
            ltout => \c0.n14322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11334_2_lut_3_lut_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__40600\,
            in1 => \_gnd_net_\,
            in2 => \N__39205\,
            in3 => \N__42799\,
            lcout => \c0.n14871\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20360_4_lut_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010100010"
        )
    port map (
            in0 => \N__40456\,
            in1 => \N__51367\,
            in2 => \N__39190\,
            in3 => \N__39139\,
            lcout => \c0.n23975\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1631_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__47563\,
            in1 => \N__39160\,
            in2 => \N__52246\,
            in3 => \N__39148\,
            lcout => \c0.n17602\,
            ltout => \c0.n17602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_3_lut_4_lut_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100100010"
        )
    port map (
            in0 => \N__49202\,
            in1 => \N__51366\,
            in2 => \N__40084\,
            in3 => \N__40157\,
            lcout => \c0.n8_adj_4417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_7__6__5463_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49320\,
            in1 => \N__48734\,
            in2 => \N__42041\,
            in3 => \N__39847\,
            lcout => data_out_frame_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i26_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40039\,
            in1 => \N__42151\,
            in2 => \_gnd_net_\,
            in3 => \N__40075\,
            lcout => encoder0_position_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i8_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__39994\,
            in1 => \_gnd_net_\,
            in2 => \N__42203\,
            in3 => \N__40284\,
            lcout => encoder0_position_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_8__2__5459_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__48733\,
            in1 => \N__49321\,
            in2 => \N__39979\,
            in3 => \N__39933\,
            lcout => data_out_frame_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i25_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42150\,
            in1 => \N__39919\,
            in2 => \_gnd_net_\,
            in3 => \N__39889\,
            lcout => encoder0_position_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.byte_transmit_counter_5__I_0_Mux_6_i5_3_lut_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39846\,
            in1 => \N__48484\,
            in2 => \_gnd_net_\,
            in3 => \N__39832\,
            lcout => \c0.n5_adj_4350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i2_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39486\,
            in1 => \N__52069\,
            in2 => \_gnd_net_\,
            in3 => \N__44661\,
            lcout => control_mode_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66710\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1686_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__42375\,
            in1 => \N__40359\,
            in2 => \N__40294\,
            in3 => \N__42286\,
            lcout => \c0.n22032\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i144_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69840\,
            in1 => \N__68096\,
            in2 => \N__57444\,
            in3 => \N__68972\,
            lcout => \c0.data_in_frame_17_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4649_2_lut_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__48697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49201\,
            lcout => \c0.n8107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i25_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__69374\,
            in1 => \N__43215\,
            in2 => \_gnd_net_\,
            in3 => \N__40232\,
            lcout => data_in_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i197_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67622\,
            in1 => \N__65899\,
            in2 => \N__58938\,
            in3 => \N__63173\,
            lcout => \c0.data_in_frame_24_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i5_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40198\,
            in1 => \N__47644\,
            in2 => \_gnd_net_\,
            in3 => \N__44659\,
            lcout => control_mode_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66725\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1532_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__42744\,
            in1 => \N__42978\,
            in2 => \N__46174\,
            in3 => \N__40418\,
            lcout => \c0.n1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1684_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__40671\,
            in1 => \N__40624\,
            in2 => \N__40512\,
            in3 => \N__42610\,
            lcout => OPEN,
            ltout => \c0.n23215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1492_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__42880\,
            in1 => \N__42835\,
            in2 => \N__40174\,
            in3 => \N__40159\,
            lcout => \c0.n6_adj_4338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i18884_2_lut_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48788\,
            in2 => \_gnd_net_\,
            in3 => \N__50780\,
            lcout => \c0.n22575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_7_i3_2_lut_4_lut_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__50499\,
            in1 => \N__45178\,
            in2 => \N__50849\,
            in3 => \N__51371\,
            lcout => \c0.n3_adj_4465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1643_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__40576\,
            in1 => \N__42743\,
            in2 => \_gnd_net_\,
            in3 => \N__50498\,
            lcout => \c0.data_out_frame_0__7__N_2568\,
            ltout => \c0.data_out_frame_0__7__N_2568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1893_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110111"
        )
    port map (
            in0 => \N__40623\,
            in1 => \N__40505\,
            in2 => \N__40492\,
            in3 => \N__40670\,
            lcout => \c0.n1220\,
            ltout => \c0.n1220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_11_i3_2_lut_4_lut_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__51372\,
            in1 => \N__45331\,
            in2 => \N__40489\,
            in3 => \N__50500\,
            lcout => \c0.n3_adj_4458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14213_4_lut_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__40486\,
            in1 => \N__45081\,
            in2 => \N__46175\,
            in3 => \N__44821\,
            lcout => \c0.n5024\,
            ltout => \c0.n5024_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1592_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42584\,
            in2 => \N__40474\,
            in3 => \N__43279\,
            lcout => \c0.n21773\,
            ltout => \c0.n21773_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1458_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__42833\,
            in1 => \N__40453\,
            in2 => \N__40459\,
            in3 => \N__42884\,
            lcout => OPEN,
            ltout => \c0.n4_adj_4328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i1_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__40454\,
            in1 => \N__42955\,
            in2 => \N__40423\,
            in3 => \N__40420\,
            lcout => \c0.FRAME_MATCHER_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66752\,
            ce => 'H',
            sr => \N__40927\
        );

    \c0.FRAME_MATCHER_state_i0_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__51322\,
            in1 => \N__40393\,
            in2 => \N__40381\,
            in3 => \N__50537\,
            lcout => \c0.FRAME_MATCHER_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66752\,
            ce => 'H',
            sr => \N__40927\
        );

    \c0.i18974_4_lut_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__42793\,
            in1 => \N__40807\,
            in2 => \N__40798\,
            in3 => \N__40783\,
            lcout => \c0.n22665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1656_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__40628\,
            in1 => \N__40535\,
            in2 => \N__40597\,
            in3 => \N__42789\,
            lcout => \c0.n63_adj_4293\,
            ltout => \c0.n63_adj_4293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1670_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40749\,
            in2 => \N__40705\,
            in3 => \N__40701\,
            lcout => \c0.n21734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1528_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42611\,
            in2 => \_gnd_net_\,
            in3 => \N__42791\,
            lcout => OPEN,
            ltout => \c0.n84_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1525_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__43008\,
            in1 => \N__40687\,
            in2 => \N__40675\,
            in3 => \N__40672\,
            lcout => \c0.n7_adj_4344\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1663_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101110"
        )
    port map (
            in0 => \N__40629\,
            in1 => \N__40539\,
            in2 => \N__40598\,
            in3 => \N__42790\,
            lcout => \c0.n12992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_adj_1660_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__42792\,
            in1 => \N__40585\,
            in2 => \N__40540\,
            in3 => \N__40513\,
            lcout => \c0.n12991\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1644_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__42795\,
            in1 => \N__41146\,
            in2 => \N__42616\,
            in3 => \N__53128\,
            lcout => \c0.n8_adj_4396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i30_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41147\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52843\,
            lcout => \c0.FRAME_MATCHER_state_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66779\,
            ce => 'H',
            sr => \N__41122\
        );

    \c0.i1_2_lut_4_lut_adj_1779_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__42796\,
            in1 => \N__41003\,
            in2 => \N__42545\,
            in3 => \N__53129\,
            lcout => \c0.n21338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1646_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__53130\,
            in1 => \N__42615\,
            in2 => \N__41052\,
            in3 => \N__42797\,
            lcout => \c0.n8_adj_4398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1683_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__42825\,
            in1 => \N__43007\,
            in2 => \N__42886\,
            in3 => \N__42794\,
            lcout => \c0.n21737\,
            ltout => \c0.n21737_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1780_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__42538\,
            in1 => \N__42798\,
            in2 => \N__41107\,
            in3 => \N__41099\,
            lcout => \c0.n21340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i19_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41048\,
            in2 => \_gnd_net_\,
            in3 => \N__52845\,
            lcout => \c0.FRAME_MATCHER_state_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66791\,
            ce => 'H',
            sr => \N__41020\
        );

    \c0.FRAME_MATCHER_state_i12_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42928\,
            lcout => \c0.FRAME_MATCHER_state_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66801\,
            ce => 'H',
            sr => \N__42898\
        );

    \c0.FRAME_MATCHER_state_i5_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52848\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40996\,
            lcout => \c0.FRAME_MATCHER_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66811\,
            ce => 'H',
            sr => \N__40966\
        );

    \c0.i1_2_lut_3_lut_adj_1760_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__43393\,
            in1 => \N__53177\,
            in2 => \_gnd_net_\,
            in3 => \N__53022\,
            lcout => \c0.n21358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i132_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66013\,
            in1 => \N__68167\,
            in2 => \N__58130\,
            in3 => \N__64883\,
            lcout => \c0.data_in_frame_16_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66636\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20141_4_lut_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43921\,
            in1 => \N__50388\,
            in2 => \N__48168\,
            in3 => \N__43878\,
            lcout => \c0.n23836\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i4_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66014\,
            in1 => \N__60759\,
            in2 => \N__48153\,
            in3 => \N__64884\,
            lcout => \c0.data_in_frame_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66636\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1633_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43818\,
            in1 => \N__48046\,
            in2 => \N__52068\,
            in3 => \N__44698\,
            lcout => OPEN,
            ltout => \c0.n38_adj_4407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__41239\,
            in1 => \N__54420\,
            in2 => \N__41170\,
            in3 => \N__44166\,
            lcout => OPEN,
            ltout => \c0.n43_adj_4410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__41197\,
            in1 => \N__41167\,
            in2 => \N__41161\,
            in3 => \N__43549\,
            lcout => \FRAME_MATCHER_state_31_N_2976_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i65_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__69555\,
            in1 => \N__62379\,
            in2 => \N__65991\,
            in3 => \N__51938\,
            lcout => \c0.data_in_frame_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1855_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47906\,
            in1 => \N__51800\,
            in2 => \N__51942\,
            in3 => \N__51979\,
            lcout => \c0.n22443\,
            ltout => \c0.n22443_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1219_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52546\,
            in1 => \N__51819\,
            in2 => \N__41158\,
            in3 => \N__47844\,
            lcout => \c0.n13287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1301_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54747\,
            in2 => \_gnd_net_\,
            in3 => \N__54663\,
            lcout => \c0.n22283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1541_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41178\,
            in2 => \_gnd_net_\,
            in3 => \N__44099\,
            lcout => \c0.n21986\,
            ltout => \c0.n21986_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1715_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47623\,
            in1 => \N__48028\,
            in2 => \N__41182\,
            in3 => \N__47993\,
            lcout => \c0.n13180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3725_2_lut_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41278\,
            in2 => \_gnd_net_\,
            in3 => \N__53328\,
            lcout => \c0.n6404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i49_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41179\,
            in1 => \N__69556\,
            in2 => \_gnd_net_\,
            in3 => \N__49707\,
            lcout => data_in_frame_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66640\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i43_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62187\,
            in1 => \N__60766\,
            in2 => \N__43630\,
            in3 => \N__68354\,
            lcout => \c0.data_in_frame_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i29_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__60761\,
            in1 => \N__63226\,
            in2 => \N__43609\,
            in3 => \N__67460\,
            lcout => \c0.data_in_frame_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1538_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43591\,
            in1 => \N__43690\,
            in2 => \N__47788\,
            in3 => \N__43605\,
            lcout => \c0.n13237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i30_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__60762\,
            in1 => \N__67458\,
            in2 => \N__67209\,
            in3 => \N__47997\,
            lcout => \c0.data_in_frame_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i11_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69844\,
            in1 => \N__60764\,
            in2 => \N__52058\,
            in3 => \N__68353\,
            lcout => data_in_frame_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i31_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__60763\,
            in1 => \N__67459\,
            in2 => \N__44104\,
            in3 => \N__65582\,
            lcout => \c0.data_in_frame_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i12_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69845\,
            in1 => \N__60765\,
            in2 => \N__48047\,
            in3 => \N__64894\,
            lcout => data_in_frame_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i14_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__60760\,
            in1 => \N__69846\,
            in2 => \N__67208\,
            in3 => \N__47631\,
            lcout => data_in_frame_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1668_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47624\,
            in1 => \N__44297\,
            in2 => \N__43684\,
            in3 => \N__43810\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1601_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41254\,
            in1 => \N__41208\,
            in2 => \N__41188\,
            in3 => \N__44079\,
            lcout => \c0.n13086\,
            ltout => \c0.n13086_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47446\,
            in2 => \N__41185\,
            in3 => \N__47901\,
            lcout => \c0.n6_adj_4220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1593_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43724\,
            in2 => \_gnd_net_\,
            in3 => \N__43868\,
            lcout => \c0.n21893\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i18_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69231\,
            in1 => \N__63716\,
            in2 => \N__43729\,
            in3 => \N__60843\,
            lcout => \c0.data_in_frame_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i34_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__60842\,
            in1 => \N__44080\,
            in2 => \N__64551\,
            in3 => \N__63864\,
            lcout => \c0.data_in_frame_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i1_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__43869\,
            in1 => \N__69563\,
            in2 => \N__66012\,
            in3 => \N__60844\,
            lcout => \c0.data_in_frame_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1831_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51801\,
            in1 => \N__51978\,
            in2 => \N__47907\,
            in3 => \N__47239\,
            lcout => \c0.n22280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i51_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__68355\,
            in1 => \N__49691\,
            in2 => \_gnd_net_\,
            in3 => \N__43771\,
            lcout => data_in_frame_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i16_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69847\,
            in1 => \N__68958\,
            in2 => \N__44309\,
            in3 => \N__60835\,
            lcout => data_in_frame_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i15_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__60834\,
            in1 => \N__65674\,
            in2 => \N__69794\,
            in3 => \N__43817\,
            lcout => data_in_frame_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1634_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43728\,
            lcout => \c0.n25_adj_4408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1625_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47802\,
            in1 => \N__50413\,
            in2 => \N__41227\,
            in3 => \N__47246\,
            lcout => \c0.n16_adj_4401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1602_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__41209\,
            in1 => \N__43735\,
            in2 => \N__41581\,
            in3 => \N__44298\,
            lcout => \c0.n13043\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i56_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49692\,
            in1 => \N__68957\,
            in2 => \_gnd_net_\,
            in3 => \N__44255\,
            lcout => data_in_frame_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66660\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__44263\,
            in1 => \N__48088\,
            in2 => \N__51649\,
            in3 => \N__44449\,
            lcout => \c0.n44_adj_4409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1587_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44136\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43899\,
            lcout => \c0.n21791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i37_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__60849\,
            in1 => \N__64550\,
            in2 => \N__43756\,
            in3 => \N__63206\,
            lcout => \c0.data_in_frame_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i19_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69226\,
            in1 => \N__60850\,
            in2 => \N__44344\,
            in3 => \N__68426\,
            lcout => \c0.data_in_frame_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1575_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43833\,
            in1 => \N__44197\,
            in2 => \N__44185\,
            in3 => \N__43752\,
            lcout => \c0.n21934\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i20_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69227\,
            in1 => \N__60851\,
            in2 => \N__44048\,
            in3 => \N__64824\,
            lcout => \c0.data_in_frame_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i2_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__60848\,
            in1 => \N__43918\,
            in2 => \N__66015\,
            in3 => \N__63850\,
            lcout => \c0.data_in_frame_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i23_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__50381\,
            in1 => \N__60852\,
            in2 => \N__69244\,
            in3 => \N__65673\,
            lcout => \c0.data_in_frame_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i167_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__65672\,
            in1 => \N__68018\,
            in2 => \N__41277\,
            in3 => \N__64523\,
            lcout => \c0.data_in_frame_20_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1650_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__56605\,
            in1 => \N__56465\,
            in2 => \N__56748\,
            in3 => \N__60642\,
            lcout => n21744,
            ltout => \n21744_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i52_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64826\,
            in2 => \N__41257\,
            in3 => \N__41253\,
            lcout => data_in_frame_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i168_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__68017\,
            in1 => \N__64519\,
            in2 => \N__68973\,
            in3 => \N__53321\,
            lcout => \c0.data_in_frame_20_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i170_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62185\,
            in1 => \N__68019\,
            in2 => \N__53279\,
            in3 => \N__63855\,
            lcout => \c0.data_in_frame_21_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i42_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__63854\,
            in1 => \N__60644\,
            in2 => \N__44383\,
            in3 => \N__62186\,
            lcout => \c0.data_in_frame_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i40_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__60643\,
            in1 => \N__68940\,
            in2 => \N__64552\,
            in3 => \N__44401\,
            lcout => \c0.data_in_frame_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i63_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__54746\,
            in1 => \N__60645\,
            in2 => \N__68671\,
            in3 => \N__65671\,
            lcout => \c0.data_in_frame_7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66676\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i18_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42238\,
            in1 => \N__41305\,
            in2 => \_gnd_net_\,
            in3 => \N__41746\,
            lcout => encoder0_position_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1430_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41744\,
            lcout => \c0.n21816\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__46048\,
            in1 => \N__47320\,
            in2 => \N__45077\,
            in3 => \N__44728\,
            lcout => \c0.n21740\,
            ltout => \c0.n21740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i5_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__65932\,
            in1 => \N__63170\,
            in2 => \N__41281\,
            in3 => \N__50321\,
            lcout => \c0.data_in_frame_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_12_i3_2_lut_4_lut_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51470\,
            in1 => \N__51096\,
            in2 => \N__45384\,
            in3 => \N__50660\,
            lcout => \c0.n3_adj_4456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1459_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41745\,
            in1 => \N__41700\,
            in2 => \_gnd_net_\,
            in3 => \N__41650\,
            lcout => \c0.n21813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_4_i3_2_lut_4_lut_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51463\,
            in1 => \N__51011\,
            in2 => \N__45085\,
            in3 => \N__50664\,
            lcout => \c0.n3_adj_4470\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i54_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__67161\,
            in1 => \N__49693\,
            in2 => \_gnd_net_\,
            in3 => \N__41577\,
            lcout => data_in_frame_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66702\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_14_i3_2_lut_4_lut_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51464\,
            in1 => \N__51012\,
            in2 => \N__45439\,
            in3 => \N__50665\,
            lcout => \c0.n3_adj_4453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_8_i3_2_lut_4_lut_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__50666\,
            in1 => \N__45229\,
            in2 => \N__51089\,
            in3 => \N__51465\,
            lcout => \c0.n3_adj_4463\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i6_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41534\,
            in1 => \N__41492\,
            in2 => \_gnd_net_\,
            in3 => \N__41563\,
            lcout => \c0.tx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66702\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.tx.r_Clock_Count__i8_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__41512\,
            in1 => \N__41327\,
            in2 => \N__41497\,
            in3 => \N__41386\,
            lcout => \r_Clock_Count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66702\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i21_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41889\,
            in1 => \N__43157\,
            in2 => \_gnd_net_\,
            in3 => \N__41992\,
            lcout => data_in_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i210_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__63815\,
            in1 => \N__58766\,
            in2 => \N__69245\,
            in3 => \N__67610\,
            lcout => \c0.data_in_frame_26_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.count_i0_i22_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42265\,
            in1 => \N__42232\,
            in2 => \_gnd_net_\,
            in3 => \N__42030\,
            lcout => encoder0_position_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i13_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41993\,
            in1 => \N__43169\,
            in2 => \_gnd_net_\,
            in3 => \N__41950\,
            lcout => data_in_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14264_2_lut_3_lut_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__41923\,
            in1 => \N__43156\,
            in2 => \_gnd_net_\,
            in3 => \N__50929\,
            lcout => \c0.n17790\,
            ltout => \c0.n17790_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_adj_1895_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__45069\,
            in1 => \N__46054\,
            in2 => \N__41899\,
            in3 => \N__47323\,
            lcout => \c0.n21775\,
            ltout => \c0.n21775_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i218_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__50191\,
            in1 => \N__67407\,
            in2 => \N__41896\,
            in3 => \N__63816\,
            lcout => \c0.data_in_frame_27_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i29_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__63188\,
            in1 => \N__43170\,
            in2 => \_gnd_net_\,
            in3 => \N__41888\,
            lcout => data_in_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1562_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__42638\,
            in1 => \N__56599\,
            in2 => \N__56749\,
            in3 => \N__56466\,
            lcout => \c0.n19783\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i1_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41843\,
            in1 => \N__47700\,
            in2 => \_gnd_net_\,
            in3 => \N__44654\,
            lcout => control_mode_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i3_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41784\,
            in1 => \N__48058\,
            in2 => \_gnd_net_\,
            in3 => \N__44655\,
            lcout => control_mode_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i183_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__65698\,
            in1 => \N__62729\,
            in2 => \_gnd_net_\,
            in3 => \N__59200\,
            lcout => data_in_frame_22_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i4_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__54421\,
            in1 => \_gnd_net_\,
            in2 => \N__44662\,
            in3 => \N__42385\,
            lcout => control_mode_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66730\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i7_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42336\,
            in2 => \N__44320\,
            in3 => \N__44653\,
            lcout => control_mode_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i237_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__63123\,
            in1 => \N__44559\,
            in2 => \N__62205\,
            in3 => \N__67621\,
            lcout => \c0.data_in_frame_29_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_17_i3_2_lut_4_lut_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__50650\,
            in1 => \N__51398\,
            in2 => \N__45502\,
            in3 => \N__50826\,
            lcout => \c0.n3_adj_4448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_1388_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50059\,
            in1 => \N__44863\,
            in2 => \N__53956\,
            in3 => \N__44734\,
            lcout => n23726,
            ltout => \n23726_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i6_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__43822\,
            in1 => \_gnd_net_\,
            in2 => \N__42310\,
            in3 => \N__42293\,
            lcout => control_mode_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i235_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__67620\,
            in1 => \N__68395\,
            in2 => \N__44899\,
            in3 => \N__62197\,
            lcout => \c0.data_in_frame_29_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66744\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_19_i3_2_lut_4_lut_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__50778\,
            in1 => \N__51388\,
            in2 => \N__45535\,
            in3 => \N__50594\,
            lcout => \c0.n3_adj_4444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i206_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69864\,
            in1 => \N__67202\,
            in2 => \N__53598\,
            in3 => \N__67623\,
            lcout => \c0.data_in_frame_25_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66758\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1581_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__44817\,
            in1 => \N__46039\,
            in2 => \_gnd_net_\,
            in3 => \N__45073\,
            lcout => \c0.n12876\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_3_lut_4_lut_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__43342\,
            in1 => \N__43363\,
            in2 => \N__48953\,
            in3 => \N__50777\,
            lcout => \c0.n21022\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_18_i3_2_lut_4_lut_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__50779\,
            in1 => \N__51389\,
            in2 => \N__45583\,
            in3 => \N__50595\,
            lcout => \c0.n3_adj_4446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i233_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__62189\,
            in1 => \N__69487\,
            in2 => \N__44791\,
            in3 => \N__67624\,
            lcout => \c0.data_in_frame_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66758\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1531_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__42786\,
            in1 => \N__42585\,
            in2 => \N__42567\,
            in3 => \N__42409\,
            lcout => \c0.n5_adj_4342\,
            ltout => \c0.n5_adj_4342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i3_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__42494\,
            in1 => \_gnd_net_\,
            in2 => \N__42550\,
            in3 => \_gnd_net_\,
            lcout => \c0.FRAME_MATCHER_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66771\,
            ce => 'H',
            sr => \N__42445\
        );

    \c0.i3_3_lut_4_lut_adj_1749_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__43362\,
            in1 => \N__43345\,
            in2 => \N__48981\,
            in3 => \N__50802\,
            lcout => \c0.n21686\,
            ltout => \c0.n21686_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_4_lut_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__42493\,
            in1 => \N__53188\,
            in2 => \N__42448\,
            in3 => \N__42787\,
            lcout => \c0.n21334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1530_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__42785\,
            in1 => \N__42429\,
            in2 => \_gnd_net_\,
            in3 => \N__43344\,
            lcout => \c0.n1_adj_4349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i48_4_lut_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__43361\,
            in1 => \N__43343\,
            in2 => \N__43306\,
            in3 => \N__43290\,
            lcout => \c0.n45_adj_4389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_0___i26_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43031\,
            in1 => \N__43171\,
            in2 => \_gnd_net_\,
            in3 => \N__63769\,
            lcout => data_in_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1534_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__42649\,
            in1 => \N__43009\,
            in2 => \N__43502\,
            in3 => \N__53026\,
            lcout => \c0.n21332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14222_2_lut_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46158\,
            in2 => \_gnd_net_\,
            in3 => \N__42971\,
            lcout => \c0.n937\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i178_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44925\,
            in1 => \N__63768\,
            in2 => \_gnd_net_\,
            in3 => \N__59210\,
            lcout => data_in_frame_22_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1757_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__42935\,
            in1 => \N__53131\,
            in2 => \_gnd_net_\,
            in3 => \N__53019\,
            lcout => \c0.n21352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i179_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__68352\,
            in1 => \N__59310\,
            in2 => \_gnd_net_\,
            in3 => \N__59211\,
            lcout => data_in_frame_22_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66795\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1747_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__42885\,
            in1 => \N__42826\,
            in2 => \_gnd_net_\,
            in3 => \N__42788\,
            lcout => \c0.n7_adj_4356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1758_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__53020\,
            in1 => \_gnd_net_\,
            in2 => \N__53174\,
            in3 => \N__43451\,
            lcout => \c0.n21354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1777_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__43531\,
            in1 => \N__53135\,
            in2 => \_gnd_net_\,
            in3 => \N__53021\,
            lcout => \c0.n21378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i240_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__68880\,
            in1 => \N__50034\,
            in2 => \N__62204\,
            in3 => \N__67685\,
            lcout => \c0.data_in_frame_29_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66795\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i28_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43532\,
            in2 => \_gnd_net_\,
            in3 => \N__52744\,
            lcout => \c0.FRAME_MATCHER_state_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66805\,
            ce => 'H',
            sr => \N__43510\
        );

    \c0.FRAME_MATCHER_state_i31_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43487\,
            in2 => \_gnd_net_\,
            in3 => \N__52844\,
            lcout => \c0.FRAME_MATCHER_state_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66817\,
            ce => 'H',
            sr => \N__43465\
        );

    \c0.FRAME_MATCHER_state_i13_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43444\,
            in2 => \_gnd_net_\,
            in3 => \N__52846\,
            lcout => \c0.FRAME_MATCHER_state_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66829\,
            ce => 'H',
            sr => \N__43420\
        );

    \c0.FRAME_MATCHER_state_i15_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43394\,
            in2 => \_gnd_net_\,
            in3 => \N__52745\,
            lcout => \c0.FRAME_MATCHER_state_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66841\,
            ce => 'H',
            sr => \N__43372\
        );

    \c0.select_365_Select_0_i3_2_lut_4_lut_LC_18_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51451\,
            in1 => \N__51190\,
            in2 => \N__56719\,
            in3 => \N__50680\,
            lcout => \c0.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_5_i3_2_lut_4_lut_LC_18_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51471\,
            in1 => \N__51122\,
            in2 => \N__47391\,
            in3 => \N__50678\,
            lcout => \c0.n3_adj_4468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1680_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47725\,
            in1 => \N__43571\,
            in2 => \N__44703\,
            in3 => \N__51683\,
            lcout => \c0.n18_adj_4370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1550_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__43572\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47509\,
            lcout => \c0.n21957\,
            ltout => \c0.n21957_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1586_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43557\,
            in1 => \N__43579\,
            in2 => \N__43582\,
            in3 => \N__52054\,
            lcout => \c0.n13099\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1557_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51684\,
            in1 => \N__44695\,
            in2 => \_gnd_net_\,
            in3 => \N__47726\,
            lcout => \c0.n22287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i28_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__60867\,
            in1 => \N__67364\,
            in2 => \N__64893\,
            in3 => \N__43573\,
            lcout => \c0.data_in_frame_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i27_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67363\,
            in1 => \N__60869\,
            in2 => \N__47736\,
            in3 => \N__68410\,
            lcout => \c0.data_in_frame_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i45_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__60868\,
            in1 => \N__63204\,
            in2 => \N__43561\,
            in3 => \N__62188\,
            lcout => \c0.data_in_frame_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i9_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__44702\,
            in1 => \N__69567\,
            in2 => \N__69777\,
            in3 => \N__60870\,
            lcout => data_in_frame_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20143_4_lut_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47540\,
            in1 => \N__44050\,
            in2 => \N__44505\,
            in3 => \N__47501\,
            lcout => \c0.n23838\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1603_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51685\,
            in1 => \N__44696\,
            in2 => \_gnd_net_\,
            in3 => \N__43644\,
            lcout => \c0.n21902\,
            ltout => \c0.n21902_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1609_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44697\,
            in1 => \N__51776\,
            in2 => \N__43651\,
            in3 => \N__47539\,
            lcout => \c0.n21992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i24_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69168\,
            in1 => \N__68956\,
            in2 => \N__47547\,
            in3 => \N__60896\,
            lcout => \c0.data_in_frame_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i25_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__60894\,
            in1 => \N__69548\,
            in2 => \N__43648\,
            in3 => \N__67379\,
            lcout => \c0.data_in_frame_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1540_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43636\,
            in1 => \N__47762\,
            in2 => \N__43629\,
            in3 => \N__47500\,
            lcout => \c0.n10_adj_4363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i7_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__60895\,
            in1 => \N__51686\,
            in2 => \N__65647\,
            in3 => \N__65969\,
            lcout => \c0.data_in_frame_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i26_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67362\,
            in1 => \N__60846\,
            in2 => \N__47767\,
            in3 => \N__63863\,
            lcout => \c0.data_in_frame_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1679_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54400\,
            in1 => \N__52034\,
            in2 => \N__47693\,
            in3 => \N__48026\,
            lcout => OPEN,
            ltout => \c0.n21879_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1566_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61092\,
            in1 => \N__47758\,
            in2 => \N__43612\,
            in3 => \N__44355\,
            lcout => \c0.n29_adj_4374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1554_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47992\,
            in2 => \_gnd_net_\,
            in3 => \N__43604\,
            lcout => \c0.n22051\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i8_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__47493\,
            in1 => \N__68955\,
            in2 => \N__66029\,
            in3 => \N__60847\,
            lcout => \c0.data_in_frame_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i38_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__60845\,
            in1 => \N__64532\,
            in2 => \N__67210\,
            in3 => \N__61093\,
            lcout => \c0.data_in_frame_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66655\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1612_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51775\,
            in2 => \N__47508\,
            in3 => \N__51687\,
            lcout => \c0.n22194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1556_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47684\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48027\,
            lcout => \c0.n22290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1590_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49597\,
            in2 => \_gnd_net_\,
            in3 => \N__43970\,
            lcout => \c0.n22258\,
            ltout => \c0.n22258_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1569_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44221\,
            in1 => \N__47615\,
            in2 => \N__43675\,
            in3 => \N__51990\,
            lcout => OPEN,
            ltout => \c0.n27_adj_4377_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1570_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43672\,
            in1 => \N__43927\,
            in2 => \N__43666\,
            in3 => \N__43696\,
            lcout => \c0.n14072\,
            ltout => \c0.n14072_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1549_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43663\,
            in3 => \N__54363\,
            lcout => \c0.n13852\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1672_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47616\,
            in1 => \N__43951\,
            in2 => \N__48208\,
            in3 => \N__43660\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1583_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43971\,
            in1 => \N__44419\,
            in2 => \N__43654\,
            in3 => \N__43809\,
            lcout => \c0.n14113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1605_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48139\,
            in2 => \_gnd_net_\,
            in3 => \N__50339\,
            lcout => \c0.n21803\,
            ltout => \c0.n21803_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1559_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43945\,
            in1 => \N__43936\,
            in2 => \N__43930\,
            in3 => \N__44014\,
            lcout => \c0.n30_adj_4371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1551_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__44336\,
            in1 => \N__43900\,
            in2 => \N__43879\,
            in3 => \_gnd_net_\,
            lcout => \c0.n13376\,
            ltout => \c0.n13376_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1560_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43806\,
            in2 => \N__43837\,
            in3 => \N__44292\,
            lcout => \c0.n22320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1669_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43808\,
            in1 => \N__43834\,
            in2 => \N__44308\,
            in3 => \N__44444\,
            lcout => \c0.n6_adj_4386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1594_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__47632\,
            in1 => \N__44293\,
            in2 => \_gnd_net_\,
            in3 => \N__43807\,
            lcout => OPEN,
            ltout => \c0.n13386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1621_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54367\,
            in1 => \N__43770\,
            in2 => \N__43759\,
            in3 => \N__44065\,
            lcout => \c0.n13033\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1607_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__43751\,
            in1 => \N__49634\,
            in2 => \N__44049\,
            in3 => \N__44012\,
            lcout => \c0.n22261\,
            ltout => \c0.n22261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1561_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44064\,
            in1 => \N__43723\,
            in2 => \N__43705\,
            in3 => \N__43702\,
            lcout => \c0.n28_adj_4372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1558_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44443\,
            in1 => \N__44103\,
            in2 => \_gnd_net_\,
            in3 => \N__44078\,
            lcout => \c0.n22218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1553_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44203\,
            in1 => \N__44398\,
            in2 => \N__44541\,
            in3 => \N__44191\,
            lcout => \c0.n21928\,
            ltout => \c0.n21928_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1542_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44053\,
            in3 => \N__44469\,
            lcout => \c0.n13861\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1595_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44038\,
            in1 => \N__44013\,
            in2 => \N__44542\,
            in3 => \N__48089\,
            lcout => \c0.n21882\,
            ltout => \c0.n21882_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1539_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43993\,
            in3 => \N__61103\,
            lcout => \c0.data_out_frame_0__7__N_2744\,
            ltout => \c0.data_out_frame_0__7__N_2744_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44362\,
            in1 => \N__48090\,
            in2 => \N__43978\,
            in3 => \N__44399\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4272_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1334_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44379\,
            in1 => \N__44251\,
            in2 => \N__43975\,
            in3 => \N__54815\,
            lcout => \c0.n22069\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i32_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__60823\,
            in1 => \N__67361\,
            in2 => \N__43972\,
            in3 => \N__68975\,
            lcout => \c0.data_in_frame_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1537_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44400\,
            in1 => \N__44378\,
            in2 => \N__48094\,
            in3 => \N__44361\,
            lcout => \c0.n4_adj_4255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_adj_1632_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__50307\,
            in1 => \N__47701\,
            in2 => \N__44343\,
            in3 => \N__44310\,
            lcout => \c0.n39_adj_4406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1330_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__44256\,
            in1 => \N__61124\,
            in2 => \_gnd_net_\,
            in3 => \N__44227\,
            lcout => \c0.n14037\,
            ltout => \c0.n14037_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1787_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__44220\,
            in1 => \_gnd_net_\,
            in2 => \N__44206\,
            in3 => \N__44468\,
            lcout => \c0.n22108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1681_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__44491\,
            in1 => \N__48154\,
            in2 => \N__44146\,
            in3 => \N__50368\,
            lcout => \c0.n6_adj_4369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1552_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44135\,
            in2 => \N__48169\,
            in3 => \N__44492\,
            lcout => \c0.n5_adj_4368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__5__I_0_2_lut_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51774\,
            in2 => \_gnd_net_\,
            in3 => \N__50306\,
            lcout => \c0.data_out_frame_29__7__N_1474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i55_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__65649\,
            in1 => \N__49674\,
            in2 => \_gnd_net_\,
            in3 => \N__44181\,
            lcout => data_in_frame_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i3_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__60715\,
            in1 => \N__65865\,
            in2 => \N__68411\,
            in3 => \N__44145\,
            lcout => \c0.data_in_frame_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i21_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69212\,
            in1 => \N__60756\,
            in2 => \N__44506\,
            in3 => \N__63171\,
            lcout => \c0.data_in_frame_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_9_i3_2_lut_4_lut_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__51444\,
            in1 => \N__50659\,
            in2 => \N__45280\,
            in3 => \N__50962\,
            lcout => \c0.n3_adj_4462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i41_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__69559\,
            in1 => \N__60757\,
            in2 => \N__44473\,
            in3 => \N__62198\,
            lcout => \c0.data_in_frame_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1202_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62590\,
            in1 => \N__65155\,
            in2 => \N__62822\,
            in3 => \N__63388\,
            lcout => \c0.n22057\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i48_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__68944\,
            in1 => \N__60758\,
            in2 => \N__62206\,
            in3 => \N__47883\,
            lcout => \c0.data_in_frame_5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_6_i3_2_lut_4_lut_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__51443\,
            in1 => \N__50658\,
            in2 => \N__47359\,
            in3 => \N__50961\,
            lcout => \c0.n3_adj_4467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1574_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47355\,
            in1 => \N__45225\,
            in2 => \N__47401\,
            in3 => \N__45534\,
            lcout => \c0.n28_adj_4381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i17_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__60755\,
            in1 => \N__69213\,
            in2 => \N__44448\,
            in3 => \N__69558\,
            lcout => \c0.data_in_frame_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i204_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__64698\,
            in1 => \N__53626\,
            in2 => \N__69866\,
            in3 => \N__67611\,
            lcout => \c0.data_in_frame_25_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i50_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__63781\,
            in1 => \N__49703\,
            in2 => \_gnd_net_\,
            in3 => \N__44415\,
            lcout => data_in_frame_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i177_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__69486\,
            in1 => \N__62815\,
            in2 => \_gnd_net_\,
            in3 => \N__59169\,
            lcout => data_in_frame_22_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i36_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__64818\,
            in1 => \N__60714\,
            in2 => \N__49642\,
            in3 => \N__64531\,
            lcout => \c0.data_in_frame_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_1176_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59883\,
            in2 => \_gnd_net_\,
            in3 => \N__57105\,
            lcout => n4,
            ltout => \n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i2_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__59694\,
            in1 => \N__68289\,
            in2 => \N__44545\,
            in3 => \N__59944\,
            lcout => rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i39_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__60713\,
            in1 => \N__65697\,
            in2 => \N__64556\,
            in3 => \N__44534\,
            lcout => \c0.data_in_frame_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i3_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__44518\,
            in1 => \N__64699\,
            in2 => \N__59710\,
            in3 => \N__56221\,
            lcout => rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66717\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_16_i3_2_lut_4_lut_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51448\,
            in1 => \N__50954\,
            in2 => \N__49897\,
            in3 => \N__50651\,
            lcout => \c0.n3_adj_4450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_adj_1466_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__46049\,
            in1 => \N__45064\,
            in2 => \N__47321\,
            in3 => \N__44723\,
            lcout => \c0.n21758\,
            ltout => \c0.n21758_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i162_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__63814\,
            in1 => \N__64527\,
            in2 => \N__44509\,
            in3 => \N__53241\,
            lcout => \c0.data_in_frame_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66731\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_4_lut_adj_1457_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__46050\,
            in1 => \N__45065\,
            in2 => \N__47322\,
            in3 => \N__44724\,
            lcout => \c0.n21749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1240_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55432\,
            in2 => \_gnd_net_\,
            in3 => \N__61430\,
            lcout => \c0.n22308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i212_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__64700\,
            in1 => \N__57987\,
            in2 => \N__69253\,
            in3 => \N__67678\,
            lcout => \c0.data_in_frame_26_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66731\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i234_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__67609\,
            in1 => \N__44880\,
            in2 => \N__62190\,
            in3 => \N__63825\,
            lcout => \c0.data_in_frame_29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1571_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45327\,
            in1 => \N__45174\,
            in2 => \N__45385\,
            in3 => \N__45435\,
            lcout => \c0.n17_adj_4378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i141_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__63145\,
            in1 => \N__67912\,
            in2 => \N__69881\,
            in3 => \N__55375\,
            lcout => \c0.data_in_frame_17_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.control_mode_i0_i0_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44591\,
            in1 => \N__44710\,
            in2 => \_gnd_net_\,
            in3 => \N__44660\,
            lcout => control_mode_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_97_i9_2_lut_3_lut_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__56467\,
            in1 => \_gnd_net_\,
            in2 => \N__56744\,
            in3 => \N__56600\,
            lcout => \c0.n9_adj_4278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i137_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69860\,
            in1 => \N__67911\,
            in2 => \N__55627\,
            in3 => \N__69491\,
            lcout => \c0.data_in_frame_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66745\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1376_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56057\,
            in1 => \N__56279\,
            in2 => \N__44560\,
            in3 => \N__53743\,
            lcout => \c0.n23523\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1362_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58609\,
            in1 => \N__65326\,
            in2 => \N__44803\,
            in3 => \N__64990\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4286_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1374_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__54016\,
            in1 => \_gnd_net_\,
            in2 => \N__44806\,
            in3 => \N__59983\,
            lcout => \c0.n23389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i190_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__68632\,
            in1 => \N__67206\,
            in2 => \N__68044\,
            in3 => \N__49919\,
            lcout => \c0.data_in_frame_23_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i227_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__67731\,
            in1 => \N__44802\,
            in2 => \N__64567\,
            in3 => \N__68394\,
            lcout => \c0.data_in_frame_28_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i230_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__64566\,
            in1 => \N__67207\,
            in2 => \N__58377\,
            in3 => \N__67733\,
            lcout => \c0.data_in_frame_28_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i203_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68393\,
            in1 => \N__69865\,
            in2 => \N__53694\,
            in3 => \N__67732\,
            lcout => \c0.data_in_frame_25_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1375_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011101101"
        )
    port map (
            in0 => \N__44790\,
            in1 => \N__44773\,
            in2 => \N__53533\,
            in3 => \N__58866\,
            lcout => OPEN,
            ltout => \c0.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1378_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__59461\,
            in1 => \N__56233\,
            in2 => \N__44755\,
            in3 => \N__44752\,
            lcout => OPEN,
            ltout => \c0.n32_adj_4295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1386_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__58357\,
            in1 => \N__54070\,
            in2 => \N__44746\,
            in3 => \N__44743\,
            lcout => \c0.n34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1367_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58867\,
            in1 => \N__55798\,
            in2 => \N__44898\,
            in3 => \N__50205\,
            lcout => OPEN,
            ltout => \c0.n23388_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1385_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__53532\,
            in1 => \N__44881\,
            in2 => \N__44866\,
            in3 => \N__64972\,
            lcout => \c0.n30_adj_4299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1577_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49822\,
            in1 => \N__45838\,
            in2 => \N__45802\,
            in3 => \N__45715\,
            lcout => \c0.n27_adj_4383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_adj_1568_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__45877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45279\,
            lcout => OPEN,
            ltout => \c0.n15_adj_4376_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1572_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50157\,
            in1 => \N__49873\,
            in2 => \N__44857\,
            in3 => \N__44854\,
            lcout => OPEN,
            ltout => \c0.n18_adj_4379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1573_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45630\,
            in1 => \N__45498\,
            in2 => \N__44845\,
            in3 => \N__45579\,
            lcout => OPEN,
            ltout => \c0.n30_adj_4380_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1579_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44842\,
            in1 => \N__44965\,
            in2 => \N__44836\,
            in3 => \N__44833\,
            lcout => \c0.n13000\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20_4_lut_adj_1731_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__66136\,
            in1 => \N__59117\,
            in2 => \N__56149\,
            in3 => \N__53560\,
            lcout => \c0.n49_adj_4488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_22_i3_2_lut_4_lut_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__50646\,
            in1 => \N__51412\,
            in2 => \N__51070\,
            in3 => \N__45675\,
            lcout => \c0.n3_adj_4438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_21_i3_2_lut_4_lut_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51413\,
            in1 => \N__50987\,
            in2 => \N__45640\,
            in3 => \N__50647\,
            lcout => \c0.n3_adj_4440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i220_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__67403\,
            in1 => \N__64823\,
            in2 => \N__56284\,
            in3 => \N__67762\,
            lcout => \c0.data_in_frame_27_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i211_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__67760\,
            in1 => \N__59118\,
            in2 => \N__69234\,
            in3 => \N__68359\,
            lcout => \c0.data_in_frame_26_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i219_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68358\,
            in1 => \N__67452\,
            in2 => \N__56058\,
            in3 => \N__67761\,
            lcout => \c0.data_in_frame_27_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1213_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59306\,
            in2 => \_gnd_net_\,
            in3 => \N__44921\,
            lcout => \c0.n22191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_23_i3_2_lut_4_lut_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51450\,
            in1 => \N__51068\,
            in2 => \N__45714\,
            in3 => \N__50649\,
            lcout => \c0.n3_adj_4436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i18920_2_lut_3_lut_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__56826\,
            in1 => \N__59655\,
            in2 => \_gnd_net_\,
            in3 => \N__56187\,
            lcout => OPEN,
            ltout => \c0.rx.n22611_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_adj_1172_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001011"
        )
    port map (
            in0 => \N__57061\,
            in1 => \N__56927\,
            in2 => \N__44905\,
            in3 => \N__57007\,
            lcout => \c0.rx.n17411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_3_lut_4_lut_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__56827\,
            in1 => \N__59653\,
            in2 => \N__56938\,
            in3 => \N__56188\,
            lcout => OPEN,
            ltout => \c0.rx.n8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i18819_4_lut_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__59654\,
            in1 => \N__57008\,
            in2 => \N__44902\,
            in3 => \N__56828\,
            lcout => \c0.rx.n14391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_24_i3_2_lut_4_lut_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51449\,
            in1 => \N__51067\,
            in2 => \N__45760\,
            in3 => \N__50648\,
            lcout => \c0.n3_adj_4435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_30_i3_2_lut_4_lut_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__51403\,
            in1 => \N__50969\,
            in2 => \N__50679\,
            in3 => \N__45943\,
            lcout => \c0.n3_adj_4426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1576_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45676\,
            in1 => \N__45903\,
            in2 => \N__45759\,
            in3 => \N__45942\,
            lcout => \c0.n29_adj_4382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_31_i3_2_lut_4_lut_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__50667\,
            in1 => \N__46147\,
            in2 => \N__51065\,
            in3 => \N__51402\,
            lcout => \c0.n3_adj_4421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_18_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_25_i3_2_lut_4_lut_LC_18_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51410\,
            in1 => \N__50973\,
            in2 => \N__45798\,
            in3 => \N__50669\,
            lcout => \c0.n3_adj_4434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_29_i3_2_lut_4_lut_LC_18_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__50668\,
            in1 => \N__51409\,
            in2 => \N__51066\,
            in3 => \N__45904\,
            lcout => \c0.n3_adj_4428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_26_i3_2_lut_4_lut_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__50980\,
            in1 => \N__51411\,
            in2 => \N__45837\,
            in3 => \N__50674\,
            lcout => \c0.n3_adj_4433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_27_i3_2_lut_4_lut_LC_18_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51475\,
            in1 => \N__50974\,
            in2 => \N__45876\,
            in3 => \N__50673\,
            lcout => \c0.n3_adj_4432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i0_LC_19_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1001011000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56630\,
            in2 => \N__44953\,
            in3 => \N__51173\,
            lcout => \c0.FRAME_MATCHER_i_0\,
            ltout => OPEN,
            carryin => \bfn_19_1_0_\,
            carryout => \c0.n19442\,
            clk => \N__66630\,
            ce => 'H',
            sr => \N__44980\
        );

    \c0.add_49_2_THRU_CRY_0_LC_19_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47190\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19442\,
            carryout => \c0.n19442_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_1_LC_19_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47215\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19442_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19442_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_2_LC_19_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47194\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19442_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19442_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_3_LC_19_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47216\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19442_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19442_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_4_LC_19_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47198\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19442_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19442_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_5_LC_19_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47217\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19442_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19442_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_2_THRU_CRY_6_LC_19_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47202\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19442_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19442_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i1_LC_19_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51100\,
            in1 => \N__56495\,
            in2 => \_gnd_net_\,
            in3 => \N__44968\,
            lcout => \c0.FRAME_MATCHER_i_1\,
            ltout => OPEN,
            carryin => \bfn_19_2_0_\,
            carryout => \c0.n19443\,
            clk => \N__66631\,
            ce => 'H',
            sr => \N__46060\
        );

    \c0.add_49_3_THRU_CRY_0_LC_19_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47177\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19443\,
            carryout => \c0.n19443_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_1_LC_19_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47212\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19443_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19443_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_2_LC_19_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47181\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19443_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19443_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_3_LC_19_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47213\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19443_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19443_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_4_LC_19_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47185\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19443_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19443_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_5_LC_19_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47214\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19443_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19443_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_3_THRU_CRY_6_LC_19_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47189\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19443_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19443_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i2_LC_19_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51191\,
            in1 => \N__56353\,
            in2 => \_gnd_net_\,
            in3 => \N__44983\,
            lcout => \c0.FRAME_MATCHER_i_2\,
            ltout => OPEN,
            carryin => \bfn_19_3_0_\,
            carryout => \c0.n19444\,
            clk => \N__66632\,
            ce => 'H',
            sr => \N__47413\
        );

    \c0.add_49_4_THRU_CRY_0_LC_19_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47164\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19444\,
            carryout => \c0.n19444_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_1_LC_19_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47209\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19444_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19444_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_2_LC_19_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47168\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19444_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19444_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_3_LC_19_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47210\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19444_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19444_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_4_LC_19_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47172\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19444_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19444_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_5_LC_19_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47211\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19444_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19444_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_4_THRU_CRY_6_LC_19_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47176\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19444_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19444_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i3_LC_19_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51160\,
            in1 => \N__45999\,
            in2 => \_gnd_net_\,
            in3 => \N__44986\,
            lcout => \c0.FRAME_MATCHER_i_3\,
            ltout => OPEN,
            carryin => \bfn_19_4_0_\,
            carryout => \c0.n19445\,
            clk => \N__66633\,
            ce => 'H',
            sr => \N__45964\
        );

    \c0.add_49_5_THRU_CRY_0_LC_19_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47151\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19445\,
            carryout => \c0.n19445_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_1_LC_19_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47206\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19445_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19445_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_2_LC_19_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47155\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19445_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19445_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_3_LC_19_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47207\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19445_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19445_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_4_LC_19_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47159\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19445_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19445_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_5_LC_19_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47208\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19445_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19445_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_5_THRU_CRY_6_LC_19_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47163\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19445_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19445_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i4_LC_19_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51175\,
            in1 => \N__45018\,
            in2 => \_gnd_net_\,
            in3 => \N__45007\,
            lcout => \c0.FRAME_MATCHER_i_4\,
            ltout => OPEN,
            carryin => \bfn_19_5_0_\,
            carryout => \c0.n19446\,
            clk => \N__66635\,
            ce => 'H',
            sr => \N__45004\
        );

    \c0.add_49_6_THRU_CRY_0_LC_19_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47063\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19446\,
            carryout => \c0.n19446_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_1_LC_19_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47148\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19446_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19446_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_2_LC_19_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47067\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19446_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19446_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_3_LC_19_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47149\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19446_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19446_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_4_LC_19_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47071\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19446_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19446_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_5_LC_19_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47150\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19446_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19446_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_6_THRU_CRY_6_LC_19_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47075\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19446_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19446_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i5_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51174\,
            in1 => \N__47380\,
            in2 => \_gnd_net_\,
            in3 => \N__45100\,
            lcout => \c0.FRAME_MATCHER_i_5\,
            ltout => OPEN,
            carryin => \bfn_19_6_0_\,
            carryout => \c0.n19447\,
            clk => \N__66637\,
            ce => 'H',
            sr => \N__45097\
        );

    \c0.add_49_7_THRU_CRY_0_LC_19_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47050\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19447\,
            carryout => \c0.n19447_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_1_LC_19_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47145\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19447_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19447_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_2_LC_19_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47054\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19447_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19447_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_3_LC_19_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47146\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19447_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19447_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_4_LC_19_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47058\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19447_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19447_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_5_LC_19_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47147\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19447_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19447_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_7_THRU_CRY_6_LC_19_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47062\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19447_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19447_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i6_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51172\,
            in1 => \N__47348\,
            in2 => \_gnd_net_\,
            in3 => \N__45118\,
            lcout => \c0.FRAME_MATCHER_i_6\,
            ltout => OPEN,
            carryin => \bfn_19_7_0_\,
            carryout => \c0.n19448\,
            clk => \N__66642\,
            ce => 'H',
            sr => \N__45115\
        );

    \c0.add_49_8_THRU_CRY_0_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47037\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19448\,
            carryout => \c0.n19448_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_1_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47142\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19448_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19448_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_2_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47041\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19448_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19448_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_3_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47143\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19448_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19448_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_4_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47045\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19448_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19448_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_5_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47144\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19448_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19448_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_8_THRU_CRY_6_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47049\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19448_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19448_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i7_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51064\,
            in1 => \N__45155\,
            in2 => \_gnd_net_\,
            in3 => \N__45139\,
            lcout => \c0.FRAME_MATCHER_i_7\,
            ltout => OPEN,
            carryin => \bfn_19_8_0_\,
            carryout => \c0.n19449\,
            clk => \N__66649\,
            ce => 'H',
            sr => \N__45136\
        );

    \c0.add_49_9_THRU_CRY_0_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47024\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19449\,
            carryout => \c0.n19449_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_1_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47139\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19449_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19449_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_2_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47028\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19449_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19449_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_3_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47140\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19449_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19449_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_4_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47032\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19449_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19449_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_5_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47141\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19449_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19449_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_9_THRU_CRY_6_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47036\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19449_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19449_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i8_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51193\,
            in1 => \N__45215\,
            in2 => \_gnd_net_\,
            in3 => \N__45196\,
            lcout => \c0.FRAME_MATCHER_i_8\,
            ltout => OPEN,
            carryin => \bfn_19_9_0_\,
            carryout => \c0.n19450\,
            clk => \N__66656\,
            ce => 'H',
            sr => \N__45193\
        );

    \c0.add_49_10_THRU_CRY_0_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46927\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19450\,
            carryout => \c0.n19450_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_1_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47021\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19450_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19450_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_2_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46931\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19450_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19450_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_3_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47022\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19450_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19450_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_4_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46935\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19450_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19450_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_5_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47023\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19450_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19450_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_10_THRU_CRY_6_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46939\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19450_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19450_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i9_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51192\,
            in1 => \N__45266\,
            in2 => \_gnd_net_\,
            in3 => \N__45250\,
            lcout => \c0.FRAME_MATCHER_i_9\,
            ltout => OPEN,
            carryin => \bfn_19_10_0_\,
            carryout => \c0.n19451\,
            clk => \N__66661\,
            ce => 'H',
            sr => \N__45247\
        );

    \c0.add_49_11_THRU_CRY_0_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46914\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19451\,
            carryout => \c0.n19451_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_1_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47018\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19451_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19451_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_2_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46918\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19451_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19451_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_3_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47019\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19451_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19451_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_4_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46922\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19451_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19451_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_5_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47020\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19451_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19451_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_11_THRU_CRY_6_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46926\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19451_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19451_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i10_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51204\,
            in1 => \N__50138\,
            in2 => \_gnd_net_\,
            in3 => \N__45232\,
            lcout => \c0.FRAME_MATCHER_i_10\,
            ltout => OPEN,
            carryin => \bfn_19_11_0_\,
            carryout => \c0.n19452\,
            clk => \N__66667\,
            ce => 'H',
            sr => \N__50122\
        );

    \c0.add_49_12_THRU_CRY_0_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46901\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19452\,
            carryout => \c0.n19452_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_1_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47015\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19452_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19452_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_2_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46905\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19452_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19452_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_3_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47016\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19452_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19452_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_4_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46909\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19452_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19452_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_5_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47017\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19452_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19452_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_12_THRU_CRY_6_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46913\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19452_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19452_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i11_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51203\,
            in1 => \N__45314\,
            in2 => \_gnd_net_\,
            in3 => \N__45301\,
            lcout => \c0.FRAME_MATCHER_i_11\,
            ltout => OPEN,
            carryin => \bfn_19_12_0_\,
            carryout => \c0.n19453\,
            clk => \N__66678\,
            ce => 'H',
            sr => \N__45298\
        );

    \c0.add_49_13_THRU_CRY_0_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46888\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19453\,
            carryout => \c0.n19453_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_1_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47012\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19453_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19453_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_2_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46892\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19453_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19453_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_3_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47013\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19453_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19453_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_4_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46896\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19453_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19453_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_5_LC_19_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__47014\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19453_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19453_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_13_THRU_CRY_6_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46900\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19453_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19453_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i12_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51205\,
            in1 => \N__45362\,
            in2 => \_gnd_net_\,
            in3 => \N__45346\,
            lcout => \c0.FRAME_MATCHER_i_12\,
            ltout => OPEN,
            carryin => \bfn_19_13_0_\,
            carryout => \c0.n19454\,
            clk => \N__66690\,
            ce => 'H',
            sr => \N__45343\
        );

    \c0.add_49_14_THRU_CRY_0_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46789\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19454\,
            carryout => \c0.n19454_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_1_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46885\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19454_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19454_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_2_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46793\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19454_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19454_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_3_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46886\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19454_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19454_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_4_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46797\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19454_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19454_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_5_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46887\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19454_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19454_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_14_THRU_CRY_6_LC_19_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46801\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19454_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19454_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i13_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51113\,
            in1 => \N__49851\,
            in2 => \_gnd_net_\,
            in3 => \N__45388\,
            lcout => \c0.FRAME_MATCHER_i_13\,
            ltout => OPEN,
            carryin => \bfn_19_14_0_\,
            carryout => \c0.n19455\,
            clk => \N__66704\,
            ce => 'H',
            sr => \N__49837\
        );

    \c0.add_49_15_THRU_CRY_0_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46776\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19455\,
            carryout => \c0.n19455_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_1_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46882\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19455_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19455_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_2_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46780\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19455_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19455_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_3_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46883\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19455_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19455_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_4_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46784\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19455_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19455_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_5_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46884\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19455_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19455_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_15_THRU_CRY_6_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46788\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19455_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19455_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i14_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51097\,
            in1 => \N__45425\,
            in2 => \_gnd_net_\,
            in3 => \N__45406\,
            lcout => \c0.FRAME_MATCHER_i_14\,
            ltout => OPEN,
            carryin => \bfn_19_15_0_\,
            carryout => \c0.n19456\,
            clk => \N__66718\,
            ce => 'H',
            sr => \N__45403\
        );

    \c0.add_49_16_THRU_CRY_0_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46763\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19456\,
            carryout => \c0.n19456_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_1_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46879\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19456_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19456_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_2_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46767\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19456_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19456_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_3_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46880\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19456_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19456_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_4_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46771\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19456_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19456_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_5_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46881\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19456_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19456_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_16_THRU_CRY_6_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46775\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19456_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19456_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i15_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51112\,
            in1 => \N__49814\,
            in2 => \_gnd_net_\,
            in3 => \N__45442\,
            lcout => \c0.FRAME_MATCHER_i_15\,
            ltout => OPEN,
            carryin => \bfn_19_16_0_\,
            carryout => \c0.n19457\,
            clk => \N__66732\,
            ce => 'H',
            sr => \N__49795\
        );

    \c0.add_49_17_THRU_CRY_0_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46750\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19457\,
            carryout => \c0.n19457_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_1_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46876\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19457_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19457_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_2_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46754\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19457_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19457_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_3_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46877\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19457_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19457_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_4_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46758\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19457_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19457_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_5_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46878\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19457_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19457_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_17_THRU_CRY_6_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46762\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19457_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19457_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i16_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__50955\,
            in1 => \N__49889\,
            in2 => \_gnd_net_\,
            in3 => \N__45454\,
            lcout => \c0.FRAME_MATCHER_i_16\,
            ltout => OPEN,
            carryin => \bfn_19_17_0_\,
            carryout => \c0.n19458\,
            clk => \N__66746\,
            ce => 'H',
            sr => \N__45451\
        );

    \c0.add_49_18_THRU_CRY_0_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46654\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19458\,
            carryout => \c0.n19458_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_1_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46747\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19458_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19458_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_2_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46658\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19458_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19458_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_3_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46748\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19458_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19458_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_4_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46662\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19458_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19458_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_5_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46749\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19458_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19458_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_18_THRU_CRY_6_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46666\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19458_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19458_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i17_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51054\,
            in1 => \N__45491\,
            in2 => \_gnd_net_\,
            in3 => \N__45472\,
            lcout => \c0.FRAME_MATCHER_i_17\,
            ltout => OPEN,
            carryin => \bfn_19_18_0_\,
            carryout => \c0.n19459\,
            clk => \N__66760\,
            ce => 'H',
            sr => \N__45469\
        );

    \c0.add_49_19_THRU_CRY_0_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46641\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19459\,
            carryout => \c0.n19459_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_1_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46744\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19459_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19459_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_2_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46645\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19459_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19459_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_3_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46745\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19459_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19459_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_4_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46649\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19459_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19459_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_5_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46746\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19459_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19459_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_19_THRU_CRY_6_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46653\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19459_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19459_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i18_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51053\,
            in1 => \N__45569\,
            in2 => \_gnd_net_\,
            in3 => \N__45550\,
            lcout => \c0.FRAME_MATCHER_i_18\,
            ltout => OPEN,
            carryin => \bfn_19_19_0_\,
            carryout => \c0.n19460\,
            clk => \N__66772\,
            ce => 'H',
            sr => \N__45547\
        );

    \c0.add_49_20_THRU_CRY_0_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46628\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19460\,
            carryout => \c0.n19460_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_1_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46741\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19460_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19460_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_2_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46632\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19460_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19460_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_3_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46742\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19460_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19460_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_4_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46636\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19460_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19460_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_5_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46743\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19460_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19460_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_20_THRU_CRY_6_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46640\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19460_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19460_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i19_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51052\,
            in1 => \N__45524\,
            in2 => \_gnd_net_\,
            in3 => \N__45505\,
            lcout => \c0.FRAME_MATCHER_i_19\,
            ltout => OPEN,
            carryin => \bfn_19_20_0_\,
            carryout => \c0.n19461\,
            clk => \N__66786\,
            ce => 'H',
            sr => \N__45601\
        );

    \c0.add_49_21_THRU_CRY_0_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46495\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19461\,
            carryout => \c0.n19461_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_1_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46619\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19461_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19461_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_2_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46499\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19461_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19461_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_3_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46620\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19461_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19461_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_4_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46503\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19461_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19461_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_5_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46621\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19461_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19461_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_21_THRU_CRY_6_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46507\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19461_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19461_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i20_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51055\,
            in1 => \N__49992\,
            in2 => \_gnd_net_\,
            in3 => \N__45586\,
            lcout => \c0.FRAME_MATCHER_i_20\,
            ltout => OPEN,
            carryin => \bfn_19_21_0_\,
            carryout => \c0.n19462\,
            clk => \N__66797\,
            ce => 'H',
            sr => \N__49981\
        );

    \c0.add_49_22_THRU_CRY_0_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46545\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19462\,
            carryout => \c0.n19462_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_1_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46625\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19462_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19462_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_2_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46549\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19462_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19462_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_3_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46626\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19462_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19462_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_4_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46553\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19462_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19462_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_5_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46627\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19462_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19462_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_22_THRU_CRY_6_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46557\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19462_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19462_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i21_LC_19_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51010\,
            in1 => \N__45629\,
            in2 => \_gnd_net_\,
            in3 => \N__45613\,
            lcout => \c0.FRAME_MATCHER_i_21\,
            ltout => OPEN,
            carryin => \bfn_19_22_0_\,
            carryout => \c0.n19463\,
            clk => \N__66806\,
            ce => 'H',
            sr => \N__45610\
        );

    \c0.add_49_23_THRU_CRY_0_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46532\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19463\,
            carryout => \c0.n19463_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_1_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46622\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19463_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19463_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_2_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46536\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19463_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19463_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_3_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46623\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19463_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19463_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_4_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46540\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19463_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19463_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_5_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46624\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19463_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19463_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_23_THRU_CRY_6_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46544\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19463_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19463_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i22_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51088\,
            in1 => \N__45674\,
            in2 => \_gnd_net_\,
            in3 => \N__45655\,
            lcout => \c0.FRAME_MATCHER_i_22\,
            ltout => OPEN,
            carryin => \bfn_19_23_0_\,
            carryout => \c0.n19464\,
            clk => \N__66818\,
            ce => 'H',
            sr => \N__45652\
        );

    \c0.add_49_24_THRU_CRY_0_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46479\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19464\,
            carryout => \c0.n19464_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_1_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46616\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19464_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19464_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_2_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46483\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19464_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19464_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_3_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46617\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19464_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19464_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_4_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46487\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19464_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19464_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_5_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19464_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19464_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_24_THRU_CRY_6_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46491\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19464_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19464_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i23_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51087\,
            in1 => \N__45707\,
            in2 => \_gnd_net_\,
            in3 => \N__45688\,
            lcout => \c0.FRAME_MATCHER_i_23\,
            ltout => OPEN,
            carryin => \bfn_19_24_0_\,
            carryout => \c0.n19465\,
            clk => \N__66830\,
            ce => 'H',
            sr => \N__45685\
        );

    \c0.add_49_25_THRU_CRY_0_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46351\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19465\,
            carryout => \c0.n19465_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_1_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46492\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19465_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19465_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_2_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46355\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19465_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19465_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_3_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46493\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19465_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19465_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_4_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46359\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19465_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19465_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_5_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46494\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19465_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19465_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_25_THRU_CRY_6_LC_19_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46363\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19465_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19465_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i24_LC_19_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51085\,
            in1 => \N__45749\,
            in2 => \_gnd_net_\,
            in3 => \N__45730\,
            lcout => \c0.FRAME_MATCHER_i_24\,
            ltout => OPEN,
            carryin => \bfn_19_25_0_\,
            carryout => \c0.n19466\,
            clk => \N__66842\,
            ce => 'H',
            sr => \N__45727\
        );

    \c0.add_49_26_THRU_CRY_0_LC_19_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46269\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19466\,
            carryout => \c0.n19466_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_1_LC_19_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46273\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19466_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19466_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_2_LC_19_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46270\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19466_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19466_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_3_LC_19_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46274\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19466_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19466_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_4_LC_19_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46271\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19466_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19466_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_5_LC_19_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46275\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19466_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19466_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_26_THRU_CRY_6_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46272\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19466_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19466_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i25_LC_19_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51086\,
            in1 => \N__45791\,
            in2 => \_gnd_net_\,
            in3 => \N__45772\,
            lcout => \c0.FRAME_MATCHER_i_25\,
            ltout => OPEN,
            carryin => \bfn_19_26_0_\,
            carryout => \c0.n19467\,
            clk => \N__66851\,
            ce => 'H',
            sr => \N__45769\
        );

    \c0.add_49_27_THRU_CRY_0_LC_19_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46262\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19467\,
            carryout => \c0.n19467_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_1_LC_19_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46266\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19467_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19467_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_2_LC_19_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46263\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19467_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19467_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_3_LC_19_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46267\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19467_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19467_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_4_LC_19_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46264\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19467_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19467_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_5_LC_19_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46268\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19467_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19467_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_27_THRU_CRY_6_LC_19_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46265\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19467_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19467_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i26_LC_19_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51099\,
            in1 => \N__45830\,
            in2 => \_gnd_net_\,
            in3 => \N__45811\,
            lcout => \c0.FRAME_MATCHER_i_26\,
            ltout => OPEN,
            carryin => \bfn_19_27_0_\,
            carryout => \c0.n19468\,
            clk => \N__66860\,
            ce => 'H',
            sr => \N__45808\
        );

    \c0.add_49_28_THRU_CRY_0_LC_19_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46276\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19468\,
            carryout => \c0.n19468_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_1_LC_19_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46280\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19468_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19468_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_2_LC_19_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46277\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19468_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19468_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_3_LC_19_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46281\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19468_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19468_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_4_LC_19_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46278\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19468_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19468_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_5_LC_19_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46282\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19468_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19468_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_28_THRU_CRY_6_LC_19_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46279\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19468_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19468_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i27_LC_19_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51130\,
            in1 => \N__45869\,
            in2 => \_gnd_net_\,
            in3 => \N__45850\,
            lcout => \c0.FRAME_MATCHER_i_27\,
            ltout => OPEN,
            carryin => \bfn_19_28_0_\,
            carryout => \c0.n19469\,
            clk => \N__66866\,
            ce => 'H',
            sr => \N__45847\
        );

    \c0.add_49_29_THRU_CRY_0_LC_19_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46379\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19469\,
            carryout => \c0.n19469_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_1_LC_19_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46508\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19469_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19469_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_2_LC_19_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46383\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19469_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19469_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_3_LC_19_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46509\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19469_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19469_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_4_LC_19_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46387\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19469_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19469_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_5_LC_19_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__46510\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19469_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19469_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_29_THRU_CRY_6_LC_19_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46391\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19469_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19469_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i28_LC_19_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51123\,
            in1 => \N__50699\,
            in2 => \_gnd_net_\,
            in3 => \N__45907\,
            lcout => \c0.FRAME_MATCHER_i_28\,
            ltout => OPEN,
            carryin => \bfn_19_29_0_\,
            carryout => \c0.n19470\,
            clk => \N__66868\,
            ce => 'H',
            sr => \N__50455\
        );

    \c0.add_49_30_THRU_CRY_0_LC_19_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46511\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19470\,
            carryout => \c0.n19470_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_1_LC_19_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46515\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19470_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19470_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_2_LC_19_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46512\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19470_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19470_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_3_LC_19_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46516\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19470_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19470_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_4_LC_19_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46513\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19470_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19470_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_5_LC_19_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46517\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19470_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19470_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_30_THRU_CRY_6_LC_19_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46514\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19470_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19470_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i29_LC_19_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51131\,
            in1 => \N__45896\,
            in2 => \_gnd_net_\,
            in3 => \N__45880\,
            lcout => \c0.FRAME_MATCHER_i_29\,
            ltout => OPEN,
            carryin => \bfn_19_30_0_\,
            carryout => \c0.n19471\,
            clk => \N__66871\,
            ce => 'H',
            sr => \N__45955\
        );

    \c0.add_49_31_THRU_CRY_0_LC_19_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46518\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19471\,
            carryout => \c0.n19471_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_1_LC_19_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46522\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19471_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19471_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_2_LC_19_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46519\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19471_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19471_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_3_LC_19_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46523\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19471_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19471_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_4_LC_19_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46520\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19471_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19471_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_5_LC_19_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46524\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19471_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19471_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_31_THRU_CRY_6_LC_19_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46521\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19471_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19471_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i30_LC_19_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51161\,
            in1 => \N__45936\,
            in2 => \_gnd_net_\,
            in3 => \N__45922\,
            lcout => \c0.FRAME_MATCHER_i_30\,
            ltout => OPEN,
            carryin => \bfn_19_31_0_\,
            carryout => \c0.n19472\,
            clk => \N__66875\,
            ce => 'H',
            sr => \N__45919\
        );

    \c0.add_49_32_THRU_CRY_0_LC_19_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46525\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19472\,
            carryout => \c0.n19472_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_1_LC_19_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46529\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19472_THRU_CRY_0_THRU_CO\,
            carryout => \c0.n19472_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_2_LC_19_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46526\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19472_THRU_CRY_1_THRU_CO\,
            carryout => \c0.n19472_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_3_LC_19_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46530\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19472_THRU_CRY_2_THRU_CO\,
            carryout => \c0.n19472_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_4_LC_19_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46527\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19472_THRU_CRY_3_THRU_CO\,
            carryout => \c0.n19472_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_5_LC_19_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46531\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19472_THRU_CRY_4_THRU_CO\,
            carryout => \c0.n19472_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.add_49_32_THRU_CRY_6_LC_19_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46528\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \c0.n19472_THRU_CRY_5_THRU_CO\,
            carryout => \c0.n19472_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_i_i31_LC_19_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__51162\,
            in1 => \N__46109\,
            in2 => \_gnd_net_\,
            in3 => \N__46180\,
            lcout => \c0.FRAME_MATCHER_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66876\,
            ce => 'H',
            sr => \N__46075\
        );

    \c0.select_365_Select_1_i3_2_lut_4_lut_LC_20_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51472\,
            in1 => \N__51189\,
            in2 => \N__56544\,
            in3 => \N__50663\,
            lcout => \c0.n3_adj_4475\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_3_i3_2_lut_4_lut_LC_20_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51474\,
            in1 => \N__51159\,
            in2 => \N__46014\,
            in3 => \N__50662\,
            lcout => \c0.n3_adj_4472\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_2_i3_2_lut_4_lut_LC_20_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51473\,
            in1 => \N__51158\,
            in2 => \N__56403\,
            in3 => \N__50661\,
            lcout => \c0.n3_adj_4474\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_96_i9_2_lut_3_lut_LC_20_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__56568\,
            in1 => \N__56394\,
            in2 => \_gnd_net_\,
            in3 => \N__56708\,
            lcout => \c0.n9_adj_4302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_86_i9_2_lut_3_lut_LC_20_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__56569\,
            in1 => \_gnd_net_\,
            in2 => \N__56743\,
            in3 => \N__56419\,
            lcout => \c0.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_92_i11_2_lut_LC_20_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47384\,
            in2 => \_gnd_net_\,
            in3 => \N__47347\,
            lcout => \c0.n11_adj_4326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52105\,
            in1 => \N__52179\,
            in2 => \N__60154\,
            in3 => \N__52143\,
            lcout => \c0.n13697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1622_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__52144\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48451\,
            lcout => \c0.n10_adj_4399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1312_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48401\,
            in2 => \_gnd_net_\,
            in3 => \N__47253\,
            lcout => \c0.n6_adj_4258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i60_LC_20_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__60889\,
            in1 => \N__68568\,
            in2 => \N__52275\,
            in3 => \N__64879\,
            lcout => \c0.data_in_frame_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1258_LC_20_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54193\,
            in2 => \_gnd_net_\,
            in3 => \N__60191\,
            lcout => \c0.n6_adj_4241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i71_LC_20_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__62509\,
            in1 => \N__52106\,
            in2 => \N__66028\,
            in3 => \N__65648\,
            lcout => \c0.data_in_frame_8_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i70_LC_20_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__67186\,
            in1 => \N__66008\,
            in2 => \N__48410\,
            in3 => \N__62510\,
            lcout => \c0.data_in_frame_8_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i88_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62374\,
            in1 => \N__69064\,
            in2 => \N__49753\,
            in3 => \N__68954\,
            lcout => \c0.data_in_frame_10_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i87_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69063\,
            in1 => \N__65576\,
            in2 => \N__60094\,
            in3 => \N__62376\,
            lcout => \c0.data_in_frame_10_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1316_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60081\,
            in2 => \_gnd_net_\,
            in3 => \N__49736\,
            lcout => \c0.n21925\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1666_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47548\,
            in1 => \N__51753\,
            in2 => \N__47524\,
            in3 => \N__51700\,
            lcout => \c0.n6_adj_4395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i22_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__67219\,
            in1 => \N__60888\,
            in2 => \N__48204\,
            in3 => \N__69065\,
            lcout => \c0.data_in_frame_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i82_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69062\,
            in1 => \N__62375\,
            in2 => \N__51547\,
            in3 => \N__63862\,
            lcout => \c0.data_in_frame_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1311_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__52098\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57712\,
            lcout => OPEN,
            ltout => \c0.n21861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1313_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47455\,
            in1 => \N__52206\,
            in2 => \N__47422\,
            in3 => \N__47419\,
            lcout => \c0.n21940\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__50439\,
            in1 => \N__51622\,
            in2 => \_gnd_net_\,
            in3 => \N__51567\,
            lcout => OPEN,
            ltout => \c0.n8_adj_4254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1290_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52274\,
            in1 => \N__47827\,
            in2 => \N__47809\,
            in3 => \N__47806\,
            lcout => \c0.n13865\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i46_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__60881\,
            in1 => \N__62148\,
            in2 => \N__47787\,
            in3 => \N__67217\,
            lcout => \c0.data_in_frame_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1614_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__47766\,
            in1 => \N__47737\,
            in2 => \N__47688\,
            in3 => \N__47707\,
            lcout => \c0.n12484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i10_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69806\,
            in1 => \N__60882\,
            in2 => \N__47689\,
            in3 => \N__63849\,
            lcout => data_in_frame_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i72_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66020\,
            in1 => \N__62542\,
            in2 => \N__57731\,
            in3 => \N__68988\,
            lcout => \c0.data_in_frame_8_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i6_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__67216\,
            in1 => \N__60883\,
            in2 => \N__51773\,
            in3 => \N__66021\,
            lcout => \c0.data_in_frame_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1662_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50341\,
            in1 => \N__48197\,
            in2 => \N__48170\,
            in3 => \N__47640\,
            lcout => OPEN,
            ltout => \c0.n13848_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1630_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010110"
        )
    port map (
            in0 => \N__47968\,
            in1 => \N__47578\,
            in2 => \N__47566\,
            in3 => \N__51970\,
            lcout => \c0.n13_adj_4405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1310_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__48233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47949\,
            lcout => \c0.n13652\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1667_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__48196\,
            in1 => \N__48158\,
            in2 => \_gnd_net_\,
            in3 => \N__50340\,
            lcout => \c0.n13398\,
            ltout => \c0.n13398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1717_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48048\,
            in1 => \N__48001\,
            in2 => \N__47971\,
            in3 => \N__47967\,
            lcout => \c0.n21794\,
            ltout => \c0.n21794_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1824_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47938\,
            in2 => \N__47911\,
            in3 => \N__48232\,
            lcout => \c0.n22239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51508\,
            in1 => \N__48364\,
            in2 => \N__52291\,
            in3 => \N__48340\,
            lcout => \c0.n44_adj_4262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i64_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__68989\,
            in1 => \N__68569\,
            in2 => \N__51919\,
            in3 => \N__60897\,
            lcout => \c0.data_in_frame_7_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1905_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__47902\,
            in1 => \N__51974\,
            in2 => \_gnd_net_\,
            in3 => \N__48351\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1308_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51914\,
            in1 => \N__48279\,
            in2 => \N__47848\,
            in3 => \N__47845\,
            lcout => \c0.n13771\,
            ltout => \c0.n13771_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1314_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48355\,
            in3 => \N__54999\,
            lcout => \c0.n4\,
            ltout => \c0.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48352\,
            in1 => \N__48383\,
            in2 => \N__48343\,
            in3 => \N__60054\,
            lcout => \c0.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1220_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__52443\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60435\,
            lcout => \c0.n21967\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1300_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48334\,
            in1 => \N__48384\,
            in2 => \N__48322\,
            in3 => \N__48292\,
            lcout => \c0.n13425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1402_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61468\,
            in1 => \N__54175\,
            in2 => \N__54478\,
            in3 => \N__48286\,
            lcout => \c0.n21170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i84_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__64836\,
            in1 => \N__62543\,
            in2 => \N__69191\,
            in3 => \N__48280\,
            lcout => \c0.data_in_frame_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66691\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1252_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48414\,
            in1 => \N__60367\,
            in2 => \N__48271\,
            in3 => \N__51856\,
            lcout => \c0.n21979\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1302_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48448\,
            in2 => \_gnd_net_\,
            in3 => \N__52171\,
            lcout => \c0.n21964\,
            ltout => \c0.n21964_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_adj_1320_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60973\,
            in1 => \N__48262\,
            in2 => \N__48244\,
            in3 => \N__48240\,
            lcout => \c0.n40_adj_4261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1259_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49755\,
            in1 => \N__49779\,
            in2 => \N__48466\,
            in3 => \N__63969\,
            lcout => \c0.n21864\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1328_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__48449\,
            in1 => \N__60520\,
            in2 => \N__48415\,
            in3 => \N__49754\,
            lcout => \c0.n22415\,
            ltout => \c0.n22415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1833_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__52107\,
            in1 => \_gnd_net_\,
            in2 => \N__48388\,
            in3 => \N__57730\,
            lcout => \c0.n6_adj_4256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i73_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69750\,
            in1 => \N__62554\,
            in2 => \N__52207\,
            in3 => \N__69557\,
            lcout => \c0.data_in_frame_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66705\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1275_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61807\,
            in2 => \_gnd_net_\,
            in3 => \N__55326\,
            lcout => \c0.n13681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i61_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__63205\,
            in1 => \N__50438\,
            in2 => \N__60887\,
            in3 => \N__68674\,
            lcout => \c0.data_in_frame_7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1841_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__61813\,
            in1 => \N__55327\,
            in2 => \_gnd_net_\,
            in3 => \N__57490\,
            lcout => \c0.n22355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i135_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__52375\,
            in1 => \N__68095\,
            in2 => \N__66019\,
            in3 => \N__65661\,
            lcout => \c0.data_in_frame_16_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i86_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69125\,
            in1 => \N__62396\,
            in2 => \N__48385\,
            in3 => \N__67163\,
            lcout => \c0.data_in_frame_10_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66719\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_3_lut_4_lut_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52534\,
            in1 => \N__54709\,
            in2 => \N__54893\,
            in3 => \N__54561\,
            lcout => \c0.n35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i142_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69695\,
            in1 => \N__68092\,
            in2 => \N__55338\,
            in3 => \N__67162\,
            lcout => \c0.data_in_frame_17_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i77_LC_20_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__63143\,
            in1 => \N__69697\,
            in2 => \N__52480\,
            in3 => \N__62430\,
            lcout => \c0.data_in_frame_9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1263_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52476\,
            in2 => \_gnd_net_\,
            in3 => \N__57643\,
            lcout => \c0.n6_adj_4243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i143_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__68091\,
            in1 => \N__69696\,
            in2 => \N__61823\,
            in3 => \N__65563\,
            lcout => \c0.data_in_frame_17_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i53_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49708\,
            in1 => \N__63144\,
            in2 => \_gnd_net_\,
            in3 => \N__49608\,
            lcout => data_in_frame_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1584_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__49654\,
            in1 => \N__49641\,
            in2 => \N__49609\,
            in3 => \N__49589\,
            lcout => \c0.n13605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i35_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68373\,
            in1 => \N__64518\,
            in2 => \N__49596\,
            in3 => \N__60727\,
            lcout => \c0.data_in_frame_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_out_frame_6__6__5471_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__49356\,
            in1 => \N__49012\,
            in2 => \N__48571\,
            in3 => \N__48480\,
            lcout => data_out_frame_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1329_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60399\,
            in2 => \_gnd_net_\,
            in3 => \N__60196\,
            lcout => OPEN,
            ltout => \c0.n22440_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1235_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52629\,
            in1 => \N__49783\,
            in2 => \N__49762\,
            in3 => \N__52608\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4229_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1860_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60101\,
            in1 => \N__49759\,
            in2 => \N__49720\,
            in3 => \N__55015\,
            lcout => \c0.n5943\,
            ltout => \c0.n5943_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1754_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55328\,
            in1 => \N__55217\,
            in2 => \N__49717\,
            in3 => \N__55303\,
            lcout => \c0.n22081\,
            ltout => \c0.n22081_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1273_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__61615\,
            in1 => \_gnd_net_\,
            in2 => \N__49714\,
            in3 => \N__55395\,
            lcout => \c0.n13457\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1894_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55396\,
            in1 => \N__61616\,
            in2 => \N__61216\,
            in3 => \N__53218\,
            lcout => \c0.n13443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1221_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52378\,
            in1 => \N__55126\,
            in2 => \_gnd_net_\,
            in3 => \N__52348\,
            lcout => \c0.n21187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1580_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55624\,
            in1 => \N__63356\,
            in2 => \N__64030\,
            in3 => \N__61603\,
            lcout => \c0.n22349\,
            ltout => \c0.n22349_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1616_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57446\,
            in1 => \N__61420\,
            in2 => \N__49711\,
            in3 => \N__55431\,
            lcout => \c0.n6_adj_4224\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1857_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55430\,
            in1 => \N__61415\,
            in2 => \_gnd_net_\,
            in3 => \N__57445\,
            lcout => OPEN,
            ltout => \c0.n21858_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1247_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55385\,
            in1 => \N__64017\,
            in2 => \N__49900\,
            in3 => \N__55623\,
            lcout => \c0.n21989\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i159_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__68007\,
            in1 => \N__67339\,
            in2 => \N__61617\,
            in3 => \N__65568\,
            lcout => \c0.data_in_frame_19_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i215_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__65567\,
            in1 => \N__69249\,
            in2 => \N__59439\,
            in3 => \N__67677\,
            lcout => \c0.data_in_frame_26_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i139_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__68006\,
            in1 => \N__69802\,
            in2 => \N__68436\,
            in3 => \N__61416\,
            lcout => \c0.data_in_frame_17_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i138_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69801\,
            in1 => \N__68008\,
            in2 => \N__64035\,
            in3 => \N__63764\,
            lcout => \c0.data_in_frame_17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1567_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50710\,
            in1 => \N__49890\,
            in2 => \N__50010\,
            in3 => \N__49857\,
            lcout => \c0.n16_adj_4375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_13_i3_2_lut_4_lut_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51433\,
            in1 => \N__51041\,
            in2 => \N__49861\,
            in3 => \N__50609\,
            lcout => \c0.n3_adj_4454\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i172_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62184\,
            in1 => \N__68067\,
            in2 => \N__49939\,
            in3 => \N__64871\,
            lcout => \c0.data_in_frame_21_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66773\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1211_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__63486\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65248\,
            lcout => \c0.n22028\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_15_i3_2_lut_4_lut_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__50610\,
            in1 => \N__49821\,
            in2 => \N__51111\,
            in3 => \N__51435\,
            lcout => \c0.n3_adj_4452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i185_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__68065\,
            in1 => \N__68670\,
            in2 => \N__63268\,
            in3 => \N__69503\,
            lcout => \c0.data_in_frame_23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66773\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i171_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62183\,
            in1 => \N__68066\,
            in2 => \N__53818\,
            in3 => \N__68369\,
            lcout => \c0.data_in_frame_21_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66773\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_20_i3_2_lut_4_lut_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51434\,
            in1 => \N__51042\,
            in2 => \N__50011\,
            in3 => \N__50611\,
            lcout => \c0.n3_adj_4442\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1369_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53602\,
            in1 => \N__65322\,
            in2 => \N__49969\,
            in3 => \N__53788\,
            lcout => \c0.n12_adj_4290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1214_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53809\,
            in2 => \_gnd_net_\,
            in3 => \N__49934\,
            lcout => \c0.n21870\,
            ltout => \c0.n21870_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1192_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50073\,
            in1 => \N__55486\,
            in2 => \N__49942\,
            in3 => \N__55540\,
            lcout => \c0.n13761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1350_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55919\,
            in1 => \N__50072\,
            in2 => \_gnd_net_\,
            in3 => \N__49920\,
            lcout => \c0.n22396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__49935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49921\,
            lcout => \c0.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i207_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69730\,
            in1 => \N__65573\,
            in2 => \N__58610\,
            in3 => \N__67707\,
            lcout => \c0.data_in_frame_25_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i191_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__65572\,
            in1 => \N__55920\,
            in2 => \N__68679\,
            in3 => \N__68069\,
            lcout => \c0.data_in_frame_23_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i189_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__68068\,
            in1 => \N__68669\,
            in2 => \N__63172\,
            in3 => \N__50074\,
            lcout => \c0.data_in_frame_23_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1195_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__53601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53728\,
            lcout => \c0.n13266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1363_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__56059\,
            in1 => \N__54135\,
            in2 => \N__53941\,
            in3 => \N__59023\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1384_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011101101"
        )
    port map (
            in0 => \N__50204\,
            in1 => \N__50017\,
            in2 => \N__50062\,
            in3 => \N__56326\,
            lcout => \c0.n22_adj_4298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i157_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__63058\,
            in1 => \N__68070\,
            in2 => \N__67402\,
            in3 => \N__55876\,
            lcout => \c0.data_in_frame_19_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_adj_1721_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53600\,
            in2 => \_gnd_net_\,
            in3 => \N__54007\,
            lcout => \c0.n10_adj_4483\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1899_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__53654\,
            in1 => \N__53979\,
            in2 => \N__66913\,
            in3 => \N__53767\,
            lcout => \c0.n21233\,
            ltout => \c0.n21233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1364_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__50047\,
            in1 => \N__50038\,
            in2 => \N__50020\,
            in3 => \N__53986\,
            lcout => \c0.n23506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i239_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__65562\,
            in1 => \N__54112\,
            in2 => \N__62202\,
            in3 => \N__67708\,
            lcout => \c0.data_in_frame_29_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1727_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50206\,
            in1 => \N__58770\,
            in2 => \N__65103\,
            in3 => \N__59419\,
            lcout => \c0.n45_adj_4486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i158_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__68140\,
            in1 => \N__67392\,
            in2 => \N__58835\,
            in3 => \N__67218\,
            lcout => \c0.data_in_frame_19_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.select_365_Select_10_i3_2_lut_4_lut_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51436\,
            in1 => \N__51069\,
            in2 => \N__50167\,
            in3 => \N__50620\,
            lcout => \c0.n3_adj_4460\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i155_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__68139\,
            in1 => \N__67391\,
            in2 => \N__56006\,
            in3 => \N__68412\,
            lcout => \c0.data_in_frame_19_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i1_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__63643\,
            in1 => \N__50106\,
            in2 => \N__59716\,
            in3 => \N__56207\,
            lcout => rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i221_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__67348\,
            in1 => \N__63092\,
            in2 => \N__55839\,
            in3 => \N__67752\,
            lcout => \c0.data_in_frame_27_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__50229\,
            in1 => \N__50259\,
            in2 => \_gnd_net_\,
            in3 => \N__50244\,
            lcout => \c0.rx.n18655\,
            ltout => \c0.rx.n18655_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i3_4_lut_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__54261\,
            in1 => \N__54284\,
            in2 => \N__50080\,
            in3 => \N__54321\,
            lcout => \c0.rx.n21704\,
            ltout => \c0.rx.n21704_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i18882_2_lut_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50077\,
            in3 => \N__59711\,
            lcout => OPEN,
            ltout => \c0.rx.n22573_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i25_4_lut_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011111001100"
        )
    port map (
            in0 => \N__57059\,
            in1 => \N__56898\,
            in2 => \N__50269\,
            in3 => \N__56835\,
            lcout => OPEN,
            ltout => \c0.rx.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i1_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50266\,
            in3 => \N__57003\,
            lcout => \r_SM_Main_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Clock_Count__i0_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54285\,
            in2 => \_gnd_net_\,
            in3 => \N__50263\,
            lcout => \c0.rx.r_Clock_Count_0\,
            ltout => OPEN,
            carryin => \bfn_20_24_0_\,
            carryout => \c0.rx.n19533\,
            clk => \N__66843\,
            ce => \N__51499\,
            sr => \N__51484\
        );

    \c0.rx.r_Clock_Count__i1_LC_20_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50260\,
            in2 => \_gnd_net_\,
            in3 => \N__50248\,
            lcout => \c0.rx.r_Clock_Count_1\,
            ltout => OPEN,
            carryin => \c0.rx.n19533\,
            carryout => \c0.rx.n19534\,
            clk => \N__66843\,
            ce => \N__51499\,
            sr => \N__51484\
        );

    \c0.rx.r_Clock_Count__i2_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50245\,
            in2 => \_gnd_net_\,
            in3 => \N__50233\,
            lcout => \c0.rx.r_Clock_Count_2\,
            ltout => OPEN,
            carryin => \c0.rx.n19534\,
            carryout => \c0.rx.n19535\,
            clk => \N__66843\,
            ce => \N__51499\,
            sr => \N__51484\
        );

    \c0.rx.r_Clock_Count__i3_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50230\,
            in2 => \_gnd_net_\,
            in3 => \N__50218\,
            lcout => \c0.rx.r_Clock_Count_3\,
            ltout => OPEN,
            carryin => \c0.rx.n19535\,
            carryout => \c0.rx.n19536\,
            clk => \N__66843\,
            ce => \N__51499\,
            sr => \N__51484\
        );

    \c0.rx.r_Clock_Count__i4_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54322\,
            in2 => \_gnd_net_\,
            in3 => \N__50215\,
            lcout => \c0.rx.r_Clock_Count_4\,
            ltout => OPEN,
            carryin => \c0.rx.n19536\,
            carryout => \c0.rx.n19537\,
            clk => \N__66843\,
            ce => \N__51499\,
            sr => \N__51484\
        );

    \c0.rx.r_Clock_Count__i5_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54043\,
            in2 => \_gnd_net_\,
            in3 => \N__50212\,
            lcout => \c0.rx.r_Clock_Count_5\,
            ltout => OPEN,
            carryin => \c0.rx.n19537\,
            carryout => \c0.rx.n19538\,
            clk => \N__66843\,
            ce => \N__51499\,
            sr => \N__51484\
        );

    \c0.rx.r_Clock_Count__i6_LC_20_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54031\,
            in2 => \_gnd_net_\,
            in3 => \N__50209\,
            lcout => \c0.rx.r_Clock_Count_6\,
            ltout => OPEN,
            carryin => \c0.rx.n19538\,
            carryout => \c0.rx.n19539\,
            clk => \N__66843\,
            ce => \N__51499\,
            sr => \N__51484\
        );

    \c0.rx.r_Clock_Count__i7_LC_20_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54055\,
            in2 => \_gnd_net_\,
            in3 => \N__51502\,
            lcout => \c0.rx.r_Clock_Count_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66843\,
            ce => \N__51499\,
            sr => \N__51484\
        );

    \c0.select_365_Select_28_i3_2_lut_4_lut_LC_20_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__51466\,
            in1 => \N__51098\,
            in2 => \N__50709\,
            in3 => \N__50621\,
            lcout => \c0.n3_adj_4430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1617_LC_21_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__51623\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51571\,
            lcout => \c0.n13555\,
            ltout => \c0.n13555_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1285_LC_21_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52510\,
            in1 => \N__50443\,
            in2 => \N__50416\,
            in3 => \N__52229\,
            lcout => \c0.n22043\,
            ltout => \c0.n22043_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1837_LC_21_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50403\,
            in1 => \N__51596\,
            in2 => \N__50392\,
            in3 => \N__54683\,
            lcout => \c0.n21097\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_87_i9_2_lut_3_lut_LC_21_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__56729\,
            in1 => \N__56582\,
            in2 => \_gnd_net_\,
            in3 => \N__56455\,
            lcout => \c0.n9_adj_4341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i33_LC_21_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64549\,
            in1 => \N__60892\,
            in2 => \N__54436\,
            in3 => \N__69568\,
            lcout => \c0.data_in_frame_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66669\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i62_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__60891\,
            in1 => \N__67142\,
            in2 => \N__51598\,
            in3 => \N__68600\,
            lcout => \c0.data_in_frame_7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66669\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__50389\,
            in1 => \N__50349\,
            in2 => \N__50281\,
            in3 => \N__51754\,
            lcout => \c0.n13488\,
            ltout => \c0.n13488_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_adj_1321_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51820\,
            in1 => \N__51592\,
            in2 => \N__51805\,
            in3 => \N__51802\,
            lcout => \c0.n39_adj_4263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i44_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__60890\,
            in1 => \N__62088\,
            in2 => \N__51630\,
            in3 => \N__64888\,
            lcout => \c0.data_in_frame_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66669\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20132_2_lut_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51755\,
            in2 => \_gnd_net_\,
            in3 => \N__51710\,
            lcout => \c0.n23827\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1821_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51631\,
            in1 => \N__54682\,
            in2 => \N__51597\,
            in3 => \N__51566\,
            lcout => OPEN,
            ltout => \c0.n20368_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1745_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51997\,
            in1 => \N__52006\,
            in2 => \N__51550\,
            in3 => \N__51837\,
            lcout => \c0.n22133\,
            ltout => \c0.n22133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1315_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57369\,
            in1 => \N__51543\,
            in2 => \N__51526\,
            in3 => \N__51892\,
            lcout => \c0.n20927\,
            ltout => \c0.n20927_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1319_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__51523\,
            in1 => \N__52330\,
            in2 => \N__51517\,
            in3 => \N__51514\,
            lcout => \c0.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1317_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__54777\,
            in1 => \_gnd_net_\,
            in2 => \N__51918\,
            in3 => \_gnd_net_\,
            lcout => \c0.n22379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1555_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52050\,
            in2 => \_gnd_net_\,
            in3 => \N__54399\,
            lcout => \c0.n22334\,
            ltout => \c0.n22334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_1408_i15_2_lut_3_lut_LC_21_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51836\,
            in2 => \N__52000\,
            in3 => \N__51996\,
            lcout => \c0.n15_adj_4404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1809_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51943\,
            in1 => \N__51910\,
            in2 => \_gnd_net_\,
            in3 => \N__54776\,
            lcout => \c0.n6_adj_4259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1296_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__51855\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54214\,
            lcout => \c0.n22270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1318_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59244\,
            in2 => \_gnd_net_\,
            in3 => \N__57889\,
            lcout => \c0.n22060\,
            ltout => \c0.n22060_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1323_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__51886\,
            in1 => \N__51877\,
            in2 => \N__51868\,
            in3 => \N__51865\,
            lcout => OPEN,
            ltout => \c0.n11_adj_4266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1324_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54588\,
            in1 => \N__57655\,
            in2 => \N__51859\,
            in3 => \N__51854\,
            lcout => OPEN,
            ltout => \c0.n22842_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1326_LC_21_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__60363\,
            in1 => \N__52309\,
            in2 => \N__51841\,
            in3 => \N__52596\,
            lcout => \c0.n15_adj_4269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i47_LC_21_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__65689\,
            in1 => \N__51838\,
            in2 => \N__62177\,
            in3 => \N__60807\,
            lcout => \c0.data_in_frame_5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1298_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59579\,
            in2 => \_gnd_net_\,
            in3 => \N__57581\,
            lcout => \c0.n22245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_4_lut_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52461\,
            in1 => \N__52132\,
            in2 => \N__52303\,
            in3 => \N__52505\,
            lcout => \c0.n38_adj_4260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1294_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61062\,
            in1 => \N__52282\,
            in2 => \N__57619\,
            in3 => \N__54601\,
            lcout => \c0.n5810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1332_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52276\,
            in2 => \_gnd_net_\,
            in3 => \N__52233\,
            lcout => \c0.n22139\,
            ltout => \c0.n22139_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1336_LC_21_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54859\,
            in1 => \N__52462\,
            in2 => \N__52210\,
            in3 => \N__61024\,
            lcout => \c0.n20135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1339_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52133\,
            in1 => \N__54894\,
            in2 => \N__52329\,
            in3 => \N__57732\,
            lcout => \c0.n10_adj_4274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1230_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52202\,
            in1 => \N__52178\,
            in2 => \_gnd_net_\,
            in3 => \N__52134\,
            lcout => \c0.n21822\,
            ltout => \c0.n21822_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1292_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57615\,
            in1 => \N__52111\,
            in2 => \N__52072\,
            in3 => \N__54600\,
            lcout => \c0.n22221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1239_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__52377\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52344\,
            lcout => \c0.n22242\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1397_LC_21_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__54174\,
            in1 => \_gnd_net_\,
            in2 => \N__61501\,
            in3 => \N__54477\,
            lcout => \c0.n22296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1261_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52426\,
            in1 => \N__57346\,
            in2 => \N__57244\,
            in3 => \N__61496\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1907_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52535\,
            in1 => \N__54710\,
            in2 => \N__52411\,
            in3 => \N__52408\,
            lcout => \c0.n13786\,
            ltout => \c0.n13786_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_4_lut_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__52376\,
            in1 => \N__57285\,
            in2 => \N__52351\,
            in3 => \N__52343\,
            lcout => \c0.n7_adj_4235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i184_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__60310\,
            in1 => \N__68987\,
            in2 => \_gnd_net_\,
            in3 => \N__59199\,
            lcout => data_in_frame_22_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i74_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69839\,
            in1 => \N__63779\,
            in2 => \N__54633\,
            in3 => \N__62501\,
            lcout => \c0.data_in_frame_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1337_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60007\,
            in2 => \_gnd_net_\,
            in3 => \N__54626\,
            lcout => \c0.n13974\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i58_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__68672\,
            in1 => \N__60806\,
            in2 => \N__54895\,
            in3 => \N__63800\,
            lcout => \c0.data_in_frame_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1873_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55102\,
            in1 => \N__55064\,
            in2 => \_gnd_net_\,
            in3 => \N__54500\,
            lcout => \c0.n6_adj_4221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i81_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__69480\,
            in1 => \N__62498\,
            in2 => \N__69192\,
            in3 => \N__54714\,
            lcout => \c0.data_in_frame_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i121_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__62496\,
            in1 => \N__68673\,
            in2 => \N__54507\,
            in3 => \N__69481\,
            lcout => \c0.data_in_frame_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i83_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__68356\,
            in1 => \N__62499\,
            in2 => \N__69193\,
            in3 => \N__52539\,
            lcout => \c0.data_in_frame_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1854_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58162\,
            in1 => \N__55118\,
            in2 => \_gnd_net_\,
            in3 => \N__57291\,
            lcout => \c0.n20402\,
            ltout => \c0.n20402_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1898_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57292\,
            in1 => \N__57325\,
            in2 => \N__52513\,
            in3 => \N__58216\,
            lcout => \c0.n21834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i79_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62497\,
            in1 => \N__69883\,
            in2 => \N__52509\,
            in3 => \N__65670\,
            lcout => \c0.data_in_frame_9_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66734\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1333_LC_21_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52475\,
            in2 => \_gnd_net_\,
            in3 => \N__57395\,
            lcout => \c0.n21873\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1720_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__53656\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53695\,
            lcout => \c0.n22119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65761\,
            in1 => \N__52450\,
            in2 => \N__55027\,
            in3 => \N__60400\,
            lcout => OPEN,
            ltout => \c0.n18_adj_4222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52633\,
            in1 => \N__55668\,
            in2 => \N__52612\,
            in3 => \N__60103\,
            lcout => \c0.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i102_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64451\,
            in1 => \N__62428\,
            in2 => \N__60948\,
            in3 => \N__67171\,
            lcout => \c0.data_in_frame_12_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i76_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__62427\,
            in1 => \N__57396\,
            in2 => \N__69877\,
            in3 => \N__64825\,
            lcout => \c0.data_in_frame_9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i122_LC_21_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__63780\,
            in1 => \N__62429\,
            in2 => \N__68658\,
            in3 => \N__61382\,
            lcout => \c0.data_in_frame_15_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1217_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54796\,
            in1 => \N__52609\,
            in2 => \N__61360\,
            in3 => \N__52585\,
            lcout => \c0.n22003\,
            ltout => \c0.n22003_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1215_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__52576\,
            in1 => \N__55210\,
            in2 => \N__52564\,
            in3 => \N__52561\,
            lcout => \c0.n6221\,
            ltout => \c0.n6221_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1216_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52555\,
            in3 => \N__55895\,
            lcout => \c0.n22084\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i150_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__68093\,
            in1 => \N__69124\,
            in2 => \N__61579\,
            in3 => \N__67122\,
            lcout => \c0.data_in_frame_18_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66762\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i169_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62150\,
            in1 => \N__68094\,
            in2 => \N__55728\,
            in3 => \N__69537\,
            lcout => \c0.data_in_frame_21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66762\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1892_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55626\,
            in1 => \N__55557\,
            in2 => \N__64034\,
            in3 => \N__52552\,
            lcout => \c0.n22311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1866_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58838\,
            in1 => \N__58691\,
            in2 => \_gnd_net_\,
            in3 => \N__59278\,
            lcout => \c0.n22099\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i205_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__63107\,
            in1 => \N__53719\,
            in2 => \N__69882\,
            in3 => \N__67675\,
            lcout => \c0.data_in_frame_25_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66774\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1861_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54951\,
            in1 => \N__61747\,
            in2 => \_gnd_net_\,
            in3 => \N__58543\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4226_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1231_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53242\,
            in1 => \N__55156\,
            in2 => \N__53227\,
            in3 => \N__63357\,
            lcout => \c0.n23615\,
            ltout => \c0.n23615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1232_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__53224\,
            in3 => \N__65073\,
            lcout => \c0.n22100\,
            ltout => \c0.n22100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1278_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58278\,
            in1 => \N__53286\,
            in2 => \N__53221\,
            in3 => \N__53901\,
            lcout => \c0.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1226_LC_21_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53217\,
            in1 => \N__55155\,
            in2 => \N__53206\,
            in3 => \N__58542\,
            lcout => \c0.n12594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1767_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__52649\,
            in1 => \N__53196\,
            in2 => \_gnd_net_\,
            in3 => \N__53029\,
            lcout => \c0.n21366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.FRAME_MATCHER_state_i20_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52650\,
            in2 => \_gnd_net_\,
            in3 => \N__52867\,
            lcout => \c0.FRAME_MATCHER_state_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66788\,
            ce => 'H',
            sr => \N__53518\
        );

    \c0.i2_3_lut_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__53810\,
            in1 => \N__53786\,
            in2 => \_gnd_net_\,
            in3 => \N__55535\,
            lcout => \c0.n21043\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1455_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__53503\,
            in1 => \N__53475\,
            in2 => \_gnd_net_\,
            in3 => \N__53416\,
            lcout => \c0.n13379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55228\,
            in1 => \N__53862\,
            in2 => \N__53335\,
            in3 => \N__55753\,
            lcout => OPEN,
            ltout => \c0.n28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i16_4_lut_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62839\,
            in1 => \N__55261\,
            in2 => \N__53302\,
            in3 => \N__55678\,
            lcout => \c0.n23640\,
            ltout => \c0.n23640_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1903_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__60489\,
            in1 => \_gnd_net_\,
            in2 => \N__53299\,
            in3 => \N__53292\,
            lcout => \c0.n22197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__55485\,
            in1 => \N__53256\,
            in2 => \N__57972\,
            in3 => \N__55684\,
            lcout => \c0.n22305\,
            ltout => \c0.n22305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1901_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60340\,
            in2 => \N__53296\,
            in3 => \N__60312\,
            lcout => \c0.n20137\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__53293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53257\,
            lcout => \c0.n21208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1200_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53848\,
            in2 => \_gnd_net_\,
            in3 => \N__53248\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1201_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60313\,
            in1 => \N__63257\,
            in2 => \N__53821\,
            in3 => \N__64257\,
            lcout => \c0.n21160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1902_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__53817\,
            in1 => \N__53787\,
            in2 => \N__53727\,
            in3 => \N__55539\,
            lcout => \c0.n21949\,
            ltout => \c0.n21949_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1191_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__53650\,
            in1 => \_gnd_net_\,
            in2 => \N__53770\,
            in3 => \N__53762\,
            lcout => \c0.n23009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1736_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53690\,
            in1 => \N__59541\,
            in2 => \N__53766\,
            in3 => \N__64189\,
            lcout => \c0.n22157\,
            ltout => \c0.n22157_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1733_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58899\,
            in1 => \N__55807\,
            in2 => \N__53746\,
            in3 => \N__54130\,
            lcout => \c0.n20846\,
            ltout => \c0.n20846_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1734_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__54131\,
            in1 => \N__54008\,
            in2 => \N__53731\,
            in3 => \N__55794\,
            lcout => \c0.n12_adj_4491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1655_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53720\,
            in1 => \N__53689\,
            in2 => \N__53655\,
            in3 => \N__53599\,
            lcout => \c0.n22370\,
            ltout => \c0.n22370_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1735_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53548\,
            in1 => \N__53542\,
            in2 => \N__53536\,
            in3 => \N__56080\,
            lcout => \c0.n23356\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1194_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__53827\,
            in1 => \N__66097\,
            in2 => \_gnd_net_\,
            in3 => \N__54015\,
            lcout => \c0.n22145\,
            ltout => \c0.n22145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1381_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58614\,
            in1 => \N__53980\,
            in2 => \N__53968\,
            in3 => \N__66135\,
            lcout => \c0.n10_adj_4297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i238_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67705\,
            in1 => \N__62167\,
            in2 => \N__56308\,
            in3 => \N__67079\,
            lcout => \c0.data_in_frame_29_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1383_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59542\,
            in1 => \N__64588\,
            in2 => \N__59365\,
            in3 => \N__56065\,
            lcout => OPEN,
            ltout => \c0.n23335_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1387_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111110011111"
        )
    port map (
            in0 => \N__53916\,
            in1 => \N__53965\,
            in2 => \N__53959\,
            in3 => \N__58717\,
            lcout => \c0.n21_adj_4300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i236_LC_21_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__62166\,
            in1 => \N__64887\,
            in2 => \N__53940\,
            in3 => \N__67706\,
            lcout => \c0.data_in_frame_29_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i225_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67751\,
            in1 => \N__64565\,
            in2 => \N__53920\,
            in3 => \N__69538\,
            lcout => \c0.data_in_frame_28_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1196_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__53905\,
            in1 => \N__65428\,
            in2 => \N__55729\,
            in3 => \N__53866\,
            lcout => \c0.n22040\,
            ltout => \c0.n22040_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1193_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67818\,
            in1 => \N__64228\,
            in2 => \N__53839\,
            in3 => \N__53836\,
            lcout => \c0.n21099\,
            ltout => \c0.n21099_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1718_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54148\,
            in1 => \N__55829\,
            in2 => \N__54139\,
            in3 => \N__54136\,
            lcout => \c0.n22148\,
            ltout => \c0.n22148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1377_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111011110"
        )
    port map (
            in0 => \N__54111\,
            in1 => \N__54097\,
            in2 => \N__54079\,
            in3 => \N__54076\,
            lcout => \c0.n26_adj_4294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i173_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62160\,
            in1 => \N__68141\,
            in2 => \N__58337\,
            in3 => \N__63000\,
            lcout => \c0.data_in_frame_21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_1178_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59749\,
            in2 => \_gnd_net_\,
            in3 => \N__56160\,
            lcout => n12977,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_3_lut_4_lut_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__56991\,
            in1 => \N__56808\,
            in2 => \N__56910\,
            in3 => \N__57054\,
            lcout => \c0.rx.n12862\,
            ltout => \c0.rx.n12862_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_adj_1175_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__59748\,
            in1 => \_gnd_net_\,
            in2 => \N__54058\,
            in3 => \_gnd_net_\,
            lcout => n12973,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_adj_1171_LC_21_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__54054\,
            in1 => \N__54042\,
            in2 => \_gnd_net_\,
            in3 => \N__54030\,
            lcout => \c0.rx.n80\,
            ltout => \c0.rx.n80_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_4_lut_LC_21_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__54283\,
            in1 => \N__54319\,
            in2 => \N__54019\,
            in3 => \N__54300\,
            lcout => \r_SM_Main_2_N_3681_2\,
            ltout => \r_SM_Main_2_N_3681_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_4_lut_LC_21_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001010101"
        )
    port map (
            in0 => \N__56889\,
            in1 => \N__56993\,
            in2 => \N__54346\,
            in3 => \N__56818\,
            lcout => n14283,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i2_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__54320\,
            in1 => \N__54301\,
            in2 => \N__54289\,
            in3 => \N__54262\,
            lcout => \r_SM_Main_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66852\,
            ce => 'H',
            sr => \N__54250\
        );

    \c0.rx.r_Rx_Data_50_LC_22_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54232\,
            lcout => \r_Rx_Data\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i103_LC_22_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__65623\,
            in1 => \N__62432\,
            in2 => \N__54213\,
            in3 => \N__64346\,
            lcout => \c0.data_in_frame_12_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i124_LC_22_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__62431\,
            in1 => \N__68516\,
            in2 => \N__64892\,
            in3 => \N__54189\,
            lcout => \c0.data_in_frame_15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1286_LC_22_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54528\,
            in1 => \N__59245\,
            in2 => \N__56767\,
            in3 => \N__57909\,
            lcout => \c0.n22424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1242_LC_22_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61389\,
            in2 => \_gnd_net_\,
            in3 => \N__54188\,
            lcout => \c0.n22430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i133_LC_22_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66007\,
            in1 => \N__68166\,
            in2 => \N__57324\,
            in3 => \N__63177\,
            lcout => \c0.data_in_frame_16_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1267_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54447\,
            in2 => \_gnd_net_\,
            in3 => \N__54164\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1268_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54541\,
            in1 => \N__57175\,
            in2 => \N__54532\,
            in3 => \N__54529\,
            lcout => \c0.n20240\,
            ltout => \c0.n20240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1309_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58137\,
            in2 => \N__54514\,
            in3 => \N__57313\,
            lcout => \c0.n22385\,
            ltout => \c0.n22385_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1246_LC_22_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55219\,
            in1 => \N__54511\,
            in2 => \N__54481\,
            in3 => \N__61467\,
            lcout => \c0.n29_adj_4234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i118_LC_22_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__67123\,
            in1 => \N__57157\,
            in2 => \_gnd_net_\,
            in3 => \N__54467\,
            lcout => data_in_frame_14_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i80_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62377\,
            in1 => \N__69716\,
            in2 => \N__57370\,
            in3 => \N__68867\,
            lcout => \c0.data_in_frame_9_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i116_LC_22_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__64863\,
            in1 => \N__57158\,
            in2 => \_gnd_net_\,
            in3 => \N__54448\,
            lcout => data_in_frame_14_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i13_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__63175\,
            in1 => \N__69871\,
            in2 => \N__54407\,
            in3 => \N__60898\,
            lcout => data_in_frame_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1548_LC_22_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54432\,
            in2 => \_gnd_net_\,
            in3 => \N__54395\,
            lcout => \c0.n21797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i181_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__63174\,
            in1 => \N__59811\,
            in2 => \_gnd_net_\,
            in3 => \N__59198\,
            lcout => data_in_frame_22_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1269_LC_22_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57345\,
            in1 => \N__59581\,
            in2 => \N__57253\,
            in3 => \N__54778\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4245_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1853_LC_22_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54751\,
            in1 => \N__54718\,
            in2 => \N__54688\,
            in3 => \N__54684\,
            lcout => \c0.n13598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i119_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__65624\,
            in1 => \N__57159\,
            in2 => \_gnd_net_\,
            in3 => \N__55095\,
            lcout => data_in_frame_14_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1291_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60574\,
            in1 => \N__54634\,
            in2 => \_gnd_net_\,
            in3 => \N__54613\,
            lcout => \c0.n22233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i127_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__62538\,
            in1 => \N__68601\,
            in2 => \N__65696\,
            in3 => \N__57870\,
            lcout => \c0.data_in_frame_15_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i92_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67477\,
            in1 => \N__62540\,
            in2 => \N__54592\,
            in3 => \N__64862\,
            lcout => \c0.data_in_frame_11_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1340_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54587\,
            in1 => \N__54571\,
            in2 => \_gnd_net_\,
            in3 => \N__54565\,
            lcout => \c0.n4_adj_4240\,
            ltout => \c0.n4_adj_4240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_4_lut_LC_22_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57817\,
            in2 => \N__54544\,
            in3 => \N__57584\,
            lcout => \c0.n22781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1784_LC_22_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57585\,
            in1 => \N__57217\,
            in2 => \N__61894\,
            in3 => \N__59580\,
            lcout => \c0.n21126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i110_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__67124\,
            in1 => \N__62539\,
            in2 => \N__62149\,
            in3 => \N__61289\,
            lcout => \c0.data_in_frame_13_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i94_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67445\,
            in1 => \N__62500\,
            in2 => \N__57679\,
            in3 => \N__67157\,
            lcout => \c0.data_in_frame_11_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i120_LC_22_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__68865\,
            in1 => \N__57166\,
            in2 => \_gnd_net_\,
            in3 => \N__55057\,
            lcout => data_in_frame_14_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i202_LC_22_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__63826\,
            in1 => \N__69872\,
            in2 => \N__56138\,
            in3 => \N__67776\,
            lcout => \c0.data_in_frame_25_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66721\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1289_LC_22_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__57843\,
            in1 => \N__60937\,
            in2 => \_gnd_net_\,
            in3 => \N__57582\,
            lcout => \c0.n22236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1335_LC_22_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57674\,
            in2 => \_gnd_net_\,
            in3 => \N__54889\,
            lcout => \c0.n6_adj_4273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1264_LC_22_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54853\,
            in1 => \N__60996\,
            in2 => \N__54847\,
            in3 => \N__54828\,
            lcout => \c0.n21982\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1293_LC_22_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57842\,
            in2 => \_gnd_net_\,
            in3 => \N__55137\,
            lcout => \c0.n5813\,
            ltout => \c0.n5813_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1295_LC_22_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__54799\,
            in3 => \N__54906\,
            lcout => \c0.n13728\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1223_LC_22_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55097\,
            in1 => \N__54795\,
            in2 => \N__65404\,
            in3 => \N__54937\,
            lcout => \c0.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1338_LC_22_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57583\,
            in2 => \_gnd_net_\,
            in3 => \N__57540\,
            lcout => OPEN,
            ltout => \c0.n20222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1243_LC_22_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54927\,
            in1 => \N__60450\,
            in2 => \N__55018\,
            in3 => \N__55011\,
            lcout => OPEN,
            ltout => \c0.n28_adj_4232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_3_lut_4_lut_adj_1858_LC_22_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58029\,
            in1 => \N__55096\,
            in2 => \N__54985\,
            in3 => \N__55047\,
            lcout => OPEN,
            ltout => \c0.n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i17_4_lut_LC_22_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57199\,
            in1 => \N__57823\,
            in2 => \N__54982\,
            in3 => \N__54979\,
            lcout => \c0.n21238\,
            ltout => \c0.n21238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_LC_22_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__65759\,
            in1 => \N__54970\,
            in2 => \N__54958\,
            in3 => \N__54955\,
            lcout => \c0.n8_adj_4236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1392_LC_22_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__58172\,
            in1 => \N__65760\,
            in2 => \_gnd_net_\,
            in3 => \N__54936\,
            lcout => \c0.n21831\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i147_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69205\,
            in1 => \N__68111\,
            in2 => \N__57796\,
            in3 => \N__68357\,
            lcout => \c0.data_in_frame_18_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1228_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__54928\,
            in1 => \N__57529\,
            in2 => \N__55065\,
            in3 => \N__61156\,
            lcout => \c0.n22480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1238_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60030\,
            in1 => \N__61322\,
            in2 => \N__58498\,
            in3 => \N__54910\,
            lcout => \c0.n13719\,
            ltout => \c0.n13719_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1249_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61177\,
            in1 => \N__61824\,
            in2 => \N__55144\,
            in3 => \N__55141\,
            lcout => \c0.n14_adj_4238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i149_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__68109\,
            in1 => \N__69206\,
            in2 => \N__58236\,
            in3 => \N__63146\,
            lcout => \c0.data_in_frame_18_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i145_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__69482\,
            in1 => \N__68110\,
            in2 => \N__69233\,
            in3 => \N__57756\,
            lcout => \c0.data_in_frame_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1262_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55119\,
            in2 => \_gnd_net_\,
            in3 => \N__57284\,
            lcout => \c0.n20374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1676_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63918\,
            in1 => \N__63956\,
            in2 => \N__56014\,
            in3 => \N__55509\,
            lcout => \c0.n21067\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1233_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61763\,
            in2 => \_gnd_net_\,
            in3 => \N__61737\,
            lcout => \c0.n22113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3317_2_lut_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55101\,
            in2 => \_gnd_net_\,
            in3 => \N__55066\,
            lcout => \c0.n5996\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i134_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__65937\,
            in1 => \N__68162\,
            in2 => \N__58174\,
            in3 => \N__67170\,
            lcout => \c0.data_in_frame_16_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i195_LC_22_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68417\,
            in1 => \N__65938\,
            in2 => \N__65192\,
            in3 => \N__67756\,
            lcout => \c0.data_in_frame_24_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i131_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__65936\,
            in1 => \N__68161\,
            in2 => \N__58099\,
            in3 => \N__68418\,
            lcout => \c0.data_in_frame_16_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i163_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64517\,
            in1 => \N__68163\,
            in2 => \N__61773\,
            in3 => \N__68419\,
            lcout => \c0.data_in_frame_20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66763\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i140_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69867\,
            in1 => \N__68043\,
            in2 => \N__55429\,
            in3 => \N__64748\,
            lcout => \c0.data_in_frame_17_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64152\,
            in1 => \N__55249\,
            in2 => \N__60037\,
            in3 => \N__55240\,
            lcout => \c0.n20203\,
            ltout => \c0.n20203_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1255_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__55231\,
            in3 => \N__61745\,
            lcout => \c0.n21120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i148_LC_22_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__68042\,
            in1 => \N__69210\,
            in2 => \N__64819\,
            in3 => \N__62900\,
            lcout => \c0.data_in_frame_18_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i125_LC_22_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__63218\,
            in1 => \N__62505\,
            in2 => \N__68659\,
            in3 => \N__58483\,
            lcout => \c0.data_in_frame_15_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i123_LC_22_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__68628\,
            in1 => \N__62504\,
            in2 => \N__55218\,
            in3 => \N__68288\,
            lcout => \c0.data_in_frame_15_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1227_LC_22_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57489\,
            in1 => \N__55183\,
            in2 => \N__55171\,
            in3 => \N__55641\,
            lcout => \c0.n20196\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1719_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__65153\,
            in1 => \N__55447\,
            in2 => \N__59797\,
            in3 => \N__59279\,
            lcout => \c0.n21054\,
            ltout => \c0.n21054_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1722_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62631\,
            in1 => \N__58972\,
            in2 => \N__55441\,
            in3 => \N__55438\,
            lcout => \c0.n14_adj_4484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4028_2_lut_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__59534\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59401\,
            lcout => \c0.n6707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1884_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59400\,
            in1 => \N__59533\,
            in2 => \N__63475\,
            in3 => \N__65230\,
            lcout => \c0.n22323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1229_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55417\,
            in1 => \N__55394\,
            in2 => \_gnd_net_\,
            in3 => \N__55350\,
            lcout => \c0.n12596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1750_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__55351\,
            in1 => \N__55339\,
            in2 => \_gnd_net_\,
            in3 => \N__55302\,
            lcout => \c0.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61848\,
            in1 => \N__55282\,
            in2 => \N__55276\,
            in3 => \N__55497\,
            lcout => \c0.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1661_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55964\,
            in1 => \N__55896\,
            in2 => \N__58846\,
            in3 => \N__58692\,
            lcout => \c0.n20266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1280_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55534\,
            in1 => \N__55255\,
            in2 => \N__62598\,
            in3 => \N__58504\,
            lcout => \c0.n23062\,
            ltout => \c0.n23062_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1282_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__55749\,
            in1 => \_gnd_net_\,
            in2 => \N__55732\,
            in3 => \N__55724\,
            lcout => \c0.n14_adj_4251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_1399_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58429\,
            in1 => \N__55690\,
            in2 => \N__55945\,
            in3 => \N__58741\,
            lcout => \c0.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55564\,
            in1 => \N__61435\,
            in2 => \N__63957\,
            in3 => \N__58459\,
            lcout => \c0.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1222_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55672\,
            in1 => \N__60947\,
            in2 => \N__63421\,
            in3 => \N__55645\,
            lcout => OPEN,
            ltout => \c0.n16_adj_4223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1224_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55625\,
            in1 => \N__58189\,
            in2 => \N__55576\,
            in3 => \N__55573\,
            lcout => \c0.n22211\,
            ltout => \c0.n22211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1225_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55563\,
            in2 => \N__55543\,
            in3 => \N__64069\,
            lcout => \c0.n21140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1207_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56010\,
            in1 => \N__55513\,
            in2 => \_gnd_net_\,
            in3 => \N__55498\,
            lcout => \c0.n23298\,
            ltout => \c0.n23298_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1208_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__55471\,
            in1 => \N__58341\,
            in2 => \N__55462\,
            in3 => \N__58426\,
            lcout => \c0.n21200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i23_4_lut_adj_1729_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__55459\,
            in1 => \N__57952\,
            in2 => \N__55840\,
            in3 => \N__59067\,
            lcout => OPEN,
            ltout => \c0.n52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i26_4_lut_adj_1732_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63547\,
            in1 => \N__58898\,
            in2 => \N__55810\,
            in3 => \N__55774\,
            lcout => \c0.n55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1738_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58644\,
            in2 => \_gnd_net_\,
            in3 => \N__59393\,
            lcout => \c0.n13872\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1653_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58897\,
            in1 => \N__58645\,
            in2 => \N__59408\,
            in3 => \N__59019\,
            lcout => \c0.n12420\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i199_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__67758\,
            in1 => \N__65575\,
            in2 => \N__59407\,
            in3 => \N__65939\,
            lcout => \c0.data_in_frame_24_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1199_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61642\,
            in2 => \_gnd_net_\,
            in3 => \N__55783\,
            lcout => \c0.n22468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i15_3_lut_4_lut_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62791\,
            in1 => \N__58713\,
            in2 => \N__58845\,
            in3 => \N__59289\,
            lcout => \c0.n44_adj_4490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i19_4_lut_adj_1725_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__69280\,
            in1 => \N__58896\,
            in2 => \N__66096\,
            in3 => \N__59079\,
            lcout => OPEN,
            ltout => \c0.n48_adj_4485_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i24_4_lut_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58561\,
            in1 => \N__56020\,
            in2 => \N__55768\,
            in3 => \N__66908\,
            lcout => \c0.n53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1371_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55938\,
            in1 => \N__66128\,
            in2 => \N__65275\,
            in3 => \N__55765\,
            lcout => \c0.n22719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1654_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56142\,
            in1 => \N__63490\,
            in2 => \_gnd_net_\,
            in3 => \N__65247\,
            lcout => \c0.n20370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i28_4_lut_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__56107\,
            in1 => \N__56092\,
            in2 => \N__58570\,
            in3 => \N__56086\,
            lcout => \c0.n23416\,
            ltout => \c0.n23416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1380_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59080\,
            in1 => \N__63439\,
            in2 => \N__56068\,
            in3 => \N__59071\,
            lcout => \c0.n12_adj_4296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_adj_1829_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55966\,
            in1 => \N__56053\,
            in2 => \N__56283\,
            in3 => \N__55846\,
            lcout => \c0.n36_adj_4489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1659_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__55999\,
            in1 => \N__55890\,
            in2 => \N__58836\,
            in3 => \N__63900\,
            lcout => \c0.n22388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1782_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63901\,
            in1 => \N__55965\,
            in2 => \N__55897\,
            in3 => \N__63958\,
            lcout => \c0.n21037\,
            ltout => \c0.n21037_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1391_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58327\,
            in1 => \N__55924\,
            in2 => \N__55900\,
            in3 => \N__58427\,
            lcout => \c0.n13993\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1236_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__55894\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58822\,
            lcout => \c0.n13282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_adj_1370_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56322\,
            in1 => \N__56304\,
            in2 => \_gnd_net_\,
            in3 => \N__56293\,
            lcout => OPEN,
            ltout => \c0.n8_adj_4291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i20116_4_lut_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__56278\,
            in1 => \N__56248\,
            in2 => \N__56242\,
            in3 => \N__56239\,
            lcout => \c0.n23811\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i7_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__68784\,
            in1 => \N__59958\,
            in2 => \N__56220\,
            in3 => \N__59699\,
            lcout => rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i12_3_lut_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__56810\,
            in1 => \N__59698\,
            in2 => \_gnd_net_\,
            in3 => \N__56186\,
            lcout => \c0.rx.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_4_lut_4_lut_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__56992\,
            in1 => \N__56809\,
            in2 => \N__56928\,
            in3 => \N__57058\,
            lcout => n14436,
            ltout => \n14436_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i11380_3_lut_4_lut_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__59747\,
            in1 => \N__56914\,
            in2 => \N__56164\,
            in3 => \N__59957\,
            lcout => n14917,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i2_3_lut_adj_1174_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__57091\,
            in1 => \N__59863\,
            in2 => \_gnd_net_\,
            in3 => \N__56161\,
            lcout => n12970,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i2_LC_22_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__59898\,
            in1 => \N__57115\,
            in2 => \N__57101\,
            in3 => \N__59911\,
            lcout => \r_Bit_Index_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i0_LC_22_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000010101010"
        )
    port map (
            in0 => \N__59752\,
            in1 => \_gnd_net_\,
            in2 => \N__56946\,
            in3 => \N__59897\,
            lcout => \r_Bit_Index_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i15930_2_lut_LC_22_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__59751\,
            in1 => \_gnd_net_\,
            in2 => \N__59868\,
            in3 => \_gnd_net_\,
            lcout => n19619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i1_2_lut_LC_22_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59859\,
            in2 => \_gnd_net_\,
            in3 => \N__57090\,
            lcout => n91,
            ltout => \n91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.i28_3_lut_4_lut_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011001100"
        )
    port map (
            in0 => \N__59750\,
            in1 => \N__56822\,
            in2 => \N__57064\,
            in3 => \N__57060\,
            lcout => OPEN,
            ltout => \c0.rx.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_SM_Main_i0_LC_22_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001010001"
        )
    port map (
            in0 => \N__57002\,
            in1 => \N__56939\,
            in2 => \N__56845\,
            in3 => \N__56842\,
            lcout => \r_SM_Main_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_69_i9_2_lut_3_lut_LC_23_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__56718\,
            in1 => \N__56598\,
            in2 => \_gnd_net_\,
            in3 => \N__56457\,
            lcout => \c0.n9_adj_4217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1260_LC_23_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__57126\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60234\,
            lcout => \c0.n22328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1664_LC_23_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__56692\,
            in1 => \N__56597\,
            in2 => \N__56458\,
            in3 => \N__62351\,
            lcout => n21755,
            ltout => \n21755_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i114_LC_23_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63831\,
            in2 => \N__56770\,
            in3 => \N__56763\,
            lcout => data_in_frame_14_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.equal_68_i9_2_lut_3_lut_LC_23_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__56691\,
            in1 => \N__56596\,
            in2 => \_gnd_net_\,
            in3 => \N__56439\,
            lcout => \c0.n9_adj_4237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1265_LC_23_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57382\,
            in2 => \_gnd_net_\,
            in3 => \N__57365\,
            lcout => \c0.n22471\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1382_LC_23_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__57314\,
            in1 => \N__58205\,
            in2 => \_gnd_net_\,
            in3 => \N__57283\,
            lcout => \c0.n21069\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1266_LC_23_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60255\,
            in1 => \N__57940\,
            in2 => \N__57187\,
            in3 => \N__57910\,
            lcout => \c0.n22446\,
            ltout => \c0.n22446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1244_LC_23_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58497\,
            in1 => \N__57234\,
            in2 => \N__57220\,
            in3 => \N__57216\,
            lcout => \c0.n30_adj_4233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i115_LC_23_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__57186\,
            in1 => \N__57155\,
            in2 => \_gnd_net_\,
            in3 => \N__68443\,
            lcout => data_in_frame_14_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1304_LC_23_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60233\,
            in2 => \_gnd_net_\,
            in3 => \N__60254\,
            lcout => \c0.n22340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i113_LC_23_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__57924\,
            in1 => \N__57154\,
            in2 => \_gnd_net_\,
            in3 => \N__69493\,
            lcout => data_in_frame_14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i117_LC_23_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__57156\,
            in1 => \N__63176\,
            in2 => \_gnd_net_\,
            in3 => \N__57127\,
            lcout => data_in_frame_14_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i192_LC_23_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__68155\,
            in1 => \N__68591\,
            in2 => \N__65297\,
            in3 => \N__68979\,
            lcout => \c0.data_in_frame_23_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i146_LC_23_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__69203\,
            in1 => \N__68156\,
            in2 => \N__57469\,
            in3 => \N__63859\,
            lcout => \c0.data_in_frame_18_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66707\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_2_lut_3_lut_LC_23_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__57447\,
            in1 => \N__57869\,
            in2 => \_gnd_net_\,
            in3 => \N__61284\,
            lcout => \c0.n10_adj_4239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1327_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60907\,
            in1 => \N__57498\,
            in2 => \N__61290\,
            in3 => \N__57523\,
            lcout => \c0.n22464\,
            ltout => \c0.n22464_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_4_lut_adj_1785_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60383\,
            in1 => \N__60172\,
            in2 => \N__57514\,
            in3 => \N__57511\,
            lcout => \c0.n8_adj_4275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1788_LC_23_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58067\,
            in1 => \N__60232\,
            in2 => \_gnd_net_\,
            in3 => \N__60253\,
            lcout => \c0.n10_adj_4267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1250_LC_23_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57499\,
            in1 => \N__61329\,
            in2 => \N__58036\,
            in3 => \N__58068\,
            lcout => \c0.n14053\,
            ltout => \c0.n14053_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1347_LC_23_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__57468\,
            in1 => \N__61242\,
            in2 => \N__57451\,
            in3 => \N__60531\,
            lcout => OPEN,
            ltout => \c0.n23586_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1297_LC_23_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62677\,
            in1 => \N__57448\,
            in2 => \N__57406\,
            in3 => \N__61285\,
            lcout => \c0.n23426\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1288_LC_23_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__61003\,
            in1 => \N__60002\,
            in2 => \_gnd_net_\,
            in3 => \N__57403\,
            lcout => \c0.n13210\,
            ltout => \c0.n13210_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1342_LC_23_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__57736\,
            in3 => \N__57733\,
            lcout => OPEN,
            ltout => \c0.n7_adj_4277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_adj_1343_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60121\,
            in1 => \N__57691\,
            in2 => \N__57682\,
            in3 => \N__60406\,
            lcout => \c0.n21867\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i93_LC_23_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__67476\,
            in1 => \N__63124\,
            in2 => \N__61045\,
            in3 => \N__62531\,
            lcout => \c0.data_in_frame_11_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1789_LC_23_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60139\,
            in1 => \N__57605\,
            in2 => \_gnd_net_\,
            in3 => \N__60511\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1322_LC_23_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61040\,
            in1 => \N__57675\,
            in2 => \N__57658\,
            in3 => \N__57632\,
            lcout => \c0.n16_adj_4265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i95_LC_23_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__62529\,
            in1 => \N__65569\,
            in2 => \N__57639\,
            in3 => \N__67451\,
            lcout => \c0.data_in_frame_11_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i91_LC_23_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__67475\,
            in1 => \N__68437\,
            in2 => \N__57614\,
            in3 => \N__62530\,
            lcout => \c0.data_in_frame_11_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66735\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1344_LC_23_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61517\,
            in2 => \_gnd_net_\,
            in3 => \N__58098\,
            lcout => \c0.n21845\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1565_LC_23_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57850\,
            in1 => \N__57592\,
            in2 => \N__57553\,
            in3 => \N__57541\,
            lcout => \c0.n6_adj_4225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_LC_23_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__57936\,
            in1 => \N__57925\,
            in2 => \_gnd_net_\,
            in3 => \N__57908\,
            lcout => \c0.n22352\,
            ltout => \c0.n22352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1253_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57874\,
            in1 => \N__57849\,
            in2 => \N__57829\,
            in3 => \N__61235\,
            lcout => \c0.n22000\,
            ltout => \c0.n22000_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i13_4_lut_adj_1245_LC_23_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__57809\,
            in1 => \N__61172\,
            in2 => \N__57826\,
            in3 => \N__60546\,
            lcout => \c0.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i128_LC_23_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__62541\,
            in1 => \N__57810\,
            in2 => \N__68680\,
            in3 => \N__68908\,
            lcout => \c0.data_in_frame_15_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i100_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62557\,
            in1 => \N__64481\,
            in2 => \N__61500\,
            in3 => \N__64874\,
            lcout => \c0.data_in_frame_12_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_4_lut_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61254\,
            in1 => \N__61518\,
            in2 => \N__57795\,
            in3 => \N__61884\,
            lcout => OPEN,
            ltout => \c0.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1254_LC_23_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64173\,
            in1 => \N__57778\,
            in2 => \N__57769\,
            in3 => \N__58062\,
            lcout => \c0.n20246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1251_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58061\,
            in1 => \N__57766\,
            in2 => \N__57757\,
            in3 => \N__57742\,
            lcout => \c0.n13544\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1237_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58243\,
            in1 => \N__61149\,
            in2 => \N__58237\,
            in3 => \N__58212\,
            lcout => \c0.n10_adj_4230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_3_lut_4_lut_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58018\,
            in1 => \N__58185\,
            in2 => \N__58173\,
            in3 => \N__58063\,
            lcout => \c0.n18_adj_4246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_LC_23_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__58141\,
            in1 => \N__58094\,
            in2 => \_gnd_net_\,
            in3 => \N__58075\,
            lcout => \c0.n22849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i201_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__69565\,
            in1 => \N__58637\,
            in2 => \N__69878\,
            in3 => \N__67757\,
            lcout => \c0.data_in_frame_25_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i109_LC_23_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__63139\,
            in1 => \N__62058\,
            in2 => \N__58069\,
            in3 => \N__62507\,
            lcout => \c0.data_in_frame_13_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i126_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__68678\,
            in1 => \N__62506\,
            in2 => \N__58028\,
            in3 => \N__67070\,
            lcout => \c0.data_in_frame_15_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1190_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62787\,
            in1 => \N__65146\,
            in2 => \N__57997\,
            in3 => \N__57973\,
            lcout => \c0.n22402\,
            ltout => \c0.n22402_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_3_lut_4_lut_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59488\,
            in1 => \N__65061\,
            in2 => \N__57955\,
            in3 => \N__65179\,
            lcout => \c0.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i213_LC_23_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__63225\,
            in1 => \N__69204\,
            in2 => \N__59499\,
            in3 => \N__67759\,
            lcout => \c0.data_in_frame_26_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_adj_1372_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__59489\,
            in1 => \N__64947\,
            in2 => \_gnd_net_\,
            in3 => \N__58390\,
            lcout => OPEN,
            ltout => \c0.n6_adj_4292_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1379_LC_23_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65062\,
            in1 => \N__58996\,
            in2 => \N__58384\,
            in3 => \N__58381\,
            lcout => \c0.n23073\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1277_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58342\,
            in1 => \N__58300\,
            in2 => \N__61209\,
            in3 => \N__62850\,
            lcout => \c0.n24_adj_4248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1348_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62765\,
            in2 => \_gnd_net_\,
            in3 => \N__58256\,
            lcout => \c0.n21905\,
            ltout => \c0.n21905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1349_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61667\,
            in1 => \N__62893\,
            in2 => \N__58294\,
            in3 => \N__64111\,
            lcout => \c0.n20288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1270_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65719\,
            in1 => \N__66049\,
            in2 => \_gnd_net_\,
            in3 => \N__58291\,
            lcout => \c0.n22399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1739_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__58257\,
            in1 => \N__58279\,
            in2 => \N__59832\,
            in3 => \N__62702\,
            lcout => \c0.n22020\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i164_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64535\,
            in1 => \N__68086\,
            in2 => \N__58261\,
            in3 => \N__64853\,
            lcout => \c0.data_in_frame_20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i196_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__64852\,
            in1 => \N__66001\,
            in2 => \N__59006\,
            in3 => \N__67676\,
            lcout => \c0.data_in_frame_24_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1856_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__61741\,
            in1 => \N__61666\,
            in2 => \N__62706\,
            in3 => \N__58541\,
            lcout => \c0.n22458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i165_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__62766\,
            in1 => \N__63178\,
            in2 => \N__68147\,
            in3 => \N__64536\,
            lcout => \c0.data_in_frame_20_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_2_lut_4_lut_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59335\,
            in1 => \N__58446\,
            in2 => \N__63310\,
            in3 => \N__58458\,
            lcout => OPEN,
            ltout => \c0.n18_adj_4249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1279_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__65364\,
            in1 => \N__58528\,
            in2 => \N__58516\,
            in3 => \N__58513\,
            lcout => \c0.n26_adj_4250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_adj_1272_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64054\,
            in1 => \N__58490\,
            in2 => \N__63416\,
            in3 => \N__61786\,
            lcout => \c0.n23072\,
            ltout => \c0.n23072_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1274_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__58447\,
            in1 => \_gnd_net_\,
            in2 => \N__58432\,
            in3 => \N__63308\,
            lcout => \c0.n22364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1256_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62707\,
            in2 => \_gnd_net_\,
            in3 => \N__61668\,
            lcout => \c0.n21124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1284_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58428\,
            in1 => \N__63316\,
            in2 => \N__65400\,
            in3 => \N__58396\,
            lcout => \c0.n21039\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i161_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__59336\,
            in1 => \N__69560\,
            in2 => \N__68164\,
            in3 => \N__64560\,
            lcout => \c0.data_in_frame_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1356_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__58837\,
            in1 => \N__58774\,
            in2 => \_gnd_net_\,
            in3 => \N__58726\,
            lcout => \c0.n14_adj_4283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i9_4_lut_adj_1352_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60490\,
            in1 => \N__61695\,
            in2 => \N__60277\,
            in3 => \N__58740\,
            lcout => OPEN,
            ltout => \c0.n24_adj_4282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i14_4_lut_adj_1354_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59770\,
            in1 => \N__65206\,
            in2 => \N__58729\,
            in3 => \N__63238\,
            lcout => \c0.n22711\,
            ltout => \c0.n22711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1209_LC_23_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63560\,
            in2 => \N__58720\,
            in3 => \N__58712\,
            lcout => \c0.n21087\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1357_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63432\,
            in1 => \N__58696\,
            in2 => \N__58675\,
            in3 => \N__58651\,
            lcout => OPEN,
            ltout => \c0.n15_adj_4284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_adj_1359_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62599\,
            in1 => \N__63877\,
            in2 => \N__58660\,
            in3 => \N__58657\,
            lcout => \c0.n22373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1212_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__69595\,
            in2 => \_gnd_net_\,
            in3 => \N__59031\,
            lcout => \c0.n22437\,
            ltout => \c0.n22437_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i21_4_lut_adj_1730_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58643\,
            in1 => \N__58618\,
            in2 => \N__58573\,
            in3 => \N__59044\,
            lcout => \c0.n50_adj_4487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1904_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63501\,
            in1 => \N__58560\,
            in2 => \N__63546\,
            in3 => \N__59065\,
            lcout => \c0.n20537\,
            ltout => \c0.n20537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1723_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59104\,
            in1 => \N__59256\,
            in2 => \N__59095\,
            in3 => \N__59092\,
            lcout => \c0.n21890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1563_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58953\,
            in1 => \N__65193\,
            in2 => \N__65053\,
            in3 => \N__59008\,
            lcout => \c0.n13320\,
            ltout => \c0.n13320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_LC_23_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__59066\,
            in1 => \N__68712\,
            in2 => \N__59047\,
            in3 => \N__59043\,
            lcout => OPEN,
            ltout => \c0.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_4_lut_adj_1897_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__64258\,
            in1 => \N__64224\,
            in2 => \N__59035\,
            in3 => \N__59032\,
            lcout => \c0.n22314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1210_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59007\,
            in2 => \_gnd_net_\,
            in3 => \N__58952\,
            lcout => \c0.n22142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1206_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__58960\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59257\,
            lcout => \c0.n22337\,
            ltout => \c0.n22337_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1743_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__58852\,
            in1 => \N__58918\,
            in2 => \N__58906\,
            in3 => \N__58903\,
            lcout => \c0.n21095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_4_lut_adj_1651_LC_23_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59446\,
            in1 => \N__66066\,
            in2 => \N__68705\,
            in3 => \N__59409\,
            lcout => \c0.n6_adj_4418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1361_LC_23_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59500\,
            in1 => \N__64911\,
            in2 => \N__64275\,
            in3 => \N__59470\,
            lcout => OPEN,
            ltout => \c0.n10_adj_4285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_3_lut_adj_1373_LC_23_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62635\,
            in2 => \N__59464\,
            in3 => \N__65016\,
            lcout => \c0.n22995\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1741_LC_23_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59445\,
            in2 => \_gnd_net_\,
            in3 => \N__68695\,
            lcout => \c0.n22054\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1740_LC_23_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66067\,
            in2 => \_gnd_net_\,
            in3 => \N__59410\,
            lcout => \c0.n22434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1203_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__59352\,
            in1 => \N__61641\,
            in2 => \N__59317\,
            in3 => \N__59290\,
            lcout => \c0.n20596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i96_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__68785\,
            in1 => \N__62508\,
            in2 => \N__67480\,
            in3 => \N__59226\,
            lcout => \c0.data_in_frame_11_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i180_LC_23_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__64885\,
            in1 => \N__61694\,
            in2 => \_gnd_net_\,
            in3 => \N__59212\,
            lcout => data_in_frame_22_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i174_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__65357\,
            in1 => \N__66974\,
            in2 => \N__62121\,
            in3 => \N__68160\,
            lcout => \c0.data_in_frame_21_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63573\,
            in1 => \N__65356\,
            in2 => \N__59125\,
            in3 => \N__59976\,
            lcout => \c0.n22215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i156_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67471\,
            in1 => \N__68159\,
            in2 => \N__63917\,
            in3 => \N__64886\,
            lcout => \c0.data_in_frame_19_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i6_LC_23_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__65501\,
            in1 => \N__59965\,
            in2 => \N__59709\,
            in3 => \N__59939\,
            lcout => rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i4_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__62975\,
            in1 => \N__59756\,
            in2 => \N__59715\,
            in3 => \N__59592\,
            lcout => rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Bit_Index_i1_LC_23_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__59910\,
            in1 => \N__59864\,
            in2 => \N__59758\,
            in3 => \N__59899\,
            lcout => \r_Bit_Index_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1353_LC_23_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__67811\,
            in1 => \N__59833\,
            in2 => \N__62752\,
            in3 => \N__59787\,
            lcout => \c0.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.rx.r_Rx_Byte_i5_LC_23_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__59757\,
            in1 => \N__59708\,
            in2 => \N__59593\,
            in3 => \N__66975\,
            lcout => rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i97_LC_24_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64345\,
            in1 => \N__62378\,
            in2 => \N__59578\,
            in3 => \N__69502\,
            lcout => \c0.data_in_frame_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66708\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i200_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__68980\,
            in1 => \N__66030\,
            in2 => \N__59522\,
            in3 => \N__67775\,
            lcout => \c0.data_in_frame_24_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66722\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i98_LC_24_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64356\,
            in1 => \N__62525\,
            in2 => \N__60259\,
            in3 => \N__63861\,
            lcout => \c0.data_in_frame_12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66722\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i99_LC_24_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__62522\,
            in1 => \N__64357\,
            in2 => \N__68442\,
            in3 => \N__60235\,
            lcout => \c0.data_in_frame_12_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66722\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i107_LC_24_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61970\,
            in1 => \N__62524\,
            in2 => \N__60211\,
            in3 => \N__68433\,
            lcout => \c0.data_in_frame_13_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66722\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1786_LC_24_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__60207\,
            in1 => \N__61138\,
            in2 => \_gnd_net_\,
            in3 => \N__61107\,
            lcout => \c0.n22274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i106_LC_24_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__61969\,
            in1 => \N__62523\,
            in2 => \N__60195\,
            in3 => \N__63860\,
            lcout => \c0.data_in_frame_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66722\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i89_LC_24_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__67408\,
            in1 => \N__69492\,
            in2 => \N__60150\,
            in3 => \N__62527\,
            lcout => \c0.data_in_frame_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1305_LC_24_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60143\,
            in2 => \_gnd_net_\,
            in3 => \N__60512\,
            lcout => OPEN,
            ltout => \c0.n13999_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1248_LC_24_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60117\,
            in1 => \N__60102\,
            in2 => \N__60061\,
            in3 => \N__60058\,
            lcout => \c0.n13233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i75_LC_24_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__62526\,
            in1 => \N__69880\,
            in2 => \N__68441\,
            in3 => \N__60003\,
            lcout => \c0.data_in_frame_9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1346_LC_24_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60553\,
            in1 => \N__61542\,
            in2 => \N__61261\,
            in3 => \N__60535\,
            lcout => \c0.n21114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3286_2_lut_LC_24_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62671\,
            in2 => \_gnd_net_\,
            in3 => \N__61886\,
            lcout => \c0.n5965\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i90_LC_24_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__63793\,
            in1 => \N__67457\,
            in2 => \N__60519\,
            in3 => \N__62528\,
            lcout => \c0.data_in_frame_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i188_LC_24_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__68157\,
            in1 => \N__68552\,
            in2 => \N__60482\,
            in3 => \N__64873\,
            lcout => \c0.data_in_frame_23_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66750\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i186_LC_24_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__60333\,
            in1 => \N__63830\,
            in2 => \N__68590\,
            in3 => \N__68158\,
            lcout => \c0.data_in_frame_23_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66750\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_4_lut_adj_1341_LC_24_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__60451\,
            in1 => \N__60436\,
            in2 => \N__60421\,
            in3 => \N__60412\,
            lcout => \c0.n8_adj_4276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i105_LC_24_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62544\,
            in1 => \N__62120\,
            in2 => \N__60398\,
            in3 => \N__69564\,
            lcout => \c0.data_in_frame_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66750\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i104_LC_24_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__68866\,
            in1 => \N__62545\,
            in2 => \N__64458\,
            in3 => \N__60356\,
            lcout => \c0.data_in_frame_12_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66750\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1281_LC_24_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60329\,
            in2 => \_gnd_net_\,
            in3 => \N__60311\,
            lcout => \c0.n21995\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i59_LC_24_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__60863\,
            in1 => \N__68553\,
            in2 => \N__60997\,
            in3 => \N__68434\,
            lcout => \c0.data_in_frame_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66750\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i176_LC_24_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62086\,
            in1 => \N__68148\,
            in2 => \N__61202\,
            in3 => \N__68909\,
            lcout => \c0.data_in_frame_21_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1859_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__61887\,
            in1 => \N__62672\,
            in2 => \_gnd_net_\,
            in3 => \N__61176\,
            lcout => \c0.n22091\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1578_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61131\,
            in2 => \_gnd_net_\,
            in3 => \N__61111\,
            lcout => \c0.n13421\,
            ltout => \c0.n13421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i4_4_lut_adj_1287_LC_24_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61044\,
            in1 => \N__60972\,
            in2 => \N__61027\,
            in3 => \N__61023\,
            lcout => \c0.n10_adj_4252\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1303_LC_24_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__60989\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60566\,
            lcout => \c0.n22343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_4_lut_adj_1325_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__61312\,
            in1 => \N__60958\,
            in2 => \N__60949\,
            in3 => \N__61448\,
            lcout => \c0.n16_adj_4268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i57_LC_24_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__68545\,
            in1 => \N__60567\,
            in2 => \N__60893\,
            in3 => \N__69450\,
            lcout => \c0.data_in_frame_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i166_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__68143\,
            in1 => \N__64534\,
            in2 => \N__63309\,
            in3 => \N__67104\,
            lcout => \c0.data_in_frame_20_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i130_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__65992\,
            in1 => \N__68144\,
            in2 => \N__61525\,
            in3 => \N__63851\,
            lcout => \c0.data_in_frame_16_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i160_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__68142\,
            in1 => \N__67453\,
            in2 => \N__63355\,
            in3 => \N__68971\,
            lcout => \c0.data_in_frame_19_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1299_LC_24_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61343\,
            in2 => \_gnd_net_\,
            in3 => \N__61481\,
            lcout => \c0.n21975\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i5_2_lut_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61434\,
            in2 => \_gnd_net_\,
            in3 => \N__61390\,
            lcout => \c0.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i101_LC_24_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__64533\,
            in1 => \N__62556\,
            in2 => \N__61359\,
            in3 => \N__63161\,
            lcout => \c0.data_in_frame_12_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i108_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__62555\,
            in1 => \N__62087\,
            in2 => \N__61330\,
            in3 => \N__64875\,
            lcout => \c0.data_in_frame_13_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1345_LC_24_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62661\,
            in2 => \_gnd_net_\,
            in3 => \N__61294\,
            lcout => \c0.n14081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i129_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__65940\,
            in1 => \N__68145\,
            in2 => \N__61243\,
            in3 => \N__69566\,
            lcout => \c0.data_in_frame_16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1197_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63295\,
            in1 => \N__62770\,
            in2 => \N__62751\,
            in3 => \N__62698\,
            lcout => \c0.n22105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i111_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__65570\,
            in1 => \N__62503\,
            in2 => \N__62676\,
            in3 => \N__62181\,
            lcout => \c0.data_in_frame_13_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i214_LC_24_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69151\,
            in1 => \N__67103\,
            in2 => \N__62630\,
            in3 => \N__67744\,
            lcout => \c0.data_in_frame_26_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i175_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__65571\,
            in1 => \N__68146\,
            in2 => \N__62591\,
            in3 => \N__62182\,
            lcout => \c0.data_in_frame_21_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i112_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__62502\,
            in1 => \N__68970\,
            in2 => \N__62203\,
            in3 => \N__61885\,
            lcout => \c0.data_in_frame_13_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i7_3_lut_4_lut_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__61852\,
            in1 => \N__61828\,
            in2 => \N__62901\,
            in3 => \N__64207\,
            lcout => \c0.n20_adj_4247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_3_lut_4_lut_adj_1896_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__61774\,
            in1 => \N__61746\,
            in2 => \N__61708\,
            in3 => \N__61672\,
            lcout => \c0.n22007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1257_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63351\,
            in2 => \_gnd_net_\,
            in3 => \N__61618\,
            lcout => \c0.n13768\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1276_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__61578\,
            in1 => \N__61561\,
            in2 => \_gnd_net_\,
            in3 => \N__61546\,
            lcout => \c0.n14143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i154_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67469\,
            in1 => \N__68087\,
            in2 => \N__63417\,
            in3 => \N__63813\,
            lcout => \c0.data_in_frame_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i198_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67673\,
            in1 => \N__65949\,
            in2 => \N__63539\,
            in3 => \N__67063\,
            lcout => \c0.data_in_frame_24_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1283_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__63387\,
            in1 => \N__63364\,
            in2 => \N__63358\,
            in3 => \N__64123\,
            lcout => \c0.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1351_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__63304\,
            in1 => \N__62869\,
            in2 => \N__62827\,
            in3 => \N__63267\,
            lcout => \c0.n26_adj_4281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i229_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__64498\,
            in1 => \N__63106\,
            in2 => \N__64932\,
            in3 => \N__67674\,
            lcout => \c0.data_in_frame_28_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_adj_1496_LC_24_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__62902\,
            in1 => \N__64110\,
            in2 => \_gnd_net_\,
            in3 => \N__64219\,
            lcout => \c0.n22095\,
            ltout => \c0.n22095_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i12_4_lut_LC_24_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__62863\,
            in1 => \N__66048\,
            in2 => \N__62857\,
            in3 => \N__62854\,
            lcout => \c0.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1883_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62826\,
            in2 => \_gnd_net_\,
            in3 => \N__63876\,
            lcout => \c0.n22267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_adj_1198_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64244\,
            in2 => \_gnd_net_\,
            in3 => \N__64220\,
            lcout => \c0.n20406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_4_lut_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64177\,
            in1 => \N__64156\,
            in2 => \N__64135\,
            in3 => \N__64122\,
            lcout => OPEN,
            ltout => \c0.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i11_4_lut_adj_1271_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__64109\,
            in1 => \N__64084\,
            in2 => \N__64072\,
            in3 => \N__64065\,
            lcout => \c0.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i10_4_lut_adj_1218_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64048\,
            in1 => \N__64036\,
            in2 => \N__63994\,
            in3 => \N__63979\,
            lcout => \c0.n23287\,
            ltout => \c0.n23287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_4_lut_adj_1355_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__65304\,
            in1 => \N__65365\,
            in2 => \N__63922\,
            in3 => \N__63919\,
            lcout => \c0.n21921\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i194_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67791\,
            in1 => \N__66003\,
            in2 => \N__65060\,
            in3 => \N__63852\,
            lcout => \c0.data_in_frame_24_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i193_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__66002\,
            in1 => \N__69451\,
            in2 => \N__63574\,
            in3 => \N__67792\,
            lcout => \c0.data_in_frame_24_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_2_lut_3_lut_4_lut_adj_1564_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__65246\,
            in1 => \N__63538\,
            in2 => \N__63505\,
            in3 => \N__63485\,
            lcout => \c0.n22255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i8_3_lut_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65305\,
            in1 => \N__65265\,
            in2 => \_gnd_net_\,
            in3 => \N__65245\,
            lcout => \c0.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i1_4_lut_adj_1205_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__65200\,
            in1 => \N__65154\,
            in2 => \N__65113\,
            in3 => \N__65080\,
            lcout => \c0.n22455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_3_lut_adj_1365_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__65059\,
            in1 => \N__65020\,
            in2 => \_gnd_net_\,
            in3 => \N__64989\,
            lcout => OPEN,
            ltout => \c0.n8_adj_4288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i6_4_lut_adj_1368_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010110"
        )
    port map (
            in0 => \N__64599\,
            in1 => \N__64963\,
            in2 => \N__64975\,
            in3 => \N__64900\,
            lcout => \c0.n24_adj_4289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3_4_lut_adj_1366_LC_24_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__64962\,
            in1 => \N__64951\,
            in2 => \N__64933\,
            in3 => \N__64912\,
            lcout => \c0.n22997\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i228_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__64511\,
            in1 => \N__64864\,
            in2 => \N__64603\,
            in3 => \N__67794\,
            lcout => \c0.data_in_frame_28_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i232_LC_24_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67793\,
            in1 => \N__64513\,
            in2 => \N__64587\,
            in3 => \N__68883\,
            lcout => \c0.data_in_frame_28_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i231_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__64512\,
            in1 => \N__65574\,
            in2 => \N__64276\,
            in3 => \N__67795\,
            lcout => \c0.data_in_frame_28_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i224_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__66124\,
            in1 => \N__68882\,
            in2 => \N__67479\,
            in3 => \N__67750\,
            lcout => \c0.data_in_frame_27_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i223_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67748\,
            in1 => \N__67462\,
            in2 => \N__66095\,
            in3 => \N__65503\,
            lcout => \c0.data_in_frame_27_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i217_LC_24_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__69561\,
            in1 => \N__66065\,
            in2 => \N__67478\,
            in3 => \N__67749\,
            lcout => \c0.data_in_frame_27_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i3589_2_lut_LC_24_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65417\,
            in2 => \_gnd_net_\,
            in3 => \N__65378\,
            lcout => \c0.n6268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i136_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__66031\,
            in1 => \N__68137\,
            in2 => \N__65750\,
            in3 => \N__68881\,
            lcout => \c0.data_in_frame_16_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i153_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__68136\,
            in1 => \N__67461\,
            in2 => \N__65718\,
            in3 => \N__69562\,
            lcout => \c0.data_in_frame_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i151_LC_24_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__65502\,
            in1 => \N__69199\,
            in2 => \N__65424\,
            in3 => \N__68138\,
            lcout => \c0.data_in_frame_18_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i152_LC_24_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__68135\,
            in1 => \N__65379\,
            in2 => \N__69232\,
            in3 => \N__68876\,
            lcout => \c0.data_in_frame_18_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.i2_3_lut_adj_1360_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__69584\,
            in1 => \N__69269\,
            in2 => \_gnd_net_\,
            in3 => \N__65355\,
            lcout => \c0.n22123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i208_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69879\,
            in1 => \N__68938\,
            in2 => \N__69594\,
            in3 => \N__67777\,
            lcout => \c0.data_in_frame_25_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i209_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67763\,
            in1 => \N__69198\,
            in2 => \N__69279\,
            in3 => \N__69452\,
            lcout => \c0.data_in_frame_26_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i216_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__69197\,
            in1 => \N__68939\,
            in2 => \N__68713\,
            in3 => \N__67778\,
            lcout => \c0.data_in_frame_26_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i187_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__68589\,
            in1 => \N__68435\,
            in2 => \N__67819\,
            in3 => \N__68165\,
            lcout => \c0.data_in_frame_23_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \c0.data_in_frame_0__i222_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__67764\,
            in1 => \N__67470\,
            in2 => \N__66912\,
            in3 => \N__67005\,
            lcout => \c0.data_in_frame_27_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__66863\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
