// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Aug 26 01:16:35 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    inout PIN_1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    inout PIN_2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    input PIN_4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    input PIN_5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    input PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    input PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    input PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    input PIN_12 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    input PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    input PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    input PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    input PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    input PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    input PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire GND_net, VCC_net, LED_c, tx_o, tx2_o, tx_enable, tx2_enable, 
        rx_i;
    wire [25:0]blink_counter;   // verilog/TinyFPGA_B.v(64[14:27])
    
    wire n4720;
    wire [15:0]data;   // coms.v(14[14:18])
    wire [7:0]\data_out[19] ;   // coms.v(15[12:20])
    wire [7:0]\data_out[18] ;   // coms.v(15[12:20])
    
    wire n4719, n2528;
    wire [7:0]\data_out[11] ;   // coms.v(15[12:20])
    wire [7:0]\data_out[10] ;   // coms.v(15[12:20])
    
    wire n2527, n4718, n4734, n2526, n2486, n2525, n2524, n4717, 
        n2388, n2522, n2510, n2521, n2520, rx_data_ready;
    wire [7:0]rx_data;   // coms.v(167[14:21])
    wire [7:0]\data_in[19] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[18] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[17] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[16] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[15] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[14] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[13] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[12] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[11] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[10] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[9] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[8] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[7] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[6] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[5] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[4] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[3] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[2] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[1] ;   // coms.v(171[13:20])
    wire [7:0]\data_in[0] ;   // coms.v(171[13:20])
    
    wire tx2_active, n1519, n4333, n4334, n4733, n4732, n135, 
        n5818, n2519, n2512, n2508, n5424, n2511, n2484, n4731, 
        n4, n5433, n4_adj_1973, n2492, n4716, n2505, n2504, n3636, 
        n5421, n4715, n4730, n4729, n4714, n2516, n5448, n2867, 
        n2866, n2865, n2864, n2863, n2517, n2862, n2861, n2860, 
        n2859, n2858, n2857, n4728, n4727, n2856, n2455, n2855, 
        n2854, n2853, n2852, n2851, n2384, n2850, n2381, n2849, 
        n2380, n2848, n2847, n2846, n2845, n2844, n5479, n2843, 
        n2842, n2841, n2840, n2839, n2838, n2837, n2836, n2523, 
        n2835, n2834, n2833, n2830, n135_adj_1974, n134, n133, 
        n132, n131, n130, n129, n128, n127, n126, n125, n124, 
        n123, n122, n121, n120, n119, n118, n117, n116, n115, 
        n114, n113, n112, n111, n2478, n2829, n2828, n2827, 
        n2826, n2825, n110, n2824, n4_adj_1975, n2822, n5;
    wire [7:0]i_Tx_Byte;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(18[16:25])
    
    wire n26, n25, n24, n4_adj_1976, n2518, n4544, n23, n22, 
        n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, 
        n11, n10, n9, n8, n4713, n2506, n4726, n4712, n2507, 
        n21_adj_1977, n4725, n7, n6, n4724, n2514, n2661, n2660, 
        n2659, n2658, n2657, n2656, n2655, n2654, n2653, n2652, 
        n2651, n2650, n2649, n2648, n2647, n2646, n2645, n2644, 
        n2643, n2642, n2641, n2640, n2639, n2638, n2637, n2636, 
        n2635, n2634, n2633, n2632, n2631, n2630, n2629, n2628, 
        n2627, n2626, n2625, n2624, n2623, n2622, n2621, n2620, 
        n2619, n2618, n2617, n2616, n2615, n2614, n2613, n2612, 
        n2611, n2610, n2609, n2608, n2607, n2606, n2605, n2604, 
        n2603, n2602, n2601, n2600, n2599, n2598, n2597, n2596, 
        n2595, n2594, n2593, n2592, n2591, n2590, n2589, n2588, 
        n2587, n2586, n2585, n2584, n2583, n2582, n2581, n2580, 
        n2579, n2578, n2577, n2576, n2575, n2574, n2573, n2572, 
        n2571, n2570, n2569, n2568, n2567, n2566, n2565, n2564, 
        n2563, n2562, n2561, n2560, n2559, n2558, n2557, n2556, 
        n2555, n2554, n2553, n2552, n2551, n2550, n2549, n2548, 
        n2547, n2546, n2545, n2544, n2543, n2542, n2541, n2540, 
        n2539, n2538, n2537, n2536, n2535, n2534, n2533, n2532, 
        n2531, n2530, n2529, n2450, n2447, n2339, n2476, n2208, 
        n2470, n2198, n5440, n5355, n5415, n2513, n2515, n4_adj_1978, 
        n11_adj_1979, n5111, n4723, n5400, n5089, n4711, n4_adj_1980, 
        n5482, n2509, n1764, n2467, n4_adj_1981, n1991, n4_adj_1982, 
        n1757, tx_active, n4155;
    wire [2:0]r_SM_Main;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    wire [7:0]r_Tx_Data;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(34[16:25])
    
    wire n4_adj_1983, n313, n315, n4722, n8_adj_1984, n7_adj_1985, 
        n4_adj_1986, n8_adj_1987, n7_adj_1988, n2418, n2415, n317, 
        n318, n320, n321, r_Rx_Data;
    wire [2:0]r_Bit_Index_adj_1999;   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_adj_2000;   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(36[17:26])
    
    wire n1768, n5646;
    wire [2:0]r_SM_Main_2__N_1824;
    
    wire n5871;
    wire [2:0]r_SM_Main_adj_2003;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_2004;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index_adj_2005;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(33[16:27])
    
    wire n4_adj_1996, n1760, n313_adj_1997, n1579, n4721, n5364, 
        n5645, n782, n4710;
    
    VCC i2 (.Y(VCC_net));
    SB_IO tx2_output (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx2_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx2_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx2_output.PIN_TYPE = 6'b101001;
    defparam tx2_output.PULLUP = 1'b1;
    defparam tx2_output.NEG_TRIGGER = 1'b0;
    defparam tx2_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO rx_input (.PACKAGE_PIN(PIN_2), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), .D_OUT_1(GND_net), 
          .D_OUT_0(GND_net), .D_IN_0(rx_i)) /* synthesis lattice_noprune=1, syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam rx_input.PIN_TYPE = 6'b000001;
    defparam rx_input.PULLUP = 1'b1;
    defparam rx_input.NEG_TRIGGER = 1'b0;
    defparam rx_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_1), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF blink_counter_523__i0 (.Q(n26), .C(CLK_c), .D(n135_adj_1974));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 i2583_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_1980), 
            .I3(n1764), .O(n2834));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i2583_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2227_4_lut (.I0(tx_active), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n5), .O(n2478));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2227_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i2129_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4), .I3(n1760), 
            .O(n2380));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i2129_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2573_3_lut (.I0(r_Tx_Data[1]), .I1(i_Tx_Byte[1]), .I2(n1519), 
            .I3(GND_net), .O(n2824));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2130_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(r_Bit_Index_adj_1999[0]), 
            .I3(n1757), .O(n2381));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i2130_4_lut.LUT_INIT = 16'hccac;
    SB_DFF blink_counter_523__i25 (.Q(blink_counter[25]), .C(CLK_c), .D(n110));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 i2602_4_lut (.I0(\data_out[18] [1]), .I1(n4_adj_1983), .I2(n4334), 
            .I3(n5421), .O(n2853));   // coms.v(123[10] 164[6])
    defparam i2602_4_lut.LUT_INIT = 16'ha3ac;
    SB_LUT4 i2241_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2492));   // coms.v(174[10] 182[6])
    defparam i2241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2219_4_lut (.I0(n782), .I1(r_Clock_Count[3]), .I2(n318), 
            .I3(r_SM_Main[2]), .O(n2470));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2219_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 blink_counter_523_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[25]), .I3(n4734), .O(n110)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2601_4_lut (.I0(\data_out[18] [0]), .I1(n5364), .I2(n4334), 
            .I3(\data_out[10] [2]), .O(n2852));   // coms.v(123[10] 164[6])
    defparam i2601_4_lut.LUT_INIT = 16'ha3ac;
    SB_LUT4 i2216_4_lut (.I0(n782), .I1(r_Clock_Count[4]), .I2(n317), 
            .I3(r_SM_Main[2]), .O(n2467));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2216_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i2253_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2504));   // coms.v(174[10] 182[6])
    defparam i2253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2254_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2505));   // coms.v(174[10] 182[6])
    defparam i2254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2255_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2506));   // coms.v(174[10] 182[6])
    defparam i2255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2256_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2507));   // coms.v(174[10] 182[6])
    defparam i2256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2257_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2508));   // coms.v(174[10] 182[6])
    defparam i2257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2258_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2509));   // coms.v(174[10] 182[6])
    defparam i2258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[24]), .I3(n4733), .O(n111)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2259_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2510));   // coms.v(174[10] 182[6])
    defparam i2259_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_3 (.CI(n4710), .I0(GND_net), .I1(n25), 
            .CO(n4711));
    SB_LUT4 i2603_4_lut (.I0(\data_out[18] [2]), .I1(n5424), .I2(n4334), 
            .I3(n5479), .O(n2854));   // coms.v(123[10] 164[6])
    defparam i2603_4_lut.LUT_INIT = 16'ha3ac;
    SB_LUT4 blink_counter_523_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n26), 
            .I3(VCC_net), .O(n135_adj_1974)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2615_4_lut (.I0(\data_out[19] [6]), .I1(n4_adj_1986), .I2(n4334), 
            .I3(n5400), .O(n2866));   // coms.v(123[10] 164[6])
    defparam i2615_4_lut.LUT_INIT = 16'ha3ac;
    SB_LUT4 i2271_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2522));   // coms.v(174[10] 182[6])
    defparam i2271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2272_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2523));   // coms.v(174[10] 182[6])
    defparam i2272_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_14 (.CI(n4721), .I0(GND_net), .I1(n14), 
            .CO(n4722));
    SB_CARRY blink_counter_523_add_4_26 (.CI(n4733), .I0(GND_net), .I1(blink_counter[24]), 
            .CO(n4734));
    SB_LUT4 i2273_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2524));   // coms.v(174[10] 182[6])
    defparam i2273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15), .I3(n4720), .O(n124)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2577_3_lut (.I0(r_Tx_Data[5]), .I1(i_Tx_Byte[5]), .I2(n1519), 
            .I3(GND_net), .O(n2828));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2577_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_13 (.CI(n4720), .I0(GND_net), .I1(n15), 
            .CO(n4721));
    SB_LUT4 i2196_4_lut (.I0(n782), .I1(r_Clock_Count[0]), .I2(n321), 
            .I3(r_SM_Main[2]), .O(n2447));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2196_4_lut.LUT_INIT = 16'h4450;
    SB_CARRY blink_counter_523_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n26), 
            .CO(n4710));
    SB_LUT4 blink_counter_523_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[23]), .I3(n4732), .O(n112)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2604_4_lut (.I0(\data_out[18] [3]), .I1(n1579), .I2(n4334), 
            .I3(n5433), .O(n2855));   // coms.v(123[10] 164[6])
    defparam i2604_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i2133_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2384));   // coms.v(174[10] 182[6])
    defparam i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2260_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2511));   // coms.v(174[10] 182[6])
    defparam i2260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2578_3_lut (.I0(r_Tx_Data[6]), .I1(i_Tx_Byte[6]), .I2(n1519), 
            .I3(GND_net), .O(n2829));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2578_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF blink_counter_523__i24 (.Q(blink_counter[24]), .C(CLK_c), .D(n111));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i23 (.Q(blink_counter[23]), .C(CLK_c), .D(n112));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i22 (.Q(blink_counter[22]), .C(CLK_c), .D(n113));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i21 (.Q(blink_counter[21]), .C(CLK_c), .D(n114));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i20 (.Q(n6), .C(CLK_c), .D(n115));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i19 (.Q(n7), .C(CLK_c), .D(n116));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i18 (.Q(n8), .C(CLK_c), .D(n117));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i17 (.Q(n9), .C(CLK_c), .D(n118));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i16 (.Q(n10), .C(CLK_c), .D(n119));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i15 (.Q(n11), .C(CLK_c), .D(n120));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i14 (.Q(n12), .C(CLK_c), .D(n121));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 i2574_3_lut (.I0(r_Tx_Data[2]), .I1(i_Tx_Byte[2]), .I2(n1519), 
            .I3(GND_net), .O(n2825));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2574_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF blink_counter_523__i13 (.Q(n13), .C(CLK_c), .D(n122));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i12 (.Q(n14), .C(CLK_c), .D(n123));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i11 (.Q(n15), .C(CLK_c), .D(n124));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i10 (.Q(n16), .C(CLK_c), .D(n125));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i9 (.Q(n17), .C(CLK_c), .D(n126));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i8 (.Q(n18), .C(CLK_c), .D(n127));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i7 (.Q(n19), .C(CLK_c), .D(n128));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i6 (.Q(n20), .C(CLK_c), .D(n129));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i5 (.Q(n21), .C(CLK_c), .D(n130));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i4 (.Q(n22), .C(CLK_c), .D(n131));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i3 (.Q(n23), .C(CLK_c), .D(n132));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i2 (.Q(n24), .C(CLK_c), .D(n133));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_DFF blink_counter_523__i1 (.Q(n25), .C(CLK_c), .D(n134));   // verilog/TinyFPGA_B.v(71[24:41])
    SB_LUT4 i2576_3_lut (.I0(r_Tx_Data[4]), .I1(i_Tx_Byte[4]), .I2(n1519), 
            .I3(GND_net), .O(n2827));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16), .I3(n4719), .O(n125)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5300_4_lut (.I0(blink_counter[22]), .I1(blink_counter[23]), 
            .I2(blink_counter[24]), .I3(blink_counter[21]), .O(n5646));
    defparam i5300_4_lut.LUT_INIT = 16'hfec4;
    SB_LUT4 i5299_4_lut (.I0(blink_counter[23]), .I1(blink_counter[22]), 
            .I2(blink_counter[24]), .I3(blink_counter[21]), .O(n5645));
    defparam i5299_4_lut.LUT_INIT = 16'hcf08;
    SB_LUT4 i2575_3_lut (.I0(r_Tx_Data[3]), .I1(i_Tx_Byte[3]), .I2(n1519), 
            .I3(GND_net), .O(n2826));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5301_3_lut (.I0(n5645), .I1(n5646), .I2(blink_counter[25]), 
            .I3(GND_net), .O(LED_c));
    defparam i5301_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY blink_counter_523_add_4_12 (.CI(n4719), .I0(GND_net), .I1(n16), 
            .CO(n4720));
    SB_LUT4 i2605_4_lut (.I0(\data_out[18] [4]), .I1(n1768), .I2(n4334), 
            .I3(n4_adj_1981), .O(n2856));   // coms.v(123[10] 164[6])
    defparam i2605_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i2586_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4), .I3(n1764), 
            .O(n2837));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i2586_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2261_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2512));   // coms.v(174[10] 182[6])
    defparam i2261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2585_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_1980), 
            .I3(n1760), .O(n2836));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i2585_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 blink_counter_523_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17), .I3(n4718), .O(n126)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_523_add_4_25 (.CI(n4732), .I0(GND_net), .I1(blink_counter[23]), 
            .CO(n4733));
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY blink_counter_523_add_4_11 (.CI(n4718), .I0(GND_net), .I1(n17), 
            .CO(n4719));
    SB_LUT4 i2274_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2525));   // coms.v(174[10] 182[6])
    defparam i2274_3_lut.LUT_INIT = 16'hcaca;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i2262_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2513));   // coms.v(174[10] 182[6])
    defparam i2262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2263_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2514));   // coms.v(174[10] 182[6])
    defparam i2263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2264_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2515));   // coms.v(174[10] 182[6])
    defparam i2264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2571_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n3636), 
            .I3(n1764), .O(n2822));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i2571_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i2579_3_lut (.I0(r_Tx_Data[7]), .I1(i_Tx_Byte[7]), .I2(n1519), 
            .I3(GND_net), .O(n2830));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2265_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2516));   // coms.v(174[10] 182[6])
    defparam i2265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2266_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2517));   // coms.v(174[10] 182[6])
    defparam i2266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2606_4_lut (.I0(\data_out[18] [5]), .I1(n4_adj_1996), .I2(n4334), 
            .I3(n5433), .O(n2857));   // coms.v(123[10] 164[6])
    defparam i2606_4_lut.LUT_INIT = 16'ha3ac;
    SB_LUT4 i2235_4_lut (.I0(tx2_active), .I1(r_SM_Main_adj_2003[1]), .I2(r_SM_Main_adj_2003[2]), 
            .I3(n4_adj_1973), .O(n2486));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2235_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i2609_4_lut (.I0(\data_out[19] [0]), .I1(n7_adj_1988), .I2(n4334), 
            .I3(n8_adj_1987), .O(n2860));   // coms.v(123[10] 164[6])
    defparam i2609_4_lut.LUT_INIT = 16'ha3ac;
    SB_LUT4 i2267_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2518));   // coms.v(174[10] 182[6])
    defparam i2267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2607_4_lut (.I0(\data_out[18] [6]), .I1(\data_out[10] [4]), 
            .I2(n4334), .I3(n4_adj_1976), .O(n2858));   // coms.v(123[10] 164[6])
    defparam i2607_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 blink_counter_523_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[22]), .I3(n4731), .O(n113)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_523_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18), .I3(n4717), .O(n127)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_523_add_4_24 (.CI(n4731), .I0(GND_net), .I1(blink_counter[22]), 
            .CO(n4732));
    SB_LUT4 i5552_4_lut (.I0(\data_out[10] [5]), .I1(n5364), .I2(n1768), 
            .I3(n5482), .O(n5871));   // coms.v(123[10] 164[6])
    defparam i5552_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main_adj_2000[2]), .I1(r_SM_Main_adj_2000[1]), 
            .I2(n2198), .I3(rx_data_ready), .O(n5089));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_SM_Main_adj_2000[2]), .I1(r_SM_Main_adj_2000[1]), 
            .I2(r_SM_Main_adj_2000[0]), .I3(r_SM_Main_2__N_1824[2]), .O(n5355));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i2612_4_lut (.I0(\data_out[19] [3]), .I1(n1991), .I2(n4334), 
            .I3(n5440), .O(n2863));   // coms.v(123[10] 164[6])
    defparam i2612_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i2268_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2519));   // coms.v(174[10] 182[6])
    defparam i2268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2275_3_lut (.I0(\data_in[3] [0]), .I1(\data_in[4] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2526));   // coms.v(174[10] 182[6])
    defparam i2275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2297_3_lut (.I0(\data_in[5] [6]), .I1(\data_in[6] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2548));   // coms.v(174[10] 182[6])
    defparam i2297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2303_3_lut (.I0(\data_in[6] [4]), .I1(\data_in[7] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2554));   // coms.v(174[10] 182[6])
    defparam i2303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2302_3_lut (.I0(\data_in[6] [3]), .I1(\data_in[7] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2553));   // coms.v(174[10] 182[6])
    defparam i2302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2301_3_lut (.I0(\data_in[6] [2]), .I1(\data_in[7] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2552));   // coms.v(174[10] 182[6])
    defparam i2301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2300_3_lut (.I0(\data_in[6] [1]), .I1(\data_in[7] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2551));   // coms.v(174[10] 182[6])
    defparam i2300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2299_3_lut (.I0(\data_in[6] [0]), .I1(\data_in[7] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2550));   // coms.v(174[10] 182[6])
    defparam i2299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2298_3_lut (.I0(\data_in[5] [7]), .I1(\data_in[6] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2549));   // coms.v(174[10] 182[6])
    defparam i2298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2269_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2520));   // coms.v(174[10] 182[6])
    defparam i2269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2616_4_lut (.I0(\data_out[19] [7]), .I1(n135), .I2(n4334), 
            .I3(n5482), .O(n2867));   // coms.v(123[10] 164[6])
    defparam i2616_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i2337_3_lut (.I0(\data_in[10] [6]), .I1(\data_in[11] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2588));   // coms.v(174[10] 182[6])
    defparam i2337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2370_3_lut (.I0(\data_in[14] [7]), .I1(\data_in[15] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2621));   // coms.v(174[10] 182[6])
    defparam i2370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(blink_counter[21]), .I3(n4730), .O(n114)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_523_add_4_23 (.CI(n4730), .I0(GND_net), .I1(blink_counter[21]), 
            .CO(n4731));
    SB_LUT4 i2376_3_lut (.I0(\data_in[15] [5]), .I1(\data_in[16] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2627));   // coms.v(174[10] 182[6])
    defparam i2376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2375_3_lut (.I0(\data_in[15] [4]), .I1(\data_in[16] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2626));   // coms.v(174[10] 182[6])
    defparam i2375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2374_3_lut (.I0(\data_in[15] [3]), .I1(\data_in[16] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2625));   // coms.v(174[10] 182[6])
    defparam i2374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6), .I3(n4729), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_3_lut_4_lut_4_lut (.I0(r_SM_Main_adj_2000[2]), .I1(r_SM_Main_adj_2000[1]), 
            .I2(r_SM_Main_adj_2000[0]), .I3(r_SM_Main_2__N_1824[2]), .O(n2198));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i13_3_lut_4_lut_4_lut.LUT_INIT = 16'h4303;
    SB_LUT4 i2373_3_lut (.I0(\data_in[15] [2]), .I1(\data_in[16] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2624));   // coms.v(174[10] 182[6])
    defparam i2373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2372_3_lut (.I0(\data_in[15] [1]), .I1(\data_in[16] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2623));   // coms.v(174[10] 182[6])
    defparam i2372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2610_4_lut (.I0(\data_out[19] [1]), .I1(n7_adj_1985), .I2(n4334), 
            .I3(n8_adj_1984), .O(n2861));   // coms.v(123[10] 164[6])
    defparam i2610_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i2613_4_lut (.I0(\data_out[19] [4]), .I1(n4_adj_1975), .I2(n4334), 
            .I3(n5448), .O(n2864));   // coms.v(123[10] 164[6])
    defparam i2613_4_lut.LUT_INIT = 16'ha3ac;
    SB_LUT4 i2611_4_lut (.I0(\data_out[19] [2]), .I1(n4_adj_1982), .I2(n4334), 
            .I3(n5440), .O(n2862));   // coms.v(123[10] 164[6])
    defparam i2611_4_lut.LUT_INIT = 16'ha3ac;
    SB_LUT4 i2371_3_lut (.I0(\data_in[15] [0]), .I1(\data_in[16] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2622));   // coms.v(174[10] 182[6])
    defparam i2371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2614_4_lut (.I0(\data_out[19] [5]), .I1(n4_adj_1978), .I2(n4334), 
            .I3(n5415), .O(n2865));   // coms.v(123[10] 164[6])
    defparam i2614_4_lut.LUT_INIT = 16'ha3ac;
    SB_LUT4 i2407_3_lut (.I0(\data_in[19] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2658));   // coms.v(174[10] 182[6])
    defparam i2407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2406_3_lut (.I0(\data_in[19] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2657));   // coms.v(174[10] 182[6])
    defparam i2406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2405_3_lut (.I0(\data_in[19] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2656));   // coms.v(174[10] 182[6])
    defparam i2405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2404_3_lut (.I0(\data_in[19] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2655));   // coms.v(174[10] 182[6])
    defparam i2404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2403_3_lut (.I0(\data_in[19] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2654));   // coms.v(174[10] 182[6])
    defparam i2403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2402_3_lut (.I0(\data_in[18] [7]), .I1(\data_in[19] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2653));   // coms.v(174[10] 182[6])
    defparam i2402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2401_3_lut (.I0(\data_in[18] [6]), .I1(\data_in[19] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2652));   // coms.v(174[10] 182[6])
    defparam i2401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2400_3_lut (.I0(\data_in[18] [5]), .I1(\data_in[19] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2651));   // coms.v(174[10] 182[6])
    defparam i2400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2399_3_lut (.I0(\data_in[18] [4]), .I1(\data_in[19] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2650));   // coms.v(174[10] 182[6])
    defparam i2399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2398_3_lut (.I0(\data_in[18] [3]), .I1(\data_in[19] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2649));   // coms.v(174[10] 182[6])
    defparam i2398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2397_3_lut (.I0(\data_in[18] [2]), .I1(\data_in[19] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2648));   // coms.v(174[10] 182[6])
    defparam i2397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2396_3_lut (.I0(\data_in[18] [1]), .I1(\data_in[19] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2647));   // coms.v(174[10] 182[6])
    defparam i2396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2395_3_lut (.I0(\data_in[18] [0]), .I1(\data_in[19] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2646));   // coms.v(174[10] 182[6])
    defparam i2395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2394_3_lut (.I0(\data_in[17] [7]), .I1(\data_in[18] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2645));   // coms.v(174[10] 182[6])
    defparam i2394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2393_3_lut (.I0(\data_in[17] [6]), .I1(\data_in[18] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2644));   // coms.v(174[10] 182[6])
    defparam i2393_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_10 (.CI(n4717), .I0(GND_net), .I1(n18), 
            .CO(n4718));
    SB_LUT4 i2392_3_lut (.I0(\data_in[17] [5]), .I1(\data_in[18] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2643));   // coms.v(174[10] 182[6])
    defparam i2392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2391_3_lut (.I0(\data_in[17] [4]), .I1(\data_in[18] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2642));   // coms.v(174[10] 182[6])
    defparam i2391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2390_3_lut (.I0(\data_in[17] [3]), .I1(\data_in[18] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2641));   // coms.v(174[10] 182[6])
    defparam i2390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2389_3_lut (.I0(\data_in[17] [2]), .I1(\data_in[18] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2640));   // coms.v(174[10] 182[6])
    defparam i2389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2388_3_lut (.I0(\data_in[17] [1]), .I1(\data_in[18] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2639));   // coms.v(174[10] 182[6])
    defparam i2388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2387_3_lut (.I0(\data_in[17] [0]), .I1(\data_in[18] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2638));   // coms.v(174[10] 182[6])
    defparam i2387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2386_3_lut (.I0(\data_in[16] [7]), .I1(\data_in[17] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2637));   // coms.v(174[10] 182[6])
    defparam i2386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2385_3_lut (.I0(\data_in[16] [6]), .I1(\data_in[17] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2636));   // coms.v(174[10] 182[6])
    defparam i2385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2384_3_lut (.I0(\data_in[16] [5]), .I1(\data_in[17] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2635));   // coms.v(174[10] 182[6])
    defparam i2384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2383_3_lut (.I0(\data_in[16] [4]), .I1(\data_in[17] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2634));   // coms.v(174[10] 182[6])
    defparam i2383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2382_3_lut (.I0(\data_in[16] [3]), .I1(\data_in[17] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2633));   // coms.v(174[10] 182[6])
    defparam i2382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2381_3_lut (.I0(\data_in[16] [2]), .I1(\data_in[17] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2632));   // coms.v(174[10] 182[6])
    defparam i2381_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_22 (.CI(n4729), .I0(GND_net), .I1(n6), 
            .CO(n4730));
    SB_LUT4 i2380_3_lut (.I0(\data_in[16] [1]), .I1(\data_in[17] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2631));   // coms.v(174[10] 182[6])
    defparam i2380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2408_3_lut (.I0(\data_in[19] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2659));   // coms.v(174[10] 182[6])
    defparam i2408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2379_3_lut (.I0(\data_in[16] [0]), .I1(\data_in[17] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2630));   // coms.v(174[10] 182[6])
    defparam i2379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2378_3_lut (.I0(\data_in[15] [7]), .I1(\data_in[16] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2629));   // coms.v(174[10] 182[6])
    defparam i2378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7), .I3(n4728), .O(n116)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2377_3_lut (.I0(\data_in[15] [6]), .I1(\data_in[16] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2628));   // coms.v(174[10] 182[6])
    defparam i2377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2369_3_lut (.I0(\data_in[14] [6]), .I1(\data_in[15] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2620));   // coms.v(174[10] 182[6])
    defparam i2369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2368_3_lut (.I0(\data_in[14] [5]), .I1(\data_in[15] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2619));   // coms.v(174[10] 182[6])
    defparam i2368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2367_3_lut (.I0(\data_in[14] [4]), .I1(\data_in[15] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2618));   // coms.v(174[10] 182[6])
    defparam i2367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2582_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n3636), 
            .I3(n1760), .O(n2833));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i2582_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i2366_3_lut (.I0(\data_in[14] [3]), .I1(\data_in[15] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2617));   // coms.v(174[10] 182[6])
    defparam i2366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2365_3_lut (.I0(\data_in[14] [2]), .I1(\data_in[15] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2616));   // coms.v(174[10] 182[6])
    defparam i2365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2364_3_lut (.I0(\data_in[14] [1]), .I1(\data_in[15] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2615));   // coms.v(174[10] 182[6])
    defparam i2364_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_21 (.CI(n4728), .I0(GND_net), .I1(n7), 
            .CO(n4729));
    SB_LUT4 blink_counter_523_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8), .I3(n4727), .O(n117)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_523_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(n19), 
            .I3(n4716), .O(n128)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_523_add_4_9 (.CI(n4716), .I0(GND_net), .I1(n19), 
            .CO(n4717));
    SB_LUT4 blink_counter_523_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(n20), 
            .I3(n4715), .O(n129)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_523_add_4_20 (.CI(n4727), .I0(GND_net), .I1(n8), 
            .CO(n4728));
    SB_LUT4 i2363_3_lut (.I0(\data_in[14] [0]), .I1(\data_in[15] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2614));   // coms.v(174[10] 182[6])
    defparam i2363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9), .I3(n4726), .O(n118)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2362_3_lut (.I0(\data_in[13] [7]), .I1(\data_in[14] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2613));   // coms.v(174[10] 182[6])
    defparam i2362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2361_3_lut (.I0(\data_in[13] [6]), .I1(\data_in[14] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2612));   // coms.v(174[10] 182[6])
    defparam i2361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2360_3_lut (.I0(\data_in[13] [5]), .I1(\data_in[14] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2611));   // coms.v(174[10] 182[6])
    defparam i2360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2359_3_lut (.I0(\data_in[13] [4]), .I1(\data_in[14] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2610));   // coms.v(174[10] 182[6])
    defparam i2359_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_19 (.CI(n4726), .I0(GND_net), .I1(n9), 
            .CO(n4727));
    SB_CARRY blink_counter_523_add_4_8 (.CI(n4715), .I0(GND_net), .I1(n20), 
            .CO(n4716));
    SB_LUT4 blink_counter_523_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(n21), 
            .I3(n4714), .O(n130)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2358_3_lut (.I0(\data_in[13] [3]), .I1(\data_in[14] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2609));   // coms.v(174[10] 182[6])
    defparam i2358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2357_3_lut (.I0(\data_in[13] [2]), .I1(\data_in[14] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2608));   // coms.v(174[10] 182[6])
    defparam i2357_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_7 (.CI(n4714), .I0(GND_net), .I1(n21), 
            .CO(n4715));
    SB_LUT4 blink_counter_523_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10), .I3(n4725), .O(n119)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2356_3_lut (.I0(\data_in[13] [1]), .I1(\data_in[14] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2607));   // coms.v(174[10] 182[6])
    defparam i2356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2355_3_lut (.I0(\data_in[13] [0]), .I1(\data_in[14] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2606));   // coms.v(174[10] 182[6])
    defparam i2355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2354_3_lut (.I0(\data_in[12] [7]), .I1(\data_in[13] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2605));   // coms.v(174[10] 182[6])
    defparam i2354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2353_3_lut (.I0(\data_in[12] [6]), .I1(\data_in[13] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2604));   // coms.v(174[10] 182[6])
    defparam i2353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2352_3_lut (.I0(\data_in[12] [5]), .I1(\data_in[13] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2603));   // coms.v(174[10] 182[6])
    defparam i2352_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_18 (.CI(n4725), .I0(GND_net), .I1(n10), 
            .CO(n4726));
    SB_LUT4 i2351_3_lut (.I0(\data_in[12] [4]), .I1(\data_in[13] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2602));   // coms.v(174[10] 182[6])
    defparam i2351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2350_3_lut (.I0(\data_in[12] [3]), .I1(\data_in[13] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2601));   // coms.v(174[10] 182[6])
    defparam i2350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2349_3_lut (.I0(\data_in[12] [2]), .I1(\data_in[13] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2600));   // coms.v(174[10] 182[6])
    defparam i2349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2410_3_lut (.I0(\data_in[19] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2661));   // coms.v(174[10] 182[6])
    defparam i2410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2348_3_lut (.I0(\data_in[12] [1]), .I1(\data_in[13] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2599));   // coms.v(174[10] 182[6])
    defparam i2348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2409_3_lut (.I0(\data_in[19] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2660));   // coms.v(174[10] 182[6])
    defparam i2409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2347_3_lut (.I0(\data_in[12] [0]), .I1(\data_in[13] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2598));   // coms.v(174[10] 182[6])
    defparam i2347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2346_3_lut (.I0(\data_in[11] [7]), .I1(\data_in[12] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2597));   // coms.v(174[10] 182[6])
    defparam i2346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2588_3_lut_4_lut (.I0(\data_out[10] [3]), .I1(data[11]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2839));   // coms.v(123[10] 164[6])
    defparam i2588_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2345_3_lut (.I0(\data_in[11] [6]), .I1(\data_in[12] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2596));   // coms.v(174[10] 182[6])
    defparam i2345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2344_3_lut (.I0(\data_in[11] [5]), .I1(\data_in[12] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2595));   // coms.v(174[10] 182[6])
    defparam i2344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2343_3_lut (.I0(\data_in[11] [4]), .I1(\data_in[12] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2594));   // coms.v(174[10] 182[6])
    defparam i2343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2342_3_lut (.I0(\data_in[11] [3]), .I1(\data_in[12] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2593));   // coms.v(174[10] 182[6])
    defparam i2342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2341_3_lut (.I0(\data_in[11] [2]), .I1(\data_in[12] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2592));   // coms.v(174[10] 182[6])
    defparam i2341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2608_3_lut_4_lut (.I0(\data_out[18] [7]), .I1(n5871), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2859));   // coms.v(123[10] 164[6])
    defparam i2608_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2340_3_lut (.I0(\data_in[11] [1]), .I1(\data_in[12] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2591));   // coms.v(174[10] 182[6])
    defparam i2340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2339_3_lut (.I0(\data_in[11] [0]), .I1(\data_in[12] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2590));   // coms.v(174[10] 182[6])
    defparam i2339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2338_3_lut (.I0(\data_in[10] [7]), .I1(\data_in[11] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2589));   // coms.v(174[10] 182[6])
    defparam i2338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2336_3_lut (.I0(\data_in[10] [5]), .I1(\data_in[11] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2587));   // coms.v(174[10] 182[6])
    defparam i2336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2335_3_lut (.I0(\data_in[10] [4]), .I1(\data_in[11] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2586));   // coms.v(174[10] 182[6])
    defparam i2335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2334_3_lut (.I0(\data_in[10] [3]), .I1(\data_in[11] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2585));   // coms.v(174[10] 182[6])
    defparam i2334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2333_3_lut (.I0(\data_in[10] [2]), .I1(\data_in[11] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2584));   // coms.v(174[10] 182[6])
    defparam i2333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2332_3_lut (.I0(\data_in[10] [1]), .I1(\data_in[11] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2583));   // coms.v(174[10] 182[6])
    defparam i2332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2331_3_lut (.I0(\data_in[10] [0]), .I1(\data_in[11] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2582));   // coms.v(174[10] 182[6])
    defparam i2331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2330_3_lut (.I0(\data_in[9] [7]), .I1(\data_in[10] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2581));   // coms.v(174[10] 182[6])
    defparam i2330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2329_3_lut (.I0(\data_in[9] [6]), .I1(\data_in[10] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2580));   // coms.v(174[10] 182[6])
    defparam i2329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2328_3_lut (.I0(\data_in[9] [5]), .I1(\data_in[10] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2579));   // coms.v(174[10] 182[6])
    defparam i2328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2199_3_lut (.I0(n2339), .I1(r_Bit_Index_adj_2005[0]), .I2(n2208), 
            .I3(GND_net), .O(n2450));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2199_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i2593_3_lut_4_lut (.I0(\data_out[11] [0]), .I1(data[0]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2844));   // coms.v(123[10] 164[6])
    defparam i2593_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2592_3_lut_4_lut (.I0(\data_out[10] [7]), .I1(data[15]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2843));   // coms.v(123[10] 164[6])
    defparam i2592_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2167_4_lut (.I0(n782), .I1(r_Clock_Count[6]), .I2(n315), 
            .I3(r_SM_Main[2]), .O(n2418));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2167_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_1979));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2137_4_lut (.I0(n782), .I1(r_Clock_Count[8]), .I2(n313), 
            .I3(r_SM_Main[2]), .O(n2388));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2137_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i2270_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2521));   // coms.v(174[10] 182[6])
    defparam i2270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2327_3_lut (.I0(\data_in[9] [4]), .I1(\data_in[10] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2578));   // coms.v(174[10] 182[6])
    defparam i2327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2326_3_lut (.I0(\data_in[9] [3]), .I1(\data_in[10] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2577));   // coms.v(174[10] 182[6])
    defparam i2326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2325_3_lut (.I0(\data_in[9] [2]), .I1(\data_in[10] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2576));   // coms.v(174[10] 182[6])
    defparam i2325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2324_3_lut (.I0(\data_in[9] [1]), .I1(\data_in[10] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2575));   // coms.v(174[10] 182[6])
    defparam i2324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2323_3_lut (.I0(\data_in[9] [0]), .I1(\data_in[10] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2574));   // coms.v(174[10] 182[6])
    defparam i2323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2322_3_lut (.I0(\data_in[8] [7]), .I1(\data_in[9] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2573));   // coms.v(174[10] 182[6])
    defparam i2322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2321_3_lut (.I0(\data_in[8] [6]), .I1(\data_in[9] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2572));   // coms.v(174[10] 182[6])
    defparam i2321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2320_3_lut (.I0(\data_in[8] [5]), .I1(\data_in[9] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2571));   // coms.v(174[10] 182[6])
    defparam i2320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2319_3_lut (.I0(\data_in[8] [4]), .I1(\data_in[9] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2570));   // coms.v(174[10] 182[6])
    defparam i2319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2599_3_lut_4_lut (.I0(\data_out[11] [6]), .I1(data[6]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2850));   // coms.v(123[10] 164[6])
    defparam i2599_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2318_3_lut (.I0(\data_in[8] [3]), .I1(\data_in[9] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2569));   // coms.v(174[10] 182[6])
    defparam i2318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2591_3_lut_4_lut (.I0(\data_out[10] [6]), .I1(data[14]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2842));   // coms.v(123[10] 164[6])
    defparam i2591_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2317_3_lut (.I0(\data_in[8] [2]), .I1(\data_in[9] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2568));   // coms.v(174[10] 182[6])
    defparam i2317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2316_3_lut (.I0(\data_in[8] [1]), .I1(\data_in[9] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2567));   // coms.v(174[10] 182[6])
    defparam i2316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2315_3_lut (.I0(\data_in[8] [0]), .I1(\data_in[9] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2566));   // coms.v(174[10] 182[6])
    defparam i2315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2314_3_lut (.I0(\data_in[7] [7]), .I1(\data_in[8] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2565));   // coms.v(174[10] 182[6])
    defparam i2314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2313_3_lut (.I0(\data_in[7] [6]), .I1(\data_in[8] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2564));   // coms.v(174[10] 182[6])
    defparam i2313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(n22), 
            .I3(n4713), .O(n131)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blink_counter_523_add_4_6 (.CI(n4713), .I0(GND_net), .I1(n22), 
            .CO(n4714));
    SB_LUT4 blink_counter_523_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11), .I3(n4724), .O(n120)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2312_3_lut (.I0(\data_in[7] [5]), .I1(\data_in[8] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2563));   // coms.v(174[10] 182[6])
    defparam i2312_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_17 (.CI(n4724), .I0(GND_net), .I1(n11), 
            .CO(n4725));
    SB_LUT4 i2311_3_lut (.I0(\data_in[7] [4]), .I1(\data_in[8] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2562));   // coms.v(174[10] 182[6])
    defparam i2311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2310_3_lut (.I0(\data_in[7] [3]), .I1(\data_in[8] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2561));   // coms.v(174[10] 182[6])
    defparam i2310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2309_3_lut (.I0(\data_in[7] [2]), .I1(\data_in[8] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2560));   // coms.v(174[10] 182[6])
    defparam i2309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2308_3_lut (.I0(\data_in[7] [1]), .I1(\data_in[8] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2559));   // coms.v(174[10] 182[6])
    defparam i2308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2587_3_lut_4_lut (.I0(\data_out[10] [2]), .I1(data[10]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2838));   // coms.v(123[10] 164[6])
    defparam i2587_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2307_3_lut (.I0(\data_in[7] [0]), .I1(\data_in[8] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2558));   // coms.v(174[10] 182[6])
    defparam i2307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2306_3_lut (.I0(\data_in[6] [7]), .I1(\data_in[7] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2557));   // coms.v(174[10] 182[6])
    defparam i2306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2305_3_lut (.I0(\data_in[6] [6]), .I1(\data_in[7] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2556));   // coms.v(174[10] 182[6])
    defparam i2305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2304_3_lut (.I0(\data_in[6] [5]), .I1(\data_in[7] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2555));   // coms.v(174[10] 182[6])
    defparam i2304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2296_3_lut (.I0(\data_in[5] [5]), .I1(\data_in[6] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2547));   // coms.v(174[10] 182[6])
    defparam i2296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2295_3_lut (.I0(\data_in[5] [4]), .I1(\data_in[6] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2546));   // coms.v(174[10] 182[6])
    defparam i2295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2597_3_lut_4_lut (.I0(\data_out[11] [4]), .I1(data[4]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2848));   // coms.v(123[10] 164[6])
    defparam i2597_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2294_3_lut (.I0(\data_in[5] [3]), .I1(\data_in[6] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2545));   // coms.v(174[10] 182[6])
    defparam i2294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2293_3_lut (.I0(\data_in[5] [2]), .I1(\data_in[6] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2544));   // coms.v(174[10] 182[6])
    defparam i2293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2590_3_lut_4_lut (.I0(\data_out[10] [5]), .I1(data[13]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2841));   // coms.v(123[10] 164[6])
    defparam i2590_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2292_3_lut (.I0(\data_in[5] [1]), .I1(\data_in[6] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2543));   // coms.v(174[10] 182[6])
    defparam i2292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2291_3_lut (.I0(\data_in[5] [0]), .I1(\data_in[6] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2542));   // coms.v(174[10] 182[6])
    defparam i2291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(n23), 
            .I3(n4712), .O(n132)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2290_3_lut (.I0(\data_in[4] [7]), .I1(\data_in[5] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2541));   // coms.v(174[10] 182[6])
    defparam i2290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2289_3_lut (.I0(\data_in[4] [6]), .I1(\data_in[5] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2540));   // coms.v(174[10] 182[6])
    defparam i2289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2288_3_lut (.I0(\data_in[4] [5]), .I1(\data_in[5] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2539));   // coms.v(174[10] 182[6])
    defparam i2288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2287_3_lut (.I0(\data_in[4] [4]), .I1(\data_in[5] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2538));   // coms.v(174[10] 182[6])
    defparam i2287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2286_3_lut (.I0(\data_in[4] [3]), .I1(\data_in[5] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2537));   // coms.v(174[10] 182[6])
    defparam i2286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2285_3_lut (.I0(\data_in[4] [2]), .I1(\data_in[5] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2536));   // coms.v(174[10] 182[6])
    defparam i2285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2284_3_lut (.I0(\data_in[4] [1]), .I1(\data_in[5] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2535));   // coms.v(174[10] 182[6])
    defparam i2284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2283_3_lut (.I0(\data_in[4] [0]), .I1(\data_in[5] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2534));   // coms.v(174[10] 182[6])
    defparam i2283_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_5 (.CI(n4712), .I0(GND_net), .I1(n23), 
            .CO(n4713));
    SB_LUT4 i2282_3_lut (.I0(\data_in[3] [7]), .I1(\data_in[4] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2533));   // coms.v(174[10] 182[6])
    defparam i2282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2281_3_lut (.I0(\data_in[3] [6]), .I1(\data_in[4] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2532));   // coms.v(174[10] 182[6])
    defparam i2281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12), .I3(n4723), .O(n121)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2280_3_lut (.I0(\data_in[3] [5]), .I1(\data_in[4] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2531));   // coms.v(174[10] 182[6])
    defparam i2280_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blink_counter_523_add_4_16 (.CI(n4723), .I0(GND_net), .I1(n12), 
            .CO(n4724));
    SB_LUT4 i2279_3_lut (.I0(\data_in[3] [4]), .I1(\data_in[4] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2530));   // coms.v(174[10] 182[6])
    defparam i2279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 blink_counter_523_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(n24), 
            .I3(n4711), .O(n133)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2278_3_lut (.I0(\data_in[3] [3]), .I1(\data_in[4] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2529));   // coms.v(174[10] 182[6])
    defparam i2278_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 blink_counter_523_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13), .I3(n4722), .O(n122)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2277_3_lut (.I0(\data_in[3] [2]), .I1(\data_in[4] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2528));   // coms.v(174[10] 182[6])
    defparam i2277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2276_3_lut (.I0(\data_in[3] [1]), .I1(\data_in[4] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n2527));   // coms.v(174[10] 182[6])
    defparam i2276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2233_3_lut_4_lut (.I0(\data_out[10] [0]), .I1(data[8]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2484));   // coms.v(123[10] 164[6])
    defparam i2233_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_CARRY blink_counter_523_add_4_4 (.CI(n4711), .I0(GND_net), .I1(n24), 
            .CO(n4712));
    SB_CARRY blink_counter_523_add_4_15 (.CI(n4722), .I0(GND_net), .I1(n13), 
            .CO(n4723));
    SB_LUT4 blink_counter_523_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(n25), 
            .I3(n4710), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 blink_counter_523_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14), .I3(n4721), .O(n123)) /* synthesis syn_instantiated=1 */ ;
    defparam blink_counter_523_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2225_4_lut (.I0(n782), .I1(r_Clock_Count[1]), .I2(n320), 
            .I3(r_SM_Main[2]), .O(n2476));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2225_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 i2596_3_lut_4_lut (.I0(\data_out[11] [3]), .I1(data[3]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2847));   // coms.v(123[10] 164[6])
    defparam i2596_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2589_3_lut_4_lut (.I0(\data_out[10] [4]), .I1(data[12]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2840));   // coms.v(123[10] 164[6])
    defparam i2589_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2164_4_lut (.I0(n4544), .I1(r_Clock_Count_adj_2004[8]), .I2(n313_adj_1997), 
            .I3(r_SM_Main_adj_2003[2]), .O(n2415));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2164_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i2598_3_lut_4_lut (.I0(\data_out[11] [5]), .I1(data[5]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2849));   // coms.v(123[10] 164[6])
    defparam i2598_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_4_lut (.I0(n4155), .I1(n5818), .I2(n11_adj_1979), .I3(r_SM_Main[2]), 
            .O(n5111));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut.LUT_INIT = 16'hafec;
    SB_LUT4 i2600_3_lut_4_lut (.I0(\data_out[11] [7]), .I1(data[7]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2851));   // coms.v(123[10] 164[6])
    defparam i2600_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2584_3_lut_4_lut (.I0(\data_out[10] [1]), .I1(data[9]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2835));   // coms.v(123[10] 164[6])
    defparam i2584_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2595_3_lut_4_lut (.I0(\data_out[11] [2]), .I1(data[2]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2846));   // coms.v(123[10] 164[6])
    defparam i2595_3_lut_4_lut.LUT_INIT = 16'hacaa;
    coms c0 (.CLK_c(CLK_c), .i_Tx_Byte({i_Tx_Byte[7:1], Open_0}), .\data_in[8] ({\data_in[8] }), 
         .GND_net(GND_net), .data({data}), .n2526(n2526), .\data_in[3] ({\data_in[3] }), 
         .n2839(n2839), .\data_out[10] ({\data_out[10] }), .\data_in[19] ({\data_in[19] }), 
         .\data_in[18] ({\data_in[18] }), .n2525(n2525), .\data_in[2] ({\data_in[2] }), 
         .n2524(n2524), .n2523(n2523), .n2522(n2522), .n2521(n2521), 
         .\data_out[11] ({\data_out[11] }), .n2660(n2660), .n2661(n2661), 
         .n2659(n2659), .n4(n4_adj_1986), .n2622(n2622), .\data_in[15] ({\data_in[15] }), 
         .n2623(n2623), .n2624(n2624), .n2625(n2625), .n2626(n2626), 
         .n2627(n2627), .n2621(n2621), .\data_in[14] ({\data_in[14] }), 
         .n2588(n2588), .\data_in[10] ({\data_in[10] }), .n2520(n2520), 
         .n2549(n2549), .\data_in[5] ({\data_in[5] }), .\data_in[7] ({\data_in[7] }), 
         .n2550(n2550), .\data_in[6] ({\data_in[6] }), .n2551(n2551), 
         .n2552(n2552), .n2553(n2553), .n2554(n2554), .n2548(n2548), 
         .n2519(n2519), .n21(n21_adj_1977), .n2518(n2518), .n2838(n2838), 
         .n2848(n2848), .n2847(n2847), .\data_out[18] ({\data_out[18] }), 
         .\data_out[19] ({\data_out[19] }), .n2849(n2849), .n2835(n2835), 
         .n2845(n2845), .n2865(n2865), .n2862(n2862), .n2864(n2864), 
         .n2861(n2861), .n2867(n2867), .n2863(n2863), .n2859(n2859), 
         .n2858(n2858), .n4333(n4333), .n2844(n2844), .n2860(n2860), 
         .n2843(n2843), .n2857(n2857), .n2517(n2517), .\data_in[1] ({\data_in[1] }), 
         .\data_in[4] ({\data_in[4] }), .n2850(n2850), .n2516(n2516), 
         .n2842(n2842), .n2515(n2515), .n2514(n2514), .n2513(n2513), 
         .n2512(n2512), .n4_adj_2(n4_adj_1996), .n5400(n5400), .n8(n8_adj_1987), 
         .n1768(n1768), .n2484(n2484), .n2511(n2511), .n4334(n4334), 
         .n5482(n5482), .\data_in[0] ({\data_in[0] }), .n2527(n2527), 
         .n2528(n2528), .n2529(n2529), .n2530(n2530), .n2531(n2531), 
         .n2532(n2532), .n2533(n2533), .n2534(n2534), .n2535(n2535), 
         .n2536(n2536), .n2537(n2537), .n2538(n2538), .n2539(n2539), 
         .n2540(n2540), .n2541(n2541), .n2542(n2542), .n2543(n2543), 
         .n2544(n2544), .n2545(n2545), .n2546(n2546), .n2547(n2547), 
         .n2555(n2555), .n2556(n2556), .n2557(n2557), .n2558(n2558), 
         .n2559(n2559), .n2560(n2560), .n2561(n2561), .n2562(n2562), 
         .n2563(n2563), .n2564(n2564), .n2565(n2565), .n2566(n2566), 
         .n2567(n2567), .n2568(n2568), .n2569(n2569), .n2570(n2570), 
         .n2571(n2571), .n2572(n2572), .n2573(n2573), .n2574(n2574), 
         .\data_in[9] ({\data_in[9] }), .n2575(n2575), .n2576(n2576), 
         .n2577(n2577), .n2578(n2578), .n2579(n2579), .n2580(n2580), 
         .n2581(n2581), .n2582(n2582), .n2583(n2583), .n2584(n2584), 
         .n2585(n2585), .n2586(n2586), .n2587(n2587), .n2589(n2589), 
         .n2590(n2590), .\data_in[11] ({\data_in[11] }), .n2591(n2591), 
         .n2592(n2592), .n2593(n2593), .n2594(n2594), .n2595(n2595), 
         .n2596(n2596), .n2597(n2597), .n2598(n2598), .\data_in[12] ({\data_in[12] }), 
         .n2599(n2599), .n2600(n2600), .n2601(n2601), .n2602(n2602), 
         .n2603(n2603), .n2604(n2604), .n2605(n2605), .n2606(n2606), 
         .\data_in[13] ({\data_in[13] }), .n2607(n2607), .n2608(n2608), 
         .n2609(n2609), .n2610(n2610), .n2611(n2611), .n2612(n2612), 
         .n2613(n2613), .n2614(n2614), .n2615(n2615), .n2616(n2616), 
         .n2617(n2617), .n2618(n2618), .n2619(n2619), .n2620(n2620), 
         .n2628(n2628), .n2629(n2629), .n2630(n2630), .\data_in[16] ({\data_in[16] }), 
         .n2631(n2631), .n2632(n2632), .n2633(n2633), .n2634(n2634), 
         .n2635(n2635), .n2636(n2636), .n2637(n2637), .n2638(n2638), 
         .\data_in[17] ({\data_in[17] }), .n2639(n2639), .n2640(n2640), 
         .n2641(n2641), .n2642(n2642), .n2643(n2643), .n2644(n2644), 
         .n2645(n2645), .n2646(n2646), .n2647(n2647), .n2648(n2648), 
         .n2649(n2649), .n2650(n2650), .n2651(n2651), .n2652(n2652), 
         .n2653(n2653), .n2654(n2654), .n2655(n2655), .n2656(n2656), 
         .n2657(n2657), .n2658(n2658), .n2841(n2841), .n2856(n2856), 
         .tx_active(tx_active), .tx_o(tx_o), .tx_enable(tx_enable), .n4155(n4155), 
         .n2384(n2384), .n4_adj_3(n4_adj_1982), .n5415(n5415), .n2855(n2855), 
         .n4_adj_4(n4_adj_1978), .n1991(n1991), .n2866(n2866), .n2840(n2840), 
         .n2851(n2851), .n2854(n2854), .n2510(n2510), .n2846(n2846), 
         .n2509(n2509), .n2508(n2508), .n2507(n2507), .n2506(n2506), 
         .n2505(n2505), .n2504(n2504), .n2852(n2852), .n5440(n5440), 
         .n2492(n2492), .n2853(n2853), .n4_adj_5(n4_adj_1975), .n5479(n5479), 
         .n1579(n1579), .VCC_net(VCC_net), .n4_adj_6(n4_adj_1976), .n7(n7_adj_1988), 
         .n5421(n5421), .n5448(n5448), .n135(n135), .tx2_active(tx2_active), 
         .n7_adj_7(n7_adj_1985), .n5364(n5364), .n4_adj_8(n4_adj_1983), 
         .n5424(n5424), .n8_adj_9(n8_adj_1984), .n5433(n5433), .n4_adj_10(n4_adj_1981), 
         .r_SM_Main({r_SM_Main}), .\r_Clock_Count[1] (r_Clock_Count[1]), 
         .n2388(n2388), .\r_Clock_Count[8] (r_Clock_Count[8]), .n2418(n2418), 
         .\r_Clock_Count[6] (r_Clock_Count[6]), .n321(n321), .\r_Clock_Count[0] (r_Clock_Count[0]), 
         .n1519(n1519), .n2826(n2826), .\r_Tx_Data[3] (r_Tx_Data[3]), 
         .n2827(n2827), .\r_Tx_Data[4] (r_Tx_Data[4]), .n2447(n2447), 
         .\r_Tx_Data[1] (r_Tx_Data[1]), .\r_Tx_Data[2] (r_Tx_Data[2]), .n2825(n2825), 
         .n2824(n2824), .n2830(n2830), .\r_Tx_Data[7] (r_Tx_Data[7]), 
         .n2829(n2829), .\r_Tx_Data[6] (r_Tx_Data[6]), .n2478(n2478), 
         .n2476(n2476), .n2828(n2828), .\r_Tx_Data[5] (r_Tx_Data[5]), 
         .\r_Clock_Count[3] (r_Clock_Count[3]), .\r_Clock_Count[4] (r_Clock_Count[4]), 
         .n2467(n2467), .n2470(n2470), .n313(n313), .n315(n315), .n317(n317), 
         .n11(n11_adj_1979), .n782(n782), .n318(n318), .n5111(n5111), 
         .n320(n320), .n5818(n5818), .n5(n5), .n2450(n2450), .\r_Bit_Index[0] (r_Bit_Index_adj_2005[0]), 
         .\r_SM_Main[2]_adj_11 (r_SM_Main_adj_2003[2]), .\r_SM_Main[1]_adj_12 (r_SM_Main_adj_2003[1]), 
         .n4544(n4544), .n2486(n2486), .n313_adj_13(n313_adj_1997), .\r_Clock_Count[8]_adj_14 (r_Clock_Count_adj_2004[8]), 
         .tx2_o(tx2_o), .n4_adj_15(n4_adj_1973), .n2208(n2208), .n2339(n2339), 
         .n2415(n2415), .tx2_enable(tx2_enable), .\r_Bit_Index[0]_adj_16 (r_Bit_Index_adj_1999[0]), 
         .n1757(n1757), .n2836(n2836), .rx_data({rx_data}), .r_SM_Main_adj_22({r_SM_Main_adj_2000}), 
         .\r_SM_Main_2__N_1824[2] (r_SM_Main_2__N_1824[2]), .n2837(n2837), 
         .n2834(n2834), .n2833(n2833), .n1764(n1764), .n4_adj_20(n4), 
         .n5089(n5089), .rx_data_ready(rx_data_ready), .n1760(n1760), 
         .n4_adj_21(n4_adj_1980), .n2822(n2822), .r_Rx_Data(r_Rx_Data), 
         .rx_i(rx_i), .n3636(n3636), .n5355(n5355), .n2381(n2381), .n2380(n2380), 
         .n2455(n2455)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(77[8] 84[4])
    SB_LUT4 i2594_3_lut_4_lut (.I0(\data_out[11] [1]), .I1(data[1]), .I2(n21_adj_1977), 
            .I3(n4333), .O(n2845));   // coms.v(123[10] 164[6])
    defparam i2594_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2204_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(r_Bit_Index_adj_1999[0]), 
            .I3(n1757), .O(n2455));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i2204_4_lut.LUT_INIT = 16'hccca;
    
endmodule
//
// Verilog Description of module coms
//

module coms (CLK_c, i_Tx_Byte, \data_in[8] , GND_net, data, n2526, 
            \data_in[3] , n2839, \data_out[10] , \data_in[19] , \data_in[18] , 
            n2525, \data_in[2] , n2524, n2523, n2522, n2521, \data_out[11] , 
            n2660, n2661, n2659, n4, n2622, \data_in[15] , n2623, 
            n2624, n2625, n2626, n2627, n2621, \data_in[14] , n2588, 
            \data_in[10] , n2520, n2549, \data_in[5] , \data_in[7] , 
            n2550, \data_in[6] , n2551, n2552, n2553, n2554, n2548, 
            n2519, n21, n2518, n2838, n2848, n2847, \data_out[18] , 
            \data_out[19] , n2849, n2835, n2845, n2865, n2862, n2864, 
            n2861, n2867, n2863, n2859, n2858, n4333, n2844, n2860, 
            n2843, n2857, n2517, \data_in[1] , \data_in[4] , n2850, 
            n2516, n2842, n2515, n2514, n2513, n2512, n4_adj_2, 
            n5400, n8, n1768, n2484, n2511, n4334, n5482, \data_in[0] , 
            n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
            n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
            n2543, n2544, n2545, n2546, n2547, n2555, n2556, n2557, 
            n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, 
            n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, 
            n2574, \data_in[9] , n2575, n2576, n2577, n2578, n2579, 
            n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, 
            n2589, n2590, \data_in[11] , n2591, n2592, n2593, n2594, 
            n2595, n2596, n2597, n2598, \data_in[12] , n2599, n2600, 
            n2601, n2602, n2603, n2604, n2605, n2606, \data_in[13] , 
            n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, 
            n2615, n2616, n2617, n2618, n2619, n2620, n2628, n2629, 
            n2630, \data_in[16] , n2631, n2632, n2633, n2634, n2635, 
            n2636, n2637, n2638, \data_in[17] , n2639, n2640, n2641, 
            n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, 
            n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, 
            n2658, n2841, n2856, tx_active, tx_o, tx_enable, n4155, 
            n2384, n4_adj_3, n5415, n2855, n4_adj_4, n1991, n2866, 
            n2840, n2851, n2854, n2510, n2846, n2509, n2508, n2507, 
            n2506, n2505, n2504, n2852, n5440, n2492, n2853, n4_adj_5, 
            n5479, n1579, VCC_net, n4_adj_6, n7, n5421, n5448, 
            n135, tx2_active, n7_adj_7, n5364, n4_adj_8, n5424, 
            n8_adj_9, n5433, n4_adj_10, r_SM_Main, \r_Clock_Count[1] , 
            n2388, \r_Clock_Count[8] , n2418, \r_Clock_Count[6] , n321, 
            \r_Clock_Count[0] , n1519, n2826, \r_Tx_Data[3] , n2827, 
            \r_Tx_Data[4] , n2447, \r_Tx_Data[1] , \r_Tx_Data[2] , n2825, 
            n2824, n2830, \r_Tx_Data[7] , n2829, \r_Tx_Data[6] , n2478, 
            n2476, n2828, \r_Tx_Data[5] , \r_Clock_Count[3] , \r_Clock_Count[4] , 
            n2467, n2470, n313, n315, n317, n11, n782, n318, 
            n5111, n320, n5818, n5, n2450, \r_Bit_Index[0] , \r_SM_Main[2]_adj_11 , 
            \r_SM_Main[1]_adj_12 , n4544, n2486, n313_adj_13, \r_Clock_Count[8]_adj_14 , 
            tx2_o, n4_adj_15, n2208, n2339, n2415, tx2_enable, \r_Bit_Index[0]_adj_16 , 
            n1757, n2836, rx_data, r_SM_Main_adj_22, \r_SM_Main_2__N_1824[2] , 
            n2837, n2834, n2833, n1764, n4_adj_20, n5089, rx_data_ready, 
            n1760, n4_adj_21, n2822, r_Rx_Data, rx_i, n3636, n5355, 
            n2381, n2380, n2455) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input CLK_c;
    output [7:0]i_Tx_Byte;
    output [7:0]\data_in[8] ;
    input GND_net;
    output [15:0]data;
    input n2526;
    output [7:0]\data_in[3] ;
    input n2839;
    output [7:0]\data_out[10] ;
    output [7:0]\data_in[19] ;
    output [7:0]\data_in[18] ;
    input n2525;
    output [7:0]\data_in[2] ;
    input n2524;
    input n2523;
    input n2522;
    input n2521;
    output [7:0]\data_out[11] ;
    input n2660;
    input n2661;
    input n2659;
    output n4;
    input n2622;
    output [7:0]\data_in[15] ;
    input n2623;
    input n2624;
    input n2625;
    input n2626;
    input n2627;
    input n2621;
    output [7:0]\data_in[14] ;
    input n2588;
    output [7:0]\data_in[10] ;
    input n2520;
    input n2549;
    output [7:0]\data_in[5] ;
    output [7:0]\data_in[7] ;
    input n2550;
    output [7:0]\data_in[6] ;
    input n2551;
    input n2552;
    input n2553;
    input n2554;
    input n2548;
    input n2519;
    output n21;
    input n2518;
    input n2838;
    input n2848;
    input n2847;
    output [7:0]\data_out[18] ;
    output [7:0]\data_out[19] ;
    input n2849;
    input n2835;
    input n2845;
    input n2865;
    input n2862;
    input n2864;
    input n2861;
    input n2867;
    input n2863;
    input n2859;
    input n2858;
    output n4333;
    input n2844;
    input n2860;
    input n2843;
    input n2857;
    input n2517;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[4] ;
    input n2850;
    input n2516;
    input n2842;
    input n2515;
    input n2514;
    input n2513;
    input n2512;
    output n4_adj_2;
    output n5400;
    output n8;
    output n1768;
    input n2484;
    input n2511;
    output n4334;
    output n5482;
    output [7:0]\data_in[0] ;
    input n2527;
    input n2528;
    input n2529;
    input n2530;
    input n2531;
    input n2532;
    input n2533;
    input n2534;
    input n2535;
    input n2536;
    input n2537;
    input n2538;
    input n2539;
    input n2540;
    input n2541;
    input n2542;
    input n2543;
    input n2544;
    input n2545;
    input n2546;
    input n2547;
    input n2555;
    input n2556;
    input n2557;
    input n2558;
    input n2559;
    input n2560;
    input n2561;
    input n2562;
    input n2563;
    input n2564;
    input n2565;
    input n2566;
    input n2567;
    input n2568;
    input n2569;
    input n2570;
    input n2571;
    input n2572;
    input n2573;
    input n2574;
    output [7:0]\data_in[9] ;
    input n2575;
    input n2576;
    input n2577;
    input n2578;
    input n2579;
    input n2580;
    input n2581;
    input n2582;
    input n2583;
    input n2584;
    input n2585;
    input n2586;
    input n2587;
    input n2589;
    input n2590;
    output [7:0]\data_in[11] ;
    input n2591;
    input n2592;
    input n2593;
    input n2594;
    input n2595;
    input n2596;
    input n2597;
    input n2598;
    output [7:0]\data_in[12] ;
    input n2599;
    input n2600;
    input n2601;
    input n2602;
    input n2603;
    input n2604;
    input n2605;
    input n2606;
    output [7:0]\data_in[13] ;
    input n2607;
    input n2608;
    input n2609;
    input n2610;
    input n2611;
    input n2612;
    input n2613;
    input n2614;
    input n2615;
    input n2616;
    input n2617;
    input n2618;
    input n2619;
    input n2620;
    input n2628;
    input n2629;
    input n2630;
    output [7:0]\data_in[16] ;
    input n2631;
    input n2632;
    input n2633;
    input n2634;
    input n2635;
    input n2636;
    input n2637;
    input n2638;
    output [7:0]\data_in[17] ;
    input n2639;
    input n2640;
    input n2641;
    input n2642;
    input n2643;
    input n2644;
    input n2645;
    input n2646;
    input n2647;
    input n2648;
    input n2649;
    input n2650;
    input n2651;
    input n2652;
    input n2653;
    input n2654;
    input n2655;
    input n2656;
    input n2657;
    input n2658;
    input n2841;
    input n2856;
    output tx_active;
    output tx_o;
    output tx_enable;
    output n4155;
    input n2384;
    output n4_adj_3;
    output n5415;
    input n2855;
    output n4_adj_4;
    output n1991;
    input n2866;
    input n2840;
    input n2851;
    input n2854;
    input n2510;
    input n2846;
    input n2509;
    input n2508;
    input n2507;
    input n2506;
    input n2505;
    input n2504;
    input n2852;
    output n5440;
    input n2492;
    input n2853;
    output n4_adj_5;
    output n5479;
    output n1579;
    input VCC_net;
    output n4_adj_6;
    output n7;
    output n5421;
    output n5448;
    output n135;
    output tx2_active;
    output n7_adj_7;
    output n5364;
    output n4_adj_8;
    output n5424;
    output n8_adj_9;
    output n5433;
    output n4_adj_10;
    output [2:0]r_SM_Main;
    output \r_Clock_Count[1] ;
    input n2388;
    output \r_Clock_Count[8] ;
    input n2418;
    output \r_Clock_Count[6] ;
    output n321;
    output \r_Clock_Count[0] ;
    output n1519;
    input n2826;
    output \r_Tx_Data[3] ;
    input n2827;
    output \r_Tx_Data[4] ;
    input n2447;
    output \r_Tx_Data[1] ;
    output \r_Tx_Data[2] ;
    input n2825;
    input n2824;
    input n2830;
    output \r_Tx_Data[7] ;
    input n2829;
    output \r_Tx_Data[6] ;
    input n2478;
    input n2476;
    input n2828;
    output \r_Tx_Data[5] ;
    output \r_Clock_Count[3] ;
    output \r_Clock_Count[4] ;
    input n2467;
    input n2470;
    output n313;
    output n315;
    output n317;
    input n11;
    output n782;
    output n318;
    input n5111;
    output n320;
    output n5818;
    output n5;
    input n2450;
    output \r_Bit_Index[0] ;
    output \r_SM_Main[2]_adj_11 ;
    output \r_SM_Main[1]_adj_12 ;
    output n4544;
    input n2486;
    output n313_adj_13;
    output \r_Clock_Count[8]_adj_14 ;
    output tx2_o;
    output n4_adj_15;
    output n2208;
    output n2339;
    input n2415;
    output tx2_enable;
    output \r_Bit_Index[0]_adj_16 ;
    output n1757;
    input n2836;
    output [7:0]rx_data;
    output [2:0]r_SM_Main_adj_22;
    output \r_SM_Main_2__N_1824[2] ;
    input n2837;
    input n2834;
    input n2833;
    output n1764;
    output n4_adj_20;
    input n5089;
    output rx_data_ready;
    output n1760;
    output n4_adj_21;
    input n2822;
    output r_Rx_Data;
    input rx_i;
    output n3636;
    input n5355;
    input n2381;
    input n2380;
    input n2455;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [10:0]n1;
    wire [10:0]delay_counter;   // coms.v(121[13:26])
    
    wire n6135;
    wire [143:0]data_in_field;   // coms.v(113[33:46])
    wire [7:0]byte_transmit_counter2;   // coms.v(185[13:35])
    
    wire n5746, n1729, \FRAME_MATCHER.wait_for_transmission , n2732, 
        n5743, n6129, n4748, n4749;
    wire [15:0]n69;
    
    wire n4747, \FRAME_MATCHER.wait_for_transmission_N_909 , n4735, n5740, 
        n5737, n6132, n2788, n6123, n5752, n2789, n2783, n2784, 
        n2785, n2786, n2787, n6117, n2731, n5755, n5381, n2012, 
        n5403, n20, n6111, n5758, n1979, n2092, n1892, n19, 
        n5500, n18, n2149, n2065, n21_c, n2030, n20_adj_1870, 
        n16, n5491, n5577, n2095, n1908, n2021, n16_adj_1871, 
        n15;
    wire [7:0]tx_transmit_N_568;
    
    wire n81_adj_1872, n95, n2872, n5503, n5443, n5524, n17, n2800, 
        n6105, n16_adj_1873, n2730, n5761, n2873, n6099, n6102, 
        tx_transmit, n106, n4813, n2804, n4763, n4762, n6093, 
        n1948, n5397, n5512, n22, n2729, n2009, n5378, n12, 
        n2728, n2782, n4746, n5767, n2776, n5593, n42, n48, 
        n43, n45, n44, n46, n52, n2777, n2778, n2779, n2780, 
        n2781, n4761, tx_active_prev, n50_adj_1875;
    wire [7:0]byte_transmit_counter;   // coms.v(13[12:33])
    
    wire n5853, n5551, n5557, n5554, n5581, n47, n5488, n1886, 
        n5489, n22_adj_1876, n6087, n5770, n1955, n27;
    wire [7:0]\data_in_frame[18] ;   // coms.v(172[13:26])
    wire [7:0]\data_in_frame[19] ;   // coms.v(172[13:26])
    
    wire n6081, n6084, n4745, n6075, n24, n2775, n5773, n4760, 
        n5375, n30, n24_adj_1877, n32, n6069, n6072, n5536, n20_adj_1878, 
        n5572, n5586, n24_adj_1879, n6063, n5776, n2662, n2664, 
        n2665, n2727, n31, n6057, n1866, n1814, n10, n6060, 
        n6018, n1081;
    wire [7:0]tx2_data;   // coms.v(188[14:22])
    
    wire n2726, n2874, n4744, n2725, n2724, n2723, n16_adj_1880, 
        n2039, n5412, n22_adj_1881, n2722, n4759, n5569, n20_adj_1882, 
        n2875, n2721, n2720, n2107, n24_adj_1884, n5384, n5476, 
        n5427, n5521, n24_adj_1885, n2152, n23, n2719, n5545, 
        n22_adj_1886, n1855, n25, n5466, n5519, n4743, n2718, 
        n2792, n2717, n2716, n2715, n3703, n3689, n6, n5560, 
        n18_adj_1887, n20_adj_1888, n2811, n1926, n5494, n5394, 
        n5527, n19_adj_1889, n22_adj_1890, n2796, n2810, n2714, 
        n9, n1508, n5810, n1198;
    wire [7:0]tx_data;   // coms.v(16[14:21])
    
    wire n9_adj_1891, n5845, n5570, n4709, n2077, n40, n5539, 
        n5548, n45_adj_1892, n2871, n2870, n15_adj_1893, n1251, 
        n2807, n2869, n5388, n44_adj_1894, n34, n48_adj_1895, n2713, 
        n41, n31_adj_1896, n47_adj_1897, n5840, n2293, n13, n5497, 
        n12_adj_1898, n5567, n1253, n5837, n5563, n5590, n49, 
        n5430, n5506, n5575, n14, n1917, n13_adj_1899, n2806, 
        n2712, n37, n35, n31_adj_1900, n32_adj_1901, n5582, n6312, 
        n17_adj_1902, n22_adj_1903, n18_adj_1904, n5542, n5589, n2711, 
        n2710, n2385, n20_adj_1905, n5574, n9_adj_1906, n25_adj_1907, 
        n2709, n2803, n2708, n17_adj_1908, n28, n15_adj_1909, n2802, 
        n27_adj_1910, n29, n4703, n4704, n2707, n2706, n2799, 
        n9_adj_1911, n5833, n2798, n989, n2808, n2705, n31_adj_1912, 
        n17_adj_1913, n22_adj_1914, n5830, n2704, n2703, n2702, 
        n2812, n2701, n2700, n2699, tx2_transmit_N_915;
    wire [2:0]r_SM_Main_2__N_1770;
    
    wire n4758, n2819, n2698, n2697, n2696, n2695, n2694, n2693, 
        n2692, n2691, n2134, n10_adj_1915, n2690, n2068, n6_adj_1917, 
        n6_adj_1918, n2000, n2053, n5454, n18_adj_1919, n6309, n4_adj_1920, 
        n16_adj_1921, n20_adj_1922, n4705, n4706, n1969, n2689, 
        n2074, n2688, n2687, n5469, n2686, n2125, n6_adj_1923, 
        n4708, n2685, n1835, n2104, n1913, n4742, n4757, n2684, 
        n2683, n6039, n4741, n5788, n2682, n2681, n2680, n5509, 
        n4740, n2679, n2678, n22_adj_1924, n2677, n28_adj_1925, 
        n28_adj_1926, n1965, n2676, n2675, n2674, n26, n2143, 
        n5391, n26_adj_1927, n27_adj_1928, n25_adj_1929, n24_adj_1930, 
        n6033, n2673, n2113, n25_adj_1931, n2672, n5791, n4756, 
        n2671, n2666, n2667, n2668, n2669, n2670, n2733, n2734, 
        n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, 
        n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, 
        n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
        n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
        n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, 
        n23_adj_1935, n5372, n2795, n2043, n5409, n4755, n2155, 
        n2794, n6414, n5436, n2101, n18_adj_1938, n2080, n1889, 
        n6027, n6_adj_1939, n5533, n2791, n2790, n1958, n4754, 
        n26_adj_1940, n2821, n6009, n6012, n1779, n1942, n5578, 
        n2489, n5418, n6303, n6306, n30_adj_1941, tx2_transmit_N_1031, 
        n6297, n6300, n2026, n4707, n2818, n2820, n4739, n4753, 
        n4752, n4751, n5369, n6279, n2817, n2062, n6282, n4750, 
        n6273, n5794;
    wire [4:0]n2;
    
    wire n195, n2325, n5686, n6267, n6270, n2056, n5994, n6261, 
        n4738, n6000, n6264, n6255, n5692, n6021, n2089, n6249, 
        n5695, n5797, n6243, n5698, n1973, n5997, n6237, n5701, 
        n6231, n5991, n6234, n6015, n4737, n6225, n6228, n5458, 
        n6219, n5707, n1994, n4795, n25_adj_1948, n5515, n17_adj_1950, 
        n5827, n1249, n6213, n5710, n12_adj_1951, n6207, n5713, 
        n6201, n5716, n6195, n6198, n6189, n36, n4736, n5722, 
        n2816, n6183, n5725, n2793, n6177, n5728, n2797, n6171, 
        n5731, n2801, n2805, n2809, n2813, n2814, n2815, n6165, 
        n6168, n28_adj_1955, n33, n6159, n6153, n14_adj_1957, n6147, 
        n20_adj_1958, n6150, n6141, n18_adj_1959;
    
    SB_DFF delay_counter_528__i2 (.Q(delay_counter[2]), .C(CLK_c), .D(n1[2]));   // coms.v(159[11] 161[5])
    SB_LUT4 n6135_bdd_4_lut (.I0(n6135), .I1(data_in_field[107]), .I2(data_in_field[99]), 
            .I3(byte_transmit_counter2[1]), .O(n5746));
    defparam n6135_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2481_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[8] [6]), .I3(data_in_field[70]), .O(n2732));
    defparam i2481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF delay_counter_528__i1 (.Q(delay_counter[1]), .C(CLK_c), .D(n1[1]));   // coms.v(159[11] 161[5])
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_5789 (.I0(byte_transmit_counter2[2]), 
            .I1(n5743), .I2(n5746), .I3(byte_transmit_counter2[3]), .O(n6129));
    defparam byte_transmit_counter2_2__bdd_4_lut_5789.LUT_INIT = 16'he4aa;
    SB_CARRY data_527_add_4_12 (.CI(n4748), .I0(GND_net), .I1(data[10]), 
            .CO(n4749));
    SB_LUT4 data_527_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(data[9]), 
            .I3(n4747), .O(n69[9])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_527__i15 (.Q(data[15]), .C(CLK_c), .D(n69[15]));   // coms.v(126[13:19])
    SB_DFF data_527__i14 (.Q(data[14]), .C(CLK_c), .D(n69[14]));   // coms.v(126[13:19])
    SB_DFF data_527__i13 (.Q(data[13]), .C(CLK_c), .D(n69[13]));   // coms.v(126[13:19])
    SB_DFF data_527__i12 (.Q(data[12]), .C(CLK_c), .D(n69[12]));   // coms.v(126[13:19])
    SB_DFF data_527__i11 (.Q(data[11]), .C(CLK_c), .D(n69[11]));   // coms.v(126[13:19])
    SB_DFF data_527__i10 (.Q(data[10]), .C(CLK_c), .D(n69[10]));   // coms.v(126[13:19])
    SB_DFF data_527__i9 (.Q(data[9]), .C(CLK_c), .D(n69[9]));   // coms.v(126[13:19])
    SB_DFF data_527__i8 (.Q(data[8]), .C(CLK_c), .D(n69[8]));   // coms.v(126[13:19])
    SB_DFF data_527__i7 (.Q(data[7]), .C(CLK_c), .D(n69[7]));   // coms.v(126[13:19])
    SB_DFF data_527__i6 (.Q(data[6]), .C(CLK_c), .D(n69[6]));   // coms.v(126[13:19])
    SB_DFF data_527__i5 (.Q(data[5]), .C(CLK_c), .D(n69[5]));   // coms.v(126[13:19])
    SB_DFF data_527__i4 (.Q(data[4]), .C(CLK_c), .D(n69[4]));   // coms.v(126[13:19])
    SB_DFF data_527__i3 (.Q(data[3]), .C(CLK_c), .D(n69[3]));   // coms.v(126[13:19])
    SB_DFF data_527__i2 (.Q(data[2]), .C(CLK_c), .D(n69[2]));   // coms.v(126[13:19])
    SB_DFF data_527__i1 (.Q(data[1]), .C(CLK_c), .D(n69[1]));   // coms.v(126[13:19])
    SB_CARRY byte_transmit_counter2_525_526_add_4_2 (.CI(GND_net), .I0(\FRAME_MATCHER.wait_for_transmission_N_909 ), 
            .I1(byte_transmit_counter2[0]), .CO(n4735));
    SB_CARRY data_527_add_4_11 (.CI(n4747), .I0(GND_net), .I1(data[9]), 
            .CO(n4748));
    SB_LUT4 n6129_bdd_4_lut (.I0(n6129), .I1(n5740), .I2(n5737), .I3(byte_transmit_counter2[3]), 
            .O(n6132));
    defparam n6129_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i127 (.Q(data_in_field[126]), .C(CLK_c), .D(n2788));   // coms.v(192[10] 220[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5764 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[18]), .I2(data_in_field[26]), .I3(byte_transmit_counter2[1]), 
            .O(n6123));
    defparam byte_transmit_counter2_0__bdd_4_lut_5764.LUT_INIT = 16'he4aa;
    SB_LUT4 n6123_bdd_4_lut (.I0(n6123), .I1(data_in_field[10]), .I2(data_in_field[2]), 
            .I3(byte_transmit_counter2[1]), .O(n5752));
    defparam n6123_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i128 (.Q(data_in_field[127]), .C(CLK_c), .D(n2789));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i122 (.Q(data_in_field[121]), .C(CLK_c), .D(n2783));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i123 (.Q(data_in_field[122]), .C(CLK_c), .D(n2784));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i124 (.Q(data_in_field[123]), .C(CLK_c), .D(n2785));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i125 (.Q(data_in_field[124]), .C(CLK_c), .D(n2786));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i126 (.Q(data_in_field[125]), .C(CLK_c), .D(n2787));   // coms.v(192[10] 220[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n2526));   // coms.v(174[10] 182[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5754 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[50]), .I2(data_in_field[58]), .I3(byte_transmit_counter2[1]), 
            .O(n6117));
    defparam byte_transmit_counter2_0__bdd_4_lut_5754.LUT_INIT = 16'he4aa;
    SB_LUT4 i2480_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[8] [5]), .I3(data_in_field[69]), .O(n2731));
    defparam i2480_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_0___i4 (.Q(\data_out[10] [3]), .C(CLK_c), .D(n2839));   // coms.v(123[10] 164[6])
    SB_LUT4 n6117_bdd_4_lut (.I0(n6117), .I1(data_in_field[42]), .I2(data_in_field[34]), 
            .I3(byte_transmit_counter2[1]), .O(n5755));
    defparam n6117_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut (.I0(data_in_field[131]), .I1(n5381), .I2(n2012), 
            .I3(n5403), .O(n20));   // coms.v(202[14:57])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5749 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[82]), .I2(data_in_field[90]), .I3(byte_transmit_counter2[1]), 
            .O(n6111));
    defparam byte_transmit_counter2_0__bdd_4_lut_5749.LUT_INIT = 16'he4aa;
    SB_LUT4 n6111_bdd_4_lut (.I0(n6111), .I1(data_in_field[74]), .I2(data_in_field[66]), 
            .I3(byte_transmit_counter2[1]), .O(n5758));
    defparam n6111_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut (.I0(n1979), .I1(n2092), .I2(\data_in[19] [5]), .I3(n1892), 
            .O(n19));   // coms.v(202[14:57])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n5500), .I1(n18), .I2(n2149), .I3(n2065), 
            .O(n21_c));   // coms.v(202[14:57])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n2030), .I1(n20_adj_1870), .I2(n16), .I3(n5491), 
            .O(n5577));   // coms.v(82[17:399])
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(\data_in[18] [0]), .I1(n2095), .I2(n1908), .I3(n2021), 
            .O(n16_adj_1871));   // coms.v(202[14:57])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut (.I0(n15), .I1(tx_transmit_N_568[4]), .I2(n81_adj_1872), 
            .I3(n95), .O(n2872));
    defparam i1_4_lut.LUT_INIT = 16'hc0c4;
    SB_LUT4 i7_4_lut_adj_807 (.I0(data_in_field[7]), .I1(n5503), .I2(n5443), 
            .I3(n5524), .O(n17));   // coms.v(202[14:57])
    defparam i7_4_lut_adj_807.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i139 (.Q(data_in_field[138]), .C(CLK_c), .D(n2800));   // coms.v(192[10] 220[6])
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5744 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[114]), .I2(data_in_field[122]), .I3(byte_transmit_counter2[1]), 
            .O(n6105));
    defparam byte_transmit_counter2_0__bdd_4_lut_5744.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_2_lut (.I0(\data_in[18] [6]), .I1(data_in_field[138]), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_1873));   // coms.v(93[18:87])
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(CLK_c), .D(n2525));   // coms.v(174[10] 182[6])
    SB_LUT4 i2479_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[8] [4]), .I3(data_in_field[68]), .O(n2730));
    defparam i2479_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n6105_bdd_4_lut (.I0(n6105), .I1(data_in_field[106]), .I2(data_in_field[98]), 
            .I3(byte_transmit_counter2[1]), .O(n5761));
    defparam n6105_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut (.I0(n81_adj_1872), .I1(tx_transmit_N_568[5]), .I2(GND_net), 
            .I3(GND_net), .O(n2873));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_5759 (.I0(byte_transmit_counter2[2]), 
            .I1(n5758), .I2(n5761), .I3(byte_transmit_counter2[3]), .O(n6099));
    defparam byte_transmit_counter2_2__bdd_4_lut_5759.LUT_INIT = 16'he4aa;
    SB_LUT4 n6099_bdd_4_lut (.I0(n6099), .I1(n5755), .I2(n5752), .I3(byte_transmit_counter2[3]), 
            .O(n6102));
    defparam n6099_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5643_4_lut (.I0(tx_active), .I1(tx_transmit), .I2(n106), 
            .I3(n15), .O(n4813));
    defparam i5643_4_lut.LUT_INIT = 16'h0001;
    SB_DFF data_in_frame_0___i143 (.Q(data_in_field[142]), .C(CLK_c), .D(n2804));   // coms.v(192[10] 220[6])
    SB_LUT4 delay_counter_528_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n4763), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_528_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n4762), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(CLK_c), .D(n2524));   // coms.v(174[10] 182[6])
    SB_CARRY delay_counter_528_add_4_11 (.CI(n4762), .I0(GND_net), .I1(delay_counter[9]), 
            .CO(n4763));
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5739 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[17]), .I2(data_in_field[25]), .I3(byte_transmit_counter2[1]), 
            .O(n6093));
    defparam byte_transmit_counter2_0__bdd_4_lut_5739.LUT_INIT = 16'he4aa;
    SB_LUT4 i9_4_lut_adj_808 (.I0(data_in_field[125]), .I1(n1948), .I2(n5397), 
            .I3(n5512), .O(n22));   // coms.v(93[18:87])
    defparam i9_4_lut_adj_808.LUT_INIT = 16'h6996;
    SB_LUT4 i2478_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[8] [3]), .I3(data_in_field[67]), .O(n2729));
    defparam i2478_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut (.I0(data_in_field[113]), .I1(n2009), .I2(data_in_field[141]), 
            .I3(n5378), .O(n12));   // coms.v(202[14:57])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(CLK_c), .D(n2523));   // coms.v(174[10] 182[6])
    SB_LUT4 i2477_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[8] [2]), .I3(data_in_field[66]), .O(n2728));
    defparam i2477_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n2522));   // coms.v(174[10] 182[6])
    SB_DFF data_in_frame_0___i121 (.Q(data_in_field[120]), .C(CLK_c), .D(n2782));   // coms.v(192[10] 220[6])
    SB_LUT4 data_527_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(data[8]), 
            .I3(n4746), .O(n69[8])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n6093_bdd_4_lut (.I0(n6093), .I1(data_in_field[9]), .I2(data_in_field[1]), 
            .I3(byte_transmit_counter2[1]), .O(n5767));
    defparam n6093_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i115 (.Q(data_in_field[114]), .C(CLK_c), .D(n2776));   // coms.v(192[10] 220[6])
    SB_LUT4 i21_4_lut (.I0(n5593), .I1(n42), .I2(data_in_field[42]), .I3(data_in_field[19]), 
            .O(n48));   // coms.v(202[14:57])
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut (.I0(n43), .I1(n45), .I2(n44), .I3(n46), .O(n52));   // coms.v(202[14:57])
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i116 (.Q(data_in_field[115]), .C(CLK_c), .D(n2777));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i117 (.Q(data_in_field[116]), .C(CLK_c), .D(n2778));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i118 (.Q(data_in_field[117]), .C(CLK_c), .D(n2779));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i119 (.Q(data_in_field[118]), .C(CLK_c), .D(n2780));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i120 (.Q(data_in_field[119]), .C(CLK_c), .D(n2781));   // coms.v(192[10] 220[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(CLK_c), .D(n2521));   // coms.v(174[10] 182[6])
    SB_LUT4 delay_counter_528_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n4761), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_809 (.I0(tx_active), .I1(tx_active_prev), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_1875));   // verilog/TinyFPGA_B.v(77[8] 84[4])
    defparam i1_2_lut_adj_809.LUT_INIT = 16'h4444;
    SB_LUT4 i5572_4_lut (.I0(\data_out[10] [3]), .I1(byte_transmit_counter[1]), 
            .I2(\data_out[11] [3]), .I3(byte_transmit_counter[0]), .O(n5853));
    defparam i5572_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY data_527_add_4_10 (.CI(n4746), .I0(GND_net), .I1(data[8]), 
            .CO(n4747));
    SB_LUT4 i20_4_lut (.I0(n5551), .I1(n5557), .I2(n5554), .I3(n5581), 
            .O(n47));   // coms.v(202[14:57])
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_810 (.I0(n5488), .I1(n12), .I2(n1886), .I3(\data_in[18] [1]), 
            .O(n5489));   // coms.v(202[14:57])
    defparam i6_4_lut_adj_810.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(data_in_field[10]), .I1(data_in_field[51]), .I2(data_in_field[9]), 
            .I3(GND_net), .O(n22_adj_1876));   // coms.v(202[14:57])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5729 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[49]), .I2(data_in_field[57]), .I3(byte_transmit_counter2[1]), 
            .O(n6087));
    defparam byte_transmit_counter2_0__bdd_4_lut_5729.LUT_INIT = 16'he4aa;
    SB_LUT4 n6087_bdd_4_lut (.I0(n6087), .I1(data_in_field[41]), .I2(data_in_field[33]), 
            .I3(byte_transmit_counter2[1]), .O(n5770));
    defparam n6087_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10_4_lut_adj_811 (.I0(\data_in[18] [3]), .I1(data_in_field[130]), 
            .I2(n1955), .I3(data_in_field[70]), .O(n27));   // coms.v(202[14:57])
    defparam i10_4_lut_adj_811.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5724 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_in_frame[18] [7]), .I2(\data_in_frame[19] [7]), .I3(byte_transmit_counter2[1]), 
            .O(n6081));
    defparam byte_transmit_counter2_0__bdd_4_lut_5724.LUT_INIT = 16'he4aa;
    SB_LUT4 n6081_bdd_4_lut (.I0(n6081), .I1(data_in_field[143]), .I2(data_in_field[135]), 
            .I3(byte_transmit_counter2[1]), .O(n6084));
    defparam n6081_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY delay_counter_528_add_4_10 (.CI(n4761), .I0(GND_net), .I1(delay_counter[8]), 
            .CO(n4762));
    SB_LUT4 data_527_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(data[7]), 
            .I3(n4745), .O(n69[7])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5719 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[81]), .I2(data_in_field[89]), .I3(byte_transmit_counter2[1]), 
            .O(n6075));
    defparam byte_transmit_counter2_0__bdd_4_lut_5719.LUT_INIT = 16'he4aa;
    SB_LUT4 i11_4_lut (.I0(data_in_field[86]), .I1(n22), .I2(n16_adj_1873), 
            .I3(data_in_field[73]), .O(n24));   // coms.v(93[18:87])
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i114 (.Q(data_in_field[113]), .C(CLK_c), .D(n2775));   // coms.v(192[10] 220[6])
    SB_LUT4 n6075_bdd_4_lut (.I0(n6075), .I1(data_in_field[73]), .I2(data_in_field[65]), 
            .I3(byte_transmit_counter2[1]), .O(n5773));
    defparam n6075_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 delay_counter_528_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(delay_counter[7]), 
            .I3(n4760), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut (.I0(n5375), .I1(n30), .I2(n24_adj_1877), .I3(n5381), 
            .O(n32));   // coms.v(202[14:57])
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5714 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_in_frame[18] [0]), .I2(\data_in_frame[19] [0]), .I3(byte_transmit_counter2[1]), 
            .O(n6069));
    defparam byte_transmit_counter2_0__bdd_4_lut_5714.LUT_INIT = 16'he4aa;
    SB_LUT4 n6069_bdd_4_lut (.I0(n6069), .I1(data_in_field[136]), .I2(data_in_field[128]), 
            .I3(byte_transmit_counter2[1]), .O(n6072));
    defparam n6069_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i12_4_lut (.I0(n5536), .I1(n24), .I2(n20_adj_1878), .I3(n5572), 
            .O(n5586));   // coms.v(93[18:87])
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_812 (.I0(n5489), .I1(n47), .I2(n52), .I3(n48), 
            .O(n24_adj_1879));   // coms.v(202[14:57])
    defparam i8_4_lut_adj_812.LUT_INIT = 16'hebbe;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5709 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[113]), .I2(data_in_field[121]), .I3(byte_transmit_counter2[1]), 
            .O(n6063));
    defparam byte_transmit_counter2_0__bdd_4_lut_5709.LUT_INIT = 16'he4aa;
    SB_LUT4 n6063_bdd_4_lut (.I0(n6063), .I1(data_in_field[105]), .I2(data_in_field[97]), 
            .I3(byte_transmit_counter2[1]), .O(n5776));
    defparam n6063_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_0___i159 (.Q(\data_in[19] [6]), .C(CLK_c), .D(n2660));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i160 (.Q(\data_in[19] [7]), .C(CLK_c), .D(n2661));   // coms.v(174[10] 182[6])
    SB_DFF data_in_frame_0___i2 (.Q(data_in_field[1]), .C(CLK_c), .D(n2662));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i3 (.Q(data_in_field[2]), .C(CLK_c), .D(n2664));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i4 (.Q(data_in_field[3]), .C(CLK_c), .D(n2665));   // coms.v(192[10] 220[6])
    SB_DFF data_in_0___i158 (.Q(\data_in[19] [5]), .C(CLK_c), .D(n2659));   // coms.v(174[10] 182[6])
    SB_CARRY delay_counter_528_add_4_9 (.CI(n4760), .I0(GND_net), .I1(delay_counter[7]), 
            .CO(n4761));
    SB_LUT4 i2476_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[8] [1]), .I3(data_in_field[65]), .O(n2727));
    defparam i2476_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY data_527_add_4_9 (.CI(n4745), .I0(GND_net), .I1(data[7]), 
            .CO(n4746));
    SB_LUT4 i1_2_lut_adj_813 (.I0(\data_out[11] [1]), .I1(\data_out[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // coms.v(85[17:241])
    defparam i1_2_lut_adj_813.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut (.I0(n27), .I1(data_in_field[135]), .I2(n22_adj_1876), 
            .I3(data_in_field[38]), .O(n31));   // coms.v(202[14:57])
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i121 (.Q(\data_in[15] [0]), .C(CLK_c), .D(n2622));   // coms.v(174[10] 182[6])
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_5734 (.I0(byte_transmit_counter2[2]), 
            .I1(n5773), .I2(n5776), .I3(byte_transmit_counter2[3]), .O(n6057));
    defparam byte_transmit_counter2_2__bdd_4_lut_5734.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut (.I0(\data_in[19] [2]), .I1(data_in_field[120]), .I2(n1866), 
            .I3(n1814), .O(n10));   // coms.v(202[14:57])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i122 (.Q(\data_in[15] [1]), .C(CLK_c), .D(n2623));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i123 (.Q(\data_in[15] [2]), .C(CLK_c), .D(n2624));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i124 (.Q(\data_in[15] [3]), .C(CLK_c), .D(n2625));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i125 (.Q(\data_in[15] [4]), .C(CLK_c), .D(n2626));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i126 (.Q(\data_in[15] [5]), .C(CLK_c), .D(n2627));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i120 (.Q(\data_in[14] [7]), .C(CLK_c), .D(n2621));   // coms.v(174[10] 182[6])
    SB_LUT4 n6057_bdd_4_lut (.I0(n6057), .I1(n5770), .I2(n5767), .I3(byte_transmit_counter2[3]), 
            .O(n6060));
    defparam n6057_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_0___i87 (.Q(\data_in[10] [6]), .C(CLK_c), .D(n2588));   // coms.v(174[10] 182[6])
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_0_i31_4_lut (.I0(n6018), .I1(n6072), 
            .I2(byte_transmit_counter2[4]), .I3(n1081), .O(tx2_data[0]));   // coms.v(189[35:57])
    defparam byte_transmit_counter2_4__I_0_Mux_0_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n2520));   // coms.v(174[10] 182[6])
    SB_LUT4 i2475_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[8] [0]), .I3(data_in_field[64]), .O(n2726));
    defparam i2475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_814 (.I0(n81_adj_1872), .I1(tx_transmit_N_568[6]), 
            .I2(GND_net), .I3(GND_net), .O(n2874));
    defparam i1_2_lut_adj_814.LUT_INIT = 16'h8888;
    SB_LUT4 data_527_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(data[6]), 
            .I3(n4744), .O(n69[6])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_in_0___i48 (.Q(\data_in[5] [7]), .C(CLK_c), .D(n2549));   // coms.v(174[10] 182[6])
    SB_LUT4 i2474_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[7] [7]), .I3(data_in_field[63]), .O(n2725));
    defparam i2474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2473_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[7] [6]), .I3(data_in_field[62]), .O(n2724));
    defparam i2473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i49 (.Q(\data_in[6] [0]), .C(CLK_c), .D(n2550));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i50 (.Q(\data_in[6] [1]), .C(CLK_c), .D(n2551));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i51 (.Q(\data_in[6] [2]), .C(CLK_c), .D(n2552));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i52 (.Q(\data_in[6] [3]), .C(CLK_c), .D(n2553));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i53 (.Q(\data_in[6] [4]), .C(CLK_c), .D(n2554));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i47 (.Q(\data_in[5] [6]), .C(CLK_c), .D(n2548));   // coms.v(174[10] 182[6])
    SB_LUT4 i2472_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[7] [5]), .I3(data_in_field[61]), .O(n2723));
    defparam i2472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(CLK_c), .D(n2519));   // coms.v(174[10] 182[6])
    SB_CARRY data_527_add_4_8 (.CI(n4744), .I0(GND_net), .I1(data[6]), 
            .CO(n4745));
    SB_LUT4 i3_2_lut_adj_815 (.I0(data_in_field[99]), .I1(data_in_field[64]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_1880));   // coms.v(89[18:383])
    defparam i3_2_lut_adj_815.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_816 (.I0(n2039), .I1(data_in_field[9]), .I2(data_in_field[121]), 
            .I3(n5412), .O(n22_adj_1881));   // coms.v(89[18:383])
    defparam i9_4_lut_adj_816.LUT_INIT = 16'h6996;
    SB_LUT4 i2471_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[7] [4]), .I3(data_in_field[60]), .O(n2722));
    defparam i2471_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 delay_counter_528_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(delay_counter[6]), 
            .I3(n4759), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_3_lut (.I0(n5569), .I1(data_in_field[114]), .I2(\data_in[18] [2]), 
            .I3(GND_net), .O(n20_adj_1882));   // coms.v(89[18:383])
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut (.I0(tx_active), .I1(tx_transmit), .I2(n21), 
            .I3(GND_net), .O(n81_adj_1872));   // coms.v(19[7:18])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(CLK_c), .D(n2518));   // coms.v(174[10] 182[6])
    SB_LUT4 i1_2_lut_adj_817 (.I0(n81_adj_1872), .I1(tx_transmit_N_568[7]), 
            .I2(GND_net), .I3(GND_net), .O(n2875));
    defparam i1_2_lut_adj_817.LUT_INIT = 16'h8888;
    SB_LUT4 i2470_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[7] [3]), .I3(data_in_field[59]), .O(n2721));
    defparam i2470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2469_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[7] [2]), .I3(data_in_field[58]), .O(n2720));
    defparam i2469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_818 (.I0(n2107), .I1(n22_adj_1881), .I2(n16_adj_1880), 
            .I3(data_in_field[50]), .O(n24_adj_1884));   // coms.v(89[18:383])
    defparam i11_4_lut_adj_818.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_819 (.I0(n5384), .I1(n5476), .I2(n5427), .I3(n5521), 
            .O(n24_adj_1885));   // coms.v(86[17:391])
    defparam i10_4_lut_adj_819.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_820 (.I0(data_in_field[118]), .I1(data_in_field[51]), 
            .I2(n2152), .I3(data_in_field[126]), .O(n23));   // coms.v(86[17:391])
    defparam i9_4_lut_adj_820.LUT_INIT = 16'h6996;
    SB_DFF data_out_0___i3 (.Q(\data_out[10] [2]), .C(CLK_c), .D(n2838));   // coms.v(123[10] 164[6])
    SB_LUT4 i2468_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[7] [1]), .I3(data_in_field[57]), .O(n2719));
    defparam i2468_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_821 (.I0(n5545), .I1(n22_adj_1886), .I2(data_in_field[117]), 
            .I3(n1855), .O(n25));   // coms.v(86[17:391])
    defparam i11_4_lut_adj_821.LUT_INIT = 16'h6996;
    SB_DFF data_out_0___i13 (.Q(\data_out[11] [4]), .C(CLK_c), .D(n2848));   // coms.v(123[10] 164[6])
    SB_LUT4 i5_4_lut_adj_822 (.I0(n5466), .I1(n10), .I2(data_in_field[57]), 
            .I3(data_in_field[113]), .O(n5519));   // coms.v(202[14:57])
    defparam i5_4_lut_adj_822.LUT_INIT = 16'h6996;
    SB_CARRY delay_counter_528_add_4_8 (.CI(n4759), .I0(GND_net), .I1(delay_counter[6]), 
            .CO(n4760));
    SB_LUT4 data_527_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(data[5]), 
            .I3(n4743), .O(n69[5])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2467_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[7] [0]), .I3(data_in_field[56]), .O(n2718));
    defparam i2467_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i131 (.Q(data_in_field[130]), .C(CLK_c), .D(n2792));   // coms.v(192[10] 220[6])
    SB_LUT4 i2466_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[6] [7]), .I3(data_in_field[55]), .O(n2717));
    defparam i2466_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2465_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[6] [6]), .I3(data_in_field[54]), .O(n2716));
    defparam i2465_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2464_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[6] [5]), .I3(data_in_field[53]), .O(n2715));
    defparam i2464_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_823 (.I0(n3703), .I1(\FRAME_MATCHER.wait_for_transmission_N_909 ), 
            .I2(\FRAME_MATCHER.wait_for_transmission ), .I3(n3689), .O(n6));   // coms.v(192[10] 220[6])
    defparam i14_4_lut_adj_823.LUT_INIT = 16'hf5c5;
    SB_LUT4 i9_4_lut_adj_824 (.I0(n5560), .I1(n18_adj_1887), .I2(data_in_field[101]), 
            .I3(\data_in[18] [4]), .O(n20_adj_1888));   // coms.v(202[14:57])
    defparam i9_4_lut_adj_824.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(CLK_c), 
           .D(n2811));   // coms.v(192[10] 220[6])
    SB_LUT4 i8_4_lut_adj_825 (.I0(n1926), .I1(n5494), .I2(n5394), .I3(n5527), 
            .O(n19_adj_1889));   // coms.v(202[14:57])
    defparam i8_4_lut_adj_825.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_826 (.I0(n5519), .I1(n25), .I2(n23), .I3(n24_adj_1885), 
            .O(n22_adj_1890));   // coms.v(202[14:57])
    defparam i6_4_lut_adj_826.LUT_INIT = 16'hbeeb;
    SB_DFF data_out_0___i12 (.Q(\data_out[11] [3]), .C(CLK_c), .D(n2847));   // coms.v(123[10] 164[6])
    SB_DFF data_in_frame_0___i135 (.Q(data_in_field[134]), .C(CLK_c), .D(n2796));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(CLK_c), 
           .D(n2810));   // coms.v(192[10] 220[6])
    SB_LUT4 i2463_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[6] [4]), .I3(data_in_field[52]), .O(n2714));
    defparam i2463_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i9_3_lut (.I0(\data_out[10] [0]), 
            .I1(\data_out[11] [0]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n9));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5588_4_lut (.I0(\data_out[18] [0]), .I1(n1508), .I2(\data_out[19] [0]), 
            .I3(byte_transmit_counter[0]), .O(n5810));   // coms.v(39[29:50])
    defparam i5588_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i957_4_lut (.I0(byte_transmit_counter[0]), .I1(n9), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[1]), .O(n1198));   // coms.v(39[29:50])
    defparam i957_4_lut.LUT_INIT = 16'hc50a;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_4_lut (.I0(n1198), .I1(n5810), 
            .I2(byte_transmit_counter[4]), .I3(byte_transmit_counter[2]), 
            .O(tx_data[0]));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i9_3_lut (.I0(\data_out[10] [1]), 
            .I1(\data_out[11] [1]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n9_adj_1891));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_1_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5595_4_lut (.I0(\data_out[18] [1]), .I1(byte_transmit_counter[1]), 
            .I2(\data_out[19] [1]), .I3(byte_transmit_counter[0]), .O(n5845));   // coms.v(39[29:50])
    defparam i5595_4_lut.LUT_INIT = 16'hf3bb;
    SB_LUT4 i12_4_lut_adj_827 (.I0(n5503), .I1(n24_adj_1884), .I2(n20_adj_1882), 
            .I3(n5536), .O(n5570));   // coms.v(89[18:383])
    defparam i12_4_lut_adj_827.LUT_INIT = 16'h6996;
    SB_LUT4 add_1824_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n4709), .O(tx_transmit_N_568[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1824_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut_adj_828 (.I0(data_in_field[12]), .I1(data_in_field[55]), 
            .I2(n2077), .I3(\data_in[19] [0]), .O(n40));   // coms.v(202[14:57])
    defparam i14_4_lut_adj_828.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n5521), .I1(n5539), .I2(n5527), .I3(n5548), 
            .O(n45_adj_1892));   // coms.v(202[14:57])
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_DFF byte_transmit_counter__i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
           .D(n2874));   // coms.v(123[10] 164[6])
    SB_DFF byte_transmit_counter__i3 (.Q(byte_transmit_counter[3]), .C(CLK_c), 
           .D(n2871));   // coms.v(123[10] 164[6])
    SB_DFF data_out_0___i14 (.Q(\data_out[11] [5]), .C(CLK_c), .D(n2849));   // coms.v(123[10] 164[6])
    SB_DFF byte_transmit_counter__i2 (.Q(byte_transmit_counter[2]), .C(CLK_c), 
           .D(n2870));   // coms.v(123[10] 164[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i15_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(n9_adj_1891), .I2(byte_transmit_counter[3]), .I3(byte_transmit_counter[1]), 
            .O(n15_adj_1893));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_1_i15_4_lut.LUT_INIT = 16'h4aa5;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_4_lut (.I0(n15_adj_1893), 
            .I1(n5845), .I2(byte_transmit_counter[4]), .I3(n1251), .O(i_Tx_Byte[1]));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF data_out_0___i2 (.Q(\data_out[10] [1]), .C(CLK_c), .D(n2835));   // coms.v(123[10] 164[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(CLK_c), 
           .D(n2807));   // coms.v(192[10] 220[6])
    SB_DFF byte_transmit_counter__i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
           .D(n2873));   // coms.v(123[10] 164[6])
    SB_DFF byte_transmit_counter__i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
           .D(n2869));   // coms.v(123[10] 164[6])
    SB_LUT4 i22_4_lut (.I0(n5388), .I1(n44_adj_1894), .I2(n34), .I3(n5397), 
            .O(n48_adj_1895));   // coms.v(202[14:57])
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_DFF byte_transmit_counter__i4 (.Q(byte_transmit_counter[4]), .C(CLK_c), 
           .D(n2872));   // coms.v(123[10] 164[6])
    SB_DFF data_out_0___i10 (.Q(\data_out[11] [1]), .C(CLK_c), .D(n2845));   // coms.v(123[10] 164[6])
    SB_LUT4 i2462_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[6] [3]), .I3(data_in_field[51]), .O(n2713));
    defparam i2462_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21_4_lut_adj_829 (.I0(n41), .I1(n31_adj_1896), .I2(data_in_field[61]), 
            .I3(data_in_field[20]), .O(n47_adj_1897));   // coms.v(202[14:57])
    defparam i21_4_lut_adj_829.LUT_INIT = 16'h6996;
    SB_LUT4 i5587_4_lut (.I0(\data_out[18] [2]), .I1(n1508), .I2(\data_out[19] [2]), 
            .I3(byte_transmit_counter[0]), .O(n5840));   // coms.v(39[29:50])
    defparam i5587_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_out_0___i30 (.Q(\data_out[19] [5]), .C(CLK_c), .D(n2865));   // coms.v(123[10] 164[6])
    SB_LUT4 i2044_4_lut (.I0(byte_transmit_counter[0]), .I1(\data_out[10] [2]), 
            .I2(byte_transmit_counter[3]), .I3(\data_out[11] [2]), .O(n2293));   // coms.v(39[29:50])
    defparam i2044_4_lut.LUT_INIT = 16'he545;
    SB_LUT4 i7_4_lut_adj_830 (.I0(n13), .I1(n5497), .I2(n12_adj_1898), 
            .I3(n5500), .O(n5567));   // coms.v(202[14:57])
    defparam i7_4_lut_adj_830.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_4_lut (.I0(n2293), .I1(n5840), 
            .I2(byte_transmit_counter[4]), .I3(n1253), .O(i_Tx_Byte[2]));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_4_lut.LUT_INIT = 16'hcac0;
    SB_DFF data_out_0___i27 (.Q(\data_out[19] [2]), .C(CLK_c), .D(n2862));   // coms.v(123[10] 164[6])
    SB_LUT4 i5582_4_lut (.I0(\data_out[18] [3]), .I1(byte_transmit_counter[1]), 
            .I2(\data_out[19] [3]), .I3(byte_transmit_counter[0]), .O(n5837));   // coms.v(39[29:50])
    defparam i5582_4_lut.LUT_INIT = 16'hf3bb;
    SB_DFF data_out_0___i29 (.Q(\data_out[19] [4]), .C(CLK_c), .D(n2864));   // coms.v(123[10] 164[6])
    SB_DFF data_out_0___i26 (.Q(\data_out[19] [1]), .C(CLK_c), .D(n2861));   // coms.v(123[10] 164[6])
    SB_LUT4 i23_4_lut (.I0(n45_adj_1892), .I1(n5563), .I2(n40), .I3(n5590), 
            .O(n49));   // coms.v(202[14:57])
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_831 (.I0(n5430), .I1(n5539), .I2(n5506), .I3(n5575), 
            .O(n14));   // coms.v(83[17:391])
    defparam i6_4_lut_adj_831.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_832 (.I0(\data_in[19] [4]), .I1(n1855), .I2(data_in_field[115]), 
            .I3(n1917), .O(n13_adj_1899));   // coms.v(83[17:391])
    defparam i5_4_lut_adj_832.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(CLK_c), 
           .D(n2806));   // coms.v(192[10] 220[6])
    SB_LUT4 i2461_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[6] [2]), .I3(data_in_field[50]), .O(n2712));
    defparam i2461_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_0___i32 (.Q(\data_out[19] [7]), .C(CLK_c), .D(n2867));   // coms.v(123[10] 164[6])
    SB_DFF data_out_0___i28 (.Q(\data_out[19] [3]), .C(CLK_c), .D(n2863));   // coms.v(123[10] 164[6])
    SB_LUT4 i19_4_lut_adj_833 (.I0(n37), .I1(n35), .I2(n31_adj_1900), 
            .I3(n32_adj_1901), .O(n5582));   // coms.v(82[17:399])
    defparam i19_4_lut_adj_833.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_4_lut (.I0(n6312), .I1(n5837), 
            .I2(byte_transmit_counter[4]), .I3(n1251), .O(i_Tx_Byte[3]));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_834 (.I0(n49), .I1(n5567), .I2(n47_adj_1897), 
            .I3(n48_adj_1895), .O(n17_adj_1902));   // coms.v(202[14:57])
    defparam i1_4_lut_adj_834.LUT_INIT = 16'hb77b;
    SB_DFF data_527__i0 (.Q(data[0]), .C(CLK_c), .D(n69[0]));   // coms.v(126[13:19])
    SB_LUT4 i11_4_lut_adj_835 (.I0(n5512), .I1(n22_adj_1903), .I2(n18_adj_1904), 
            .I3(n5542), .O(n5589));   // coms.v(92[18:361])
    defparam i11_4_lut_adj_835.LUT_INIT = 16'h6996;
    SB_LUT4 i2460_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[6] [1]), .I3(data_in_field[49]), .O(n2711));
    defparam i2460_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2459_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[6] [0]), .I3(data_in_field[48]), .O(n2710));
    defparam i2459_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i1 (.Q(data_in_field[0]), .C(CLK_c), .D(n2385));   // coms.v(192[10] 220[6])
    SB_LUT4 i4_4_lut_adj_836 (.I0(n5577), .I1(n21_c), .I2(n19), .I3(n20), 
            .O(n20_adj_1905));   // coms.v(202[14:57])
    defparam i4_4_lut_adj_836.LUT_INIT = 16'hd77d;
    SB_DFF delay_counter_528__i0 (.Q(delay_counter[0]), .C(CLK_c), .D(n1[0]));   // coms.v(159[11] 161[5])
    SB_LUT4 i9_4_lut_adj_837 (.I0(n17), .I1(n5557), .I2(n16_adj_1871), 
            .I3(n5572), .O(n5574));   // coms.v(202[14:57])
    defparam i9_4_lut_adj_837.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i9_3_lut (.I0(\data_out[10] [4]), 
            .I1(\data_out[11] [4]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n9_adj_1906));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_4_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut_adj_838 (.I0(n17_adj_1902), .I1(n5582), .I2(n13_adj_1899), 
            .I3(n14), .O(n25_adj_1907));   // coms.v(202[14:57])
    defparam i9_4_lut_adj_838.LUT_INIT = 16'hfeef;
    SB_LUT4 i2458_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[5] [7]), .I3(data_in_field[47]), .O(n2709));
    defparam i2458_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_0___i24 (.Q(\data_out[18] [7]), .C(CLK_c), .D(n2859));   // coms.v(123[10] 164[6])
    SB_DFF data_out_0___i23 (.Q(\data_out[18] [6]), .C(CLK_c), .D(n2858));   // coms.v(123[10] 164[6])
    SB_DFF data_in_frame_0___i142 (.Q(data_in_field[141]), .C(CLK_c), .D(n2803));   // coms.v(192[10] 220[6])
    SB_LUT4 i2457_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[5] [6]), .I3(data_in_field[46]), .O(n2708));
    defparam i2457_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out[18] [4]), 
            .I1(\data_out[19] [4]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n17_adj_1908));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_839 (.I0(n31), .I1(n24_adj_1879), .I2(n5586), 
            .I3(n32), .O(n28));   // coms.v(202[14:57])
    defparam i12_4_lut_adj_839.LUT_INIT = 16'hfdfe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i15_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n9_adj_1906), .I2(byte_transmit_counter[3]), .I3(byte_transmit_counter[2]), 
            .O(n15_adj_1909));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_4_i15_4_lut.LUT_INIT = 16'ha5d5;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i31_4_lut (.I0(n15_adj_1909), 
            .I1(n17_adj_1908), .I2(byte_transmit_counter[4]), .I3(n1508), 
            .O(i_Tx_Byte[4]));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_4_i31_4_lut.LUT_INIT = 16'hca0a;
    SB_DFF data_in_frame_0___i141 (.Q(data_in_field[140]), .C(CLK_c), .D(n2802));   // coms.v(192[10] 220[6])
    SB_LUT4 i11_4_lut_adj_840 (.I0(n5570), .I1(n22_adj_1890), .I2(n19_adj_1889), 
            .I3(n20_adj_1888), .O(n27_adj_1910));   // coms.v(202[14:57])
    defparam i11_4_lut_adj_840.LUT_INIT = 16'hdffd;
    SB_LUT4 i13_4_lut (.I0(n25_adj_1907), .I1(n5574), .I2(n20_adj_1905), 
            .I3(n5589), .O(n29));   // coms.v(202[14:57])
    defparam i13_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_1824_3 (.CI(n4703), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n4704));
    SB_LUT4 i2456_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[5] [5]), .I3(data_in_field[45]), .O(n2707));
    defparam i2456_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3459_4_lut (.I0(n29), .I1(n1729), .I2(n27_adj_1910), .I3(n28), 
            .O(n3703));
    defparam i3459_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5640_3_lut_4_lut (.I0(tx_active), .I1(tx_transmit), .I2(n15), 
            .I3(n106), .O(n4333));   // coms.v(19[7:18])
    defparam i5640_3_lut_4_lut.LUT_INIT = 16'h1110;
    SB_LUT4 i2455_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[5] [4]), .I3(data_in_field[44]), .O(n2706));
    defparam i2455_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i138 (.Q(data_in_field[137]), .C(CLK_c), .D(n2799));   // coms.v(192[10] 220[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i9_3_lut (.I0(\data_out[10] [5]), 
            .I1(\data_out[11] [5]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n9_adj_1911));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_5_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5571_4_lut (.I0(\data_out[18] [5]), .I1(n1508), .I2(\data_out[19] [5]), 
            .I3(byte_transmit_counter[0]), .O(n5833));   // coms.v(39[29:50])
    defparam i5571_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i137 (.Q(data_in_field[136]), .C(CLK_c), .D(n2798));   // coms.v(192[10] 220[6])
    SB_LUT4 i748_4_lut (.I0(byte_transmit_counter[0]), .I1(n9_adj_1911), 
            .I2(byte_transmit_counter[3]), .I3(byte_transmit_counter[1]), 
            .O(n989));   // coms.v(39[29:50])
    defparam i748_4_lut.LUT_INIT = 16'hc50a;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_4_lut (.I0(n989), .I1(n5833), 
            .I2(byte_transmit_counter[4]), .I3(byte_transmit_counter[2]), 
            .O(i_Tx_Byte[5]));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_4_lut.LUT_INIT = 16'hc0ca;
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(CLK_c), 
           .D(n2808));   // coms.v(192[10] 220[6])
    SB_LUT4 i2454_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[5] [3]), .I3(data_in_field[43]), .O(n2705));
    defparam i2454_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i35_3_lut (.I0(\data_out[10] [6]), .I1(\data_out[11] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n31_adj_1912));   // coms.v(39[29:50])
    defparam i35_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out[18] [6]), 
            .I1(\data_out[19] [6]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n17_adj_1913));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_841 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter[0]), .I3(n31_adj_1912), .O(n22_adj_1914));   // coms.v(39[29:50])
    defparam i1_4_lut_adj_841.LUT_INIT = 16'h54dc;
    SB_LUT4 i5575_3_lut (.I0(n17_adj_1913), .I1(n1251), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n5830));   // coms.v(39[29:50])
    defparam i5575_3_lut.LUT_INIT = 16'h2323;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(n5830), .I2(byte_transmit_counter[4]), .I3(n22_adj_1914), 
            .O(i_Tx_Byte[6]));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_4_lut.LUT_INIT = 16'hcacf;
    SB_LUT4 i2453_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[5] [2]), .I3(data_in_field[42]), .O(n2704));
    defparam i2453_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_0___i9 (.Q(\data_out[11] [0]), .C(CLK_c), .D(n2844));   // coms.v(123[10] 164[6])
    SB_DFF data_out_0___i25 (.Q(\data_out[19] [0]), .C(CLK_c), .D(n2860));   // coms.v(123[10] 164[6])
    SB_DFF data_out_0___i8 (.Q(\data_out[10] [7]), .C(CLK_c), .D(n2843));   // coms.v(123[10] 164[6])
    SB_LUT4 i2452_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[5] [1]), .I3(data_in_field[41]), .O(n2703));
    defparam i2452_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2451_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[5] [0]), .I3(data_in_field[40]), .O(n2702));
    defparam i2451_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(CLK_c), 
           .D(n2812));   // coms.v(192[10] 220[6])
    SB_CARRY data_527_add_4_7 (.CI(n4743), .I0(GND_net), .I1(data[5]), 
            .CO(n4744));
    SB_DFF data_out_0___i22 (.Q(\data_out[18] [5]), .C(CLK_c), .D(n2857));   // coms.v(123[10] 164[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(CLK_c), .D(n2517));   // coms.v(174[10] 182[6])
    SB_LUT4 i2450_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[4] [7]), .I3(data_in_field[39]), .O(n2701));
    defparam i2450_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_0___i15 (.Q(\data_out[11] [6]), .C(CLK_c), .D(n2850));   // coms.v(123[10] 164[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(CLK_c), .D(n2516));   // coms.v(174[10] 182[6])
    SB_DFF data_out_0___i7 (.Q(\data_out[10] [6]), .C(CLK_c), .D(n2842));   // coms.v(123[10] 164[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(CLK_c), .D(n2515));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(CLK_c), .D(n2514));   // coms.v(174[10] 182[6])
    SB_LUT4 i2449_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[4] [6]), .I3(data_in_field[38]), .O(n2700));
    defparam i2449_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(CLK_c), .D(n2513));   // coms.v(174[10] 182[6])
    SB_DFF delay_counter_528__i5 (.Q(delay_counter[5]), .C(CLK_c), .D(n1[5]));   // coms.v(159[11] 161[5])
    SB_LUT4 i2448_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[4] [5]), .I3(data_in_field[37]), .O(n2699));
    defparam i2448_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF tx2_transmit_1801 (.Q(r_SM_Main_2__N_1770[0]), .C(CLK_c), .D(tx2_transmit_N_915));   // coms.v(192[10] 220[6])
    SB_LUT4 delay_counter_528_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(delay_counter[5]), 
            .I3(n4758), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(CLK_c), 
           .D(n2819));   // coms.v(192[10] 220[6])
    SB_CARRY delay_counter_528_add_4_7 (.CI(n4758), .I0(GND_net), .I1(delay_counter[5]), 
            .CO(n4759));
    SB_DFF tx_active_prev_1793 (.Q(tx_active_prev), .C(CLK_c), .D(tx_active));   // coms.v(123[10] 164[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n2512));   // coms.v(174[10] 182[6])
    SB_LUT4 i2447_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[4] [4]), .I3(data_in_field[36]), .O(n2698));
    defparam i2447_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2446_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[4] [3]), .I3(data_in_field[35]), .O(n2697));
    defparam i2446_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2445_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[4] [2]), .I3(data_in_field[34]), .O(n2696));
    defparam i2445_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2444_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[4] [1]), .I3(data_in_field[33]), .O(n2695));
    defparam i2444_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 tx2_transmit_I_0_1818_4_lut (.I0(n3703), .I1(\FRAME_MATCHER.wait_for_transmission_N_909 ), 
            .I2(\FRAME_MATCHER.wait_for_transmission ), .I3(n3689), .O(tx2_transmit_N_915));   // coms.v(209[14] 219[8])
    defparam tx2_transmit_I_0_1818_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 i2443_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[4] [0]), .I3(data_in_field[32]), .O(n2694));
    defparam i2443_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2442_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[3] [7]), .I3(data_in_field[31]), .O(n2693));
    defparam i2442_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2441_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[3] [6]), .I3(data_in_field[30]), .O(n2692));
    defparam i2441_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_842 (.I0(tx_transmit_N_568[3]), .I1(tx_transmit_N_568[2]), 
            .I2(GND_net), .I3(GND_net), .O(n95));
    defparam i1_2_lut_adj_842.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(tx_transmit_N_568[5]), .I1(tx_transmit_N_568[7]), 
            .I2(tx_transmit_N_568[6]), .I3(GND_net), .O(n15));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2440_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[3] [5]), .I3(data_in_field[29]), .O(n2691));
    defparam i2440_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_843 (.I0(n2134), .I1(n2092), .I2(data_in_field[6]), 
            .I3(data_in_field[75]), .O(n10_adj_1915));   // coms.v(86[17:391])
    defparam i4_4_lut_adj_843.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_844 (.I0(\data_out[11] [7]), .I1(\data_out[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));
    defparam i1_2_lut_adj_844.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_845 (.I0(data_in_field[118]), .I1(data_in_field[140]), 
            .I2(GND_net), .I3(GND_net), .O(n5572));   // coms.v(93[18:87])
    defparam i1_2_lut_adj_845.LUT_INIT = 16'h6666;
    SB_LUT4 i120_2_lut (.I0(tx_transmit_N_568[4]), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n106));   // coms.v(19[7:18])
    defparam i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_846 (.I0(data_in_field[84]), .I1(data_in_field[54]), 
            .I2(GND_net), .I3(GND_net), .O(n5536));   // coms.v(89[18:383])
    defparam i1_2_lut_adj_846.LUT_INIT = 16'h6666;
    SB_LUT4 i2439_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[3] [4]), .I3(data_in_field[28]), .O(n2690));
    defparam i2439_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_847 (.I0(data_in_field[133]), .I1(data_in_field[103]), 
            .I2(GND_net), .I3(GND_net), .O(n2152));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_847.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_848 (.I0(n2068), .I1(data_in_field[99]), .I2(data_in_field[68]), 
            .I3(n6_adj_1917), .O(n5512));   // coms.v(93[18:87])
    defparam i4_4_lut_adj_848.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_849 (.I0(n2152), .I1(data_in_field[132]), .I2(data_in_field[43]), 
            .I3(n6_adj_1918), .O(n5397));   // coms.v(93[18:87])
    defparam i4_4_lut_adj_849.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(data_in_field[134]), .I1(n2000), .I2(data_in_field[142]), 
            .I3(n2053), .O(n5503));   // coms.v(89[18:383])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_850 (.I0(data_in_field[67]), .I1(data_in_field[119]), 
            .I2(data_in_field[35]), .I3(GND_net), .O(n2095));   // coms.v(202[14:57])
    defparam i2_3_lut_adj_850.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(n5400), .I1(\data_out[10] [7]), .I2(\data_out[10] [1]), 
            .I3(GND_net), .O(n8));   // coms.v(85[17:241])
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_851 (.I0(data_in_field[63]), .I1(data_in_field[93]), 
            .I2(data_in_field[64]), .I3(n5454), .O(n1892));   // coms.v(202[14:57])
    defparam i3_4_lut_adj_851.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_852 (.I0(delay_counter[7]), .I1(delay_counter[2]), 
            .I2(delay_counter[9]), .I3(delay_counter[0]), .O(n18_adj_1919));   // coms.v(135[5:24])
    defparam i7_4_lut_adj_852.LUT_INIT = 16'hfffe;
    SB_LUT4 n6309_bdd_4_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter[3]), .I3(n6309), .O(n6312));
    defparam n6309_bdd_4_lut_4_lut.LUT_INIT = 16'hfc07;
    SB_LUT4 i1_2_lut_adj_853 (.I0(data_in_field[124]), .I1(data_in_field[4]), 
            .I2(GND_net), .I3(GND_net), .O(n5563));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_853.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_854 (.I0(data_in_field[143]), .I1(data_in_field[115]), 
            .I2(GND_net), .I3(GND_net), .O(n5381));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_854.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_855 (.I0(data_in_field[61]), .I1(data_in_field[62]), 
            .I2(GND_net), .I3(GND_net), .O(n5384));   // coms.v(82[17:399])
    defparam i1_2_lut_adj_855.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_856 (.I0(data_in_field[100]), .I1(data_in_field[44]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1920));   // coms.v(83[17:391])
    defparam i1_2_lut_adj_856.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_857 (.I0(\data_out[10] [2]), .I1(\data_out[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1768));   // coms.v(79[17:503])
    defparam i1_2_lut_adj_857.LUT_INIT = 16'h6666;
    SB_DFF data_out_0___i1 (.Q(\data_out[10] [0]), .C(CLK_c), .D(n2484));   // coms.v(123[10] 164[6])
    SB_LUT4 i1_4_lut_adj_858 (.I0(data_in_field[122]), .I1(data_in_field[108]), 
            .I2(n4_adj_1920), .I3(data_in_field[2]), .O(n5593));   // coms.v(202[14:57])
    defparam i1_4_lut_adj_858.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(delay_counter[1]), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_1921));   // coms.v(135[5:24])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_859 (.I0(delay_counter[6]), .I1(n18_adj_1919), 
            .I2(delay_counter[3]), .I3(delay_counter[10]), .O(n20_adj_1922));   // coms.v(135[5:24])
    defparam i9_4_lut_adj_859.LUT_INIT = 16'hfffe;
    SB_CARRY add_1824_5 (.CI(n4705), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n4706));
    SB_LUT4 i1_2_lut_adj_860 (.I0(data_in_field[95]), .I1(data_in_field[80]), 
            .I2(GND_net), .I3(GND_net), .O(n2000));   // coms.v(89[18:383])
    defparam i1_2_lut_adj_860.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_861 (.I0(data_in_field[20]), .I1(data_in_field[34]), 
            .I2(data_in_field[132]), .I3(GND_net), .O(n1969));   // coms.v(202[14:57])
    defparam i2_3_lut_adj_861.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_862 (.I0(delay_counter[4]), .I1(n20_adj_1922), 
            .I2(n16_adj_1921), .I3(delay_counter[8]), .O(n21));   // coms.v(135[5:24])
    defparam i10_4_lut_adj_862.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_863 (.I0(data_in_field[66]), .I1(data_in_field[52]), 
            .I2(GND_net), .I3(GND_net), .O(n2021));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_863.LUT_INIT = 16'h6666;
    SB_LUT4 i2438_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[3] [3]), .I3(data_in_field[27]), .O(n2689));
    defparam i2438_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n2511));   // coms.v(174[10] 182[6])
    SB_LUT4 i3_4_lut_adj_864 (.I0(data_in_field[10]), .I1(data_in_field[40]), 
            .I2(data_in_field[26]), .I3(n2021), .O(n2074));   // coms.v(202[14:57])
    defparam i3_4_lut_adj_864.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_865 (.I0(n21), .I1(n4333), .I2(GND_net), .I3(GND_net), 
            .O(n4334));   // coms.v(135[5:24])
    defparam i1_2_lut_adj_865.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_866 (.I0(data_in_field[79]), .I1(data_in_field[49]), 
            .I2(GND_net), .I3(GND_net), .O(n5454));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_866.LUT_INIT = 16'h6666;
    SB_LUT4 i2437_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[3] [2]), .I3(data_in_field[26]), .O(n2688));
    defparam i2437_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2436_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[3] [1]), .I3(data_in_field[25]), .O(n2687));
    defparam i2436_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_867 (.I0(data_in_field[27]), .I1(n1926), .I2(GND_net), 
            .I3(GND_net), .O(n5469));   // coms.v(92[18:361])
    defparam i1_2_lut_adj_867.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_868 (.I0(n2074), .I1(data_in_field[24]), .I2(GND_net), 
            .I3(GND_net), .O(n5581));   // coms.v(82[17:399])
    defparam i1_2_lut_adj_868.LUT_INIT = 16'h6666;
    SB_LUT4 i2435_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[3] [0]), .I3(data_in_field[24]), .O(n2686));
    defparam i2435_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_869 (.I0(n2125), .I1(data_in_field[3]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_1923));   // coms.v(82[17:399])
    defparam i1_2_lut_adj_869.LUT_INIT = 16'h6666;
    SB_LUT4 add_1824_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n4708), .O(tx_transmit_N_568[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1824_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_870 (.I0(data_in_field[83]), .I1(n5469), .I2(n5454), 
            .I3(n6_adj_1923), .O(n5548));   // coms.v(82[17:399])
    defparam i4_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i2434_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[2] [7]), .I3(data_in_field[23]), .O(n2685));
    defparam i2434_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_871 (.I0(n1835), .I1(n2104), .I2(n1969), .I3(n1913), 
            .O(n5497));   // coms.v(202[14:57])
    defparam i3_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 data_527_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(data[4]), 
            .I3(n4742), .O(n69[4])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_528_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(delay_counter[4]), 
            .I3(n4757), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2433_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[2] [6]), .I3(data_in_field[22]), .O(n2684));
    defparam i2433_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2432_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[2] [5]), .I3(data_in_field[21]), .O(n2683));
    defparam i2432_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5704 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[16]), .I2(data_in_field[24]), .I3(byte_transmit_counter2[1]), 
            .O(n6039));
    defparam byte_transmit_counter2_0__bdd_4_lut_5704.LUT_INIT = 16'he4aa;
    SB_CARRY delay_counter_528_add_4_6 (.CI(n4757), .I0(GND_net), .I1(delay_counter[4]), 
            .CO(n4758));
    SB_CARRY data_527_add_4_6 (.CI(n4742), .I0(GND_net), .I1(data[4]), 
            .CO(n4743));
    SB_LUT4 add_1824_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n4704), .O(tx_transmit_N_568[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1824_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_872 (.I0(data_in_field[81]), .I1(data_in_field[111]), 
            .I2(data_in_field[47]), .I3(GND_net), .O(n2134));   // coms.v(86[17:391])
    defparam i2_3_lut_adj_872.LUT_INIT = 16'h9696;
    SB_LUT4 data_527_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(data[3]), 
            .I3(n4741), .O(n69[3])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_873 (.I0(\data_out[10] [1]), .I1(\data_out[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5482));   // coms.v(85[17:241])
    defparam i1_2_lut_adj_873.LUT_INIT = 16'h6666;
    SB_CARRY add_1824_8 (.CI(n4708), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n4709));
    SB_LUT4 n6039_bdd_4_lut (.I0(n6039), .I1(data_in_field[8]), .I2(data_in_field[0]), 
            .I3(byte_transmit_counter2[1]), .O(n5788));
    defparam n6039_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY data_527_add_4_5 (.CI(n4741), .I0(GND_net), .I1(data[3]), 
            .CO(n4742));
    SB_LUT4 i2431_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[2] [4]), .I3(data_in_field[20]), .O(n2682));
    defparam i2431_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2430_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[2] [3]), .I3(data_in_field[19]), .O(n2681));
    defparam i2430_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2429_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[2] [2]), .I3(data_in_field[18]), .O(n2680));
    defparam i2429_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_874 (.I0(n5509), .I1(data_in_field[92]), .I2(data_in_field[78]), 
            .I3(GND_net), .O(n2053));   // coms.v(89[18:383])
    defparam i2_3_lut_adj_874.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_875 (.I0(data_in_field[72]), .I1(data_in_field[42]), 
            .I2(GND_net), .I3(GND_net), .O(n2068));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_875.LUT_INIT = 16'h6666;
    SB_LUT4 data_527_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(data[2]), 
            .I3(n4740), .O(n69[2])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2428_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[2] [1]), .I3(data_in_field[17]), .O(n2679));
    defparam i2428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2427_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[2] [0]), .I3(data_in_field[16]), .O(n2678));
    defparam i2427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_2_lut (.I0(\data_in[1] [2]), .I1(\data_in[0] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_1924));   // coms.v(197[12:70])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(CLK_c), .D(n2527));   // coms.v(174[10] 182[6])
    SB_LUT4 i2426_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[1] [7]), .I3(data_in_field[15]), .O(n2677));
    defparam i2426_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_876 (.I0(\data_in[2] [6]), .I1(\data_in[3] [0]), 
            .I2(\data_in[3] [5]), .I3(\data_in[3] [4]), .O(n28_adj_1925));   // coms.v(197[12:70])
    defparam i12_4_lut_adj_876.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_877 (.I0(\data_in[1] [7]), .I1(\data_in[1] [5]), 
            .I2(\data_in[0] [6]), .I3(\data_in[0] [7]), .O(n28_adj_1926));
    defparam i12_4_lut_adj_877.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_878 (.I0(data_in_field[87]), .I1(data_in_field[128]), 
            .I2(GND_net), .I3(GND_net), .O(n1965));   // coms.v(83[17:391])
    defparam i1_2_lut_adj_878.LUT_INIT = 16'h6666;
    SB_LUT4 i2425_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[1] [6]), .I3(data_in_field[14]), .O(n2676));
    defparam i2425_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(CLK_c), .D(n2528));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(CLK_c), .D(n2529));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n2530));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(CLK_c), .D(n2531));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(CLK_c), .D(n2532));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(CLK_c), .D(n2533));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i33 (.Q(\data_in[4] [0]), .C(CLK_c), .D(n2534));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i34 (.Q(\data_in[4] [1]), .C(CLK_c), .D(n2535));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i35 (.Q(\data_in[4] [2]), .C(CLK_c), .D(n2536));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i36 (.Q(\data_in[4] [3]), .C(CLK_c), .D(n2537));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i37 (.Q(\data_in[4] [4]), .C(CLK_c), .D(n2538));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i38 (.Q(\data_in[4] [5]), .C(CLK_c), .D(n2539));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i39 (.Q(\data_in[4] [6]), .C(CLK_c), .D(n2540));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i40 (.Q(\data_in[4] [7]), .C(CLK_c), .D(n2541));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i41 (.Q(\data_in[5] [0]), .C(CLK_c), .D(n2542));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i42 (.Q(\data_in[5] [1]), .C(CLK_c), .D(n2543));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i43 (.Q(\data_in[5] [2]), .C(CLK_c), .D(n2544));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i44 (.Q(\data_in[5] [3]), .C(CLK_c), .D(n2545));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i45 (.Q(\data_in[5] [4]), .C(CLK_c), .D(n2546));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i46 (.Q(\data_in[5] [5]), .C(CLK_c), .D(n2547));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i54 (.Q(\data_in[6] [5]), .C(CLK_c), .D(n2555));   // coms.v(174[10] 182[6])
    SB_LUT4 i2_3_lut_adj_879 (.I0(data_in_field[14]), .I1(data_in_field[106]), 
            .I2(data_in_field[134]), .I3(GND_net), .O(n5554));   // coms.v(202[14:57])
    defparam i2_3_lut_adj_879.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_880 (.I0(data_in_field[56]), .I1(data_in_field[70]), 
            .I2(data_in_field[84]), .I3(GND_net), .O(n5494));   // coms.v(202[14:57])
    defparam i2_3_lut_adj_880.LUT_INIT = 16'h9696;
    SB_LUT4 i2424_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[1] [5]), .I3(data_in_field[13]), .O(n2675));
    defparam i2424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_881 (.I0(data_in_field[76]), .I1(data_in_field[126]), 
            .I2(data_in_field[112]), .I3(GND_net), .O(n5524));   // coms.v(202[14:57])
    defparam i2_3_lut_adj_881.LUT_INIT = 16'h9696;
    SB_LUT4 i2423_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[1] [4]), .I3(data_in_field[12]), .O(n2674));
    defparam i2423_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_882 (.I0(\data_in[2] [0]), .I1(\data_in[2] [3]), 
            .I2(\data_in[0] [3]), .I3(\data_in[2] [5]), .O(n26));
    defparam i10_4_lut_adj_882.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_883 (.I0(data_in_field[6]), .I1(data_in_field[104]), 
            .I2(GND_net), .I3(GND_net), .O(n2143));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_883.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_884 (.I0(n5391), .I1(n5524), .I2(n5494), .I3(n5554), 
            .O(n26_adj_1927));   // coms.v(202[14:57])
    defparam i11_4_lut_adj_884.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i55 (.Q(\data_in[6] [6]), .C(CLK_c), .D(n2556));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i56 (.Q(\data_in[6] [7]), .C(CLK_c), .D(n2557));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i57 (.Q(\data_in[7] [0]), .C(CLK_c), .D(n2558));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i58 (.Q(\data_in[7] [1]), .C(CLK_c), .D(n2559));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i59 (.Q(\data_in[7] [2]), .C(CLK_c), .D(n2560));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i60 (.Q(\data_in[7] [3]), .C(CLK_c), .D(n2561));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i61 (.Q(\data_in[7] [4]), .C(CLK_c), .D(n2562));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i62 (.Q(\data_in[7] [5]), .C(CLK_c), .D(n2563));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i63 (.Q(\data_in[7] [6]), .C(CLK_c), .D(n2564));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i64 (.Q(\data_in[7] [7]), .C(CLK_c), .D(n2565));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i65 (.Q(\data_in[8] [0]), .C(CLK_c), .D(n2566));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i66 (.Q(\data_in[8] [1]), .C(CLK_c), .D(n2567));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i67 (.Q(\data_in[8] [2]), .C(CLK_c), .D(n2568));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i68 (.Q(\data_in[8] [3]), .C(CLK_c), .D(n2569));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i69 (.Q(\data_in[8] [4]), .C(CLK_c), .D(n2570));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i70 (.Q(\data_in[8] [5]), .C(CLK_c), .D(n2571));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i71 (.Q(\data_in[8] [6]), .C(CLK_c), .D(n2572));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i72 (.Q(\data_in[8] [7]), .C(CLK_c), .D(n2573));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i73 (.Q(\data_in[9] [0]), .C(CLK_c), .D(n2574));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i74 (.Q(\data_in[9] [1]), .C(CLK_c), .D(n2575));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i75 (.Q(\data_in[9] [2]), .C(CLK_c), .D(n2576));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i76 (.Q(\data_in[9] [3]), .C(CLK_c), .D(n2577));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i77 (.Q(\data_in[9] [4]), .C(CLK_c), .D(n2578));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i78 (.Q(\data_in[9] [5]), .C(CLK_c), .D(n2579));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i79 (.Q(\data_in[9] [6]), .C(CLK_c), .D(n2580));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i80 (.Q(\data_in[9] [7]), .C(CLK_c), .D(n2581));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i81 (.Q(\data_in[10] [0]), .C(CLK_c), .D(n2582));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i82 (.Q(\data_in[10] [1]), .C(CLK_c), .D(n2583));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i83 (.Q(\data_in[10] [2]), .C(CLK_c), .D(n2584));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i84 (.Q(\data_in[10] [3]), .C(CLK_c), .D(n2585));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i85 (.Q(\data_in[10] [4]), .C(CLK_c), .D(n2586));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i86 (.Q(\data_in[10] [5]), .C(CLK_c), .D(n2587));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i88 (.Q(\data_in[10] [7]), .C(CLK_c), .D(n2589));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i89 (.Q(\data_in[11] [0]), .C(CLK_c), .D(n2590));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i90 (.Q(\data_in[11] [1]), .C(CLK_c), .D(n2591));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i91 (.Q(\data_in[11] [2]), .C(CLK_c), .D(n2592));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i92 (.Q(\data_in[11] [3]), .C(CLK_c), .D(n2593));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i93 (.Q(\data_in[11] [4]), .C(CLK_c), .D(n2594));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i94 (.Q(\data_in[11] [5]), .C(CLK_c), .D(n2595));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i95 (.Q(\data_in[11] [6]), .C(CLK_c), .D(n2596));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i96 (.Q(\data_in[11] [7]), .C(CLK_c), .D(n2597));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i97 (.Q(\data_in[12] [0]), .C(CLK_c), .D(n2598));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i98 (.Q(\data_in[12] [1]), .C(CLK_c), .D(n2599));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i99 (.Q(\data_in[12] [2]), .C(CLK_c), .D(n2600));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i100 (.Q(\data_in[12] [3]), .C(CLK_c), .D(n2601));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i101 (.Q(\data_in[12] [4]), .C(CLK_c), .D(n2602));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i102 (.Q(\data_in[12] [5]), .C(CLK_c), .D(n2603));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i103 (.Q(\data_in[12] [6]), .C(CLK_c), .D(n2604));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i104 (.Q(\data_in[12] [7]), .C(CLK_c), .D(n2605));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i105 (.Q(\data_in[13] [0]), .C(CLK_c), .D(n2606));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i106 (.Q(\data_in[13] [1]), .C(CLK_c), .D(n2607));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i107 (.Q(\data_in[13] [2]), .C(CLK_c), .D(n2608));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i108 (.Q(\data_in[13] [3]), .C(CLK_c), .D(n2609));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i109 (.Q(\data_in[13] [4]), .C(CLK_c), .D(n2610));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i110 (.Q(\data_in[13] [5]), .C(CLK_c), .D(n2611));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i111 (.Q(\data_in[13] [6]), .C(CLK_c), .D(n2612));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i112 (.Q(\data_in[13] [7]), .C(CLK_c), .D(n2613));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i113 (.Q(\data_in[14] [0]), .C(CLK_c), .D(n2614));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i114 (.Q(\data_in[14] [1]), .C(CLK_c), .D(n2615));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i115 (.Q(\data_in[14] [2]), .C(CLK_c), .D(n2616));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i116 (.Q(\data_in[14] [3]), .C(CLK_c), .D(n2617));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i117 (.Q(\data_in[14] [4]), .C(CLK_c), .D(n2618));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i118 (.Q(\data_in[14] [5]), .C(CLK_c), .D(n2619));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i119 (.Q(\data_in[14] [6]), .C(CLK_c), .D(n2620));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i127 (.Q(\data_in[15] [6]), .C(CLK_c), .D(n2628));   // coms.v(174[10] 182[6])
    SB_LUT4 i11_4_lut_adj_885 (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), 
            .I2(\data_in[0] [4]), .I3(\data_in[2] [7]), .O(n27_adj_1928));
    defparam i11_4_lut_adj_885.LUT_INIT = 16'h8000;
    SB_LUT4 i9_4_lut_adj_886 (.I0(\data_in[1] [0]), .I1(\data_in[2] [2]), 
            .I2(\data_in[1] [3]), .I3(\data_in[1] [4]), .O(n25_adj_1929));
    defparam i9_4_lut_adj_886.LUT_INIT = 16'h8000;
    SB_LUT4 i9_4_lut_adj_887 (.I0(data_in_field[91]), .I1(n1965), .I2(n2068), 
            .I3(data_in_field[46]), .O(n24_adj_1930));   // coms.v(202[14:57])
    defparam i9_4_lut_adj_887.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5685 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[48]), .I2(data_in_field[56]), .I3(byte_transmit_counter2[1]), 
            .O(n6033));
    defparam byte_transmit_counter2_0__bdd_4_lut_5685.LUT_INIT = 16'he4aa;
    SB_LUT4 i2422_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[1] [3]), .I3(data_in_field[11]), .O(n2673));
    defparam i2422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_888 (.I0(data_in_field[16]), .I1(data_in_field[1]), 
            .I2(n2113), .I3(data_in_field[74]), .O(n25_adj_1931));   // coms.v(202[14:57])
    defparam i10_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_LUT4 i2421_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[1] [2]), .I3(data_in_field[10]), .O(n2672));
    defparam i2421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n6033_bdd_4_lut (.I0(n6033), .I1(data_in_field[40]), .I2(data_in_field[32]), 
            .I3(byte_transmit_counter2[1]), .O(n5791));
    defparam n6033_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 delay_counter_528_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(delay_counter[3]), 
            .I3(n4756), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2420_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[1] [1]), .I3(data_in_field[9]), .O(n2671));
    defparam i2420_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i128 (.Q(\data_in[15] [7]), .C(CLK_c), .D(n2629));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i129 (.Q(\data_in[16] [0]), .C(CLK_c), .D(n2630));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i130 (.Q(\data_in[16] [1]), .C(CLK_c), .D(n2631));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i131 (.Q(\data_in[16] [2]), .C(CLK_c), .D(n2632));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i132 (.Q(\data_in[16] [3]), .C(CLK_c), .D(n2633));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i133 (.Q(\data_in[16] [4]), .C(CLK_c), .D(n2634));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i134 (.Q(\data_in[16] [5]), .C(CLK_c), .D(n2635));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i135 (.Q(\data_in[16] [6]), .C(CLK_c), .D(n2636));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i136 (.Q(\data_in[16] [7]), .C(CLK_c), .D(n2637));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i137 (.Q(\data_in[17] [0]), .C(CLK_c), .D(n2638));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i138 (.Q(\data_in[17] [1]), .C(CLK_c), .D(n2639));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i139 (.Q(\data_in[17] [2]), .C(CLK_c), .D(n2640));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i140 (.Q(\data_in[17] [3]), .C(CLK_c), .D(n2641));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i141 (.Q(\data_in[17] [4]), .C(CLK_c), .D(n2642));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i142 (.Q(\data_in[17] [5]), .C(CLK_c), .D(n2643));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i143 (.Q(\data_in[17] [6]), .C(CLK_c), .D(n2644));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i144 (.Q(\data_in[17] [7]), .C(CLK_c), .D(n2645));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i145 (.Q(\data_in[18] [0]), .C(CLK_c), .D(n2646));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i146 (.Q(\data_in[18] [1]), .C(CLK_c), .D(n2647));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i147 (.Q(\data_in[18] [2]), .C(CLK_c), .D(n2648));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i148 (.Q(\data_in[18] [3]), .C(CLK_c), .D(n2649));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i149 (.Q(\data_in[18] [4]), .C(CLK_c), .D(n2650));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i150 (.Q(\data_in[18] [5]), .C(CLK_c), .D(n2651));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i151 (.Q(\data_in[18] [6]), .C(CLK_c), .D(n2652));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i152 (.Q(\data_in[18] [7]), .C(CLK_c), .D(n2653));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i153 (.Q(\data_in[19] [0]), .C(CLK_c), .D(n2654));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i154 (.Q(\data_in[19] [1]), .C(CLK_c), .D(n2655));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i155 (.Q(\data_in[19] [2]), .C(CLK_c), .D(n2656));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i156 (.Q(\data_in[19] [3]), .C(CLK_c), .D(n2657));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i157 (.Q(\data_in[19] [4]), .C(CLK_c), .D(n2658));   // coms.v(174[10] 182[6])
    SB_DFF data_in_frame_0___i5 (.Q(data_in_field[4]), .C(CLK_c), .D(n2666));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i6 (.Q(data_in_field[5]), .C(CLK_c), .D(n2667));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i7 (.Q(data_in_field[6]), .C(CLK_c), .D(n2668));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i8 (.Q(data_in_field[7]), .C(CLK_c), .D(n2669));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i9 (.Q(data_in_field[8]), .C(CLK_c), .D(n2670));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i10 (.Q(data_in_field[9]), .C(CLK_c), .D(n2671));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i11 (.Q(data_in_field[10]), .C(CLK_c), .D(n2672));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i12 (.Q(data_in_field[11]), .C(CLK_c), .D(n2673));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i13 (.Q(data_in_field[12]), .C(CLK_c), .D(n2674));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i14 (.Q(data_in_field[13]), .C(CLK_c), .D(n2675));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i15 (.Q(data_in_field[14]), .C(CLK_c), .D(n2676));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i16 (.Q(data_in_field[15]), .C(CLK_c), .D(n2677));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i17 (.Q(data_in_field[16]), .C(CLK_c), .D(n2678));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i18 (.Q(data_in_field[17]), .C(CLK_c), .D(n2679));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i19 (.Q(data_in_field[18]), .C(CLK_c), .D(n2680));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i20 (.Q(data_in_field[19]), .C(CLK_c), .D(n2681));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i21 (.Q(data_in_field[20]), .C(CLK_c), .D(n2682));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i22 (.Q(data_in_field[21]), .C(CLK_c), .D(n2683));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i23 (.Q(data_in_field[22]), .C(CLK_c), .D(n2684));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i24 (.Q(data_in_field[23]), .C(CLK_c), .D(n2685));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i25 (.Q(data_in_field[24]), .C(CLK_c), .D(n2686));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i26 (.Q(data_in_field[25]), .C(CLK_c), .D(n2687));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i27 (.Q(data_in_field[26]), .C(CLK_c), .D(n2688));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i28 (.Q(data_in_field[27]), .C(CLK_c), .D(n2689));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i29 (.Q(data_in_field[28]), .C(CLK_c), .D(n2690));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i30 (.Q(data_in_field[29]), .C(CLK_c), .D(n2691));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i31 (.Q(data_in_field[30]), .C(CLK_c), .D(n2692));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i32 (.Q(data_in_field[31]), .C(CLK_c), .D(n2693));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i33 (.Q(data_in_field[32]), .C(CLK_c), .D(n2694));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i34 (.Q(data_in_field[33]), .C(CLK_c), .D(n2695));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i35 (.Q(data_in_field[34]), .C(CLK_c), .D(n2696));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i36 (.Q(data_in_field[35]), .C(CLK_c), .D(n2697));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i37 (.Q(data_in_field[36]), .C(CLK_c), .D(n2698));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i38 (.Q(data_in_field[37]), .C(CLK_c), .D(n2699));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i39 (.Q(data_in_field[38]), .C(CLK_c), .D(n2700));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i40 (.Q(data_in_field[39]), .C(CLK_c), .D(n2701));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i41 (.Q(data_in_field[40]), .C(CLK_c), .D(n2702));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i42 (.Q(data_in_field[41]), .C(CLK_c), .D(n2703));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i43 (.Q(data_in_field[42]), .C(CLK_c), .D(n2704));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i44 (.Q(data_in_field[43]), .C(CLK_c), .D(n2705));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i45 (.Q(data_in_field[44]), .C(CLK_c), .D(n2706));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i46 (.Q(data_in_field[45]), .C(CLK_c), .D(n2707));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i47 (.Q(data_in_field[46]), .C(CLK_c), .D(n2708));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i48 (.Q(data_in_field[47]), .C(CLK_c), .D(n2709));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i49 (.Q(data_in_field[48]), .C(CLK_c), .D(n2710));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i50 (.Q(data_in_field[49]), .C(CLK_c), .D(n2711));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i51 (.Q(data_in_field[50]), .C(CLK_c), .D(n2712));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i52 (.Q(data_in_field[51]), .C(CLK_c), .D(n2713));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i53 (.Q(data_in_field[52]), .C(CLK_c), .D(n2714));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i54 (.Q(data_in_field[53]), .C(CLK_c), .D(n2715));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i55 (.Q(data_in_field[54]), .C(CLK_c), .D(n2716));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i56 (.Q(data_in_field[55]), .C(CLK_c), .D(n2717));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i57 (.Q(data_in_field[56]), .C(CLK_c), .D(n2718));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i58 (.Q(data_in_field[57]), .C(CLK_c), .D(n2719));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i59 (.Q(data_in_field[58]), .C(CLK_c), .D(n2720));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i60 (.Q(data_in_field[59]), .C(CLK_c), .D(n2721));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i61 (.Q(data_in_field[60]), .C(CLK_c), .D(n2722));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i62 (.Q(data_in_field[61]), .C(CLK_c), .D(n2723));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i63 (.Q(data_in_field[62]), .C(CLK_c), .D(n2724));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i64 (.Q(data_in_field[63]), .C(CLK_c), .D(n2725));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i65 (.Q(data_in_field[64]), .C(CLK_c), .D(n2726));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i66 (.Q(data_in_field[65]), .C(CLK_c), .D(n2727));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i67 (.Q(data_in_field[66]), .C(CLK_c), .D(n2728));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i68 (.Q(data_in_field[67]), .C(CLK_c), .D(n2729));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i69 (.Q(data_in_field[68]), .C(CLK_c), .D(n2730));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i70 (.Q(data_in_field[69]), .C(CLK_c), .D(n2731));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i71 (.Q(data_in_field[70]), .C(CLK_c), .D(n2732));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i72 (.Q(data_in_field[71]), .C(CLK_c), .D(n2733));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i73 (.Q(data_in_field[72]), .C(CLK_c), .D(n2734));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i74 (.Q(data_in_field[73]), .C(CLK_c), .D(n2735));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i75 (.Q(data_in_field[74]), .C(CLK_c), .D(n2736));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i76 (.Q(data_in_field[75]), .C(CLK_c), .D(n2737));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i77 (.Q(data_in_field[76]), .C(CLK_c), .D(n2738));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i78 (.Q(data_in_field[77]), .C(CLK_c), .D(n2739));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i79 (.Q(data_in_field[78]), .C(CLK_c), .D(n2740));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i80 (.Q(data_in_field[79]), .C(CLK_c), .D(n2741));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i81 (.Q(data_in_field[80]), .C(CLK_c), .D(n2742));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i82 (.Q(data_in_field[81]), .C(CLK_c), .D(n2743));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i83 (.Q(data_in_field[82]), .C(CLK_c), .D(n2744));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i84 (.Q(data_in_field[83]), .C(CLK_c), .D(n2745));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i85 (.Q(data_in_field[84]), .C(CLK_c), .D(n2746));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i86 (.Q(data_in_field[85]), .C(CLK_c), .D(n2747));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i87 (.Q(data_in_field[86]), .C(CLK_c), .D(n2748));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i88 (.Q(data_in_field[87]), .C(CLK_c), .D(n2749));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i89 (.Q(data_in_field[88]), .C(CLK_c), .D(n2750));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i90 (.Q(data_in_field[89]), .C(CLK_c), .D(n2751));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i91 (.Q(data_in_field[90]), .C(CLK_c), .D(n2752));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i92 (.Q(data_in_field[91]), .C(CLK_c), .D(n2753));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i93 (.Q(data_in_field[92]), .C(CLK_c), .D(n2754));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i94 (.Q(data_in_field[93]), .C(CLK_c), .D(n2755));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i95 (.Q(data_in_field[94]), .C(CLK_c), .D(n2756));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i96 (.Q(data_in_field[95]), .C(CLK_c), .D(n2757));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i97 (.Q(data_in_field[96]), .C(CLK_c), .D(n2758));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i98 (.Q(data_in_field[97]), .C(CLK_c), .D(n2759));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i99 (.Q(data_in_field[98]), .C(CLK_c), .D(n2760));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i100 (.Q(data_in_field[99]), .C(CLK_c), .D(n2761));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i101 (.Q(data_in_field[100]), .C(CLK_c), .D(n2762));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i102 (.Q(data_in_field[101]), .C(CLK_c), .D(n2763));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i103 (.Q(data_in_field[102]), .C(CLK_c), .D(n2764));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i104 (.Q(data_in_field[103]), .C(CLK_c), .D(n2765));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i105 (.Q(data_in_field[104]), .C(CLK_c), .D(n2766));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i106 (.Q(data_in_field[105]), .C(CLK_c), .D(n2767));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i107 (.Q(data_in_field[106]), .C(CLK_c), .D(n2768));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i108 (.Q(data_in_field[107]), .C(CLK_c), .D(n2769));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i109 (.Q(data_in_field[108]), .C(CLK_c), .D(n2770));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i110 (.Q(data_in_field[109]), .C(CLK_c), .D(n2771));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i111 (.Q(data_in_field[110]), .C(CLK_c), .D(n2772));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i112 (.Q(data_in_field[111]), .C(CLK_c), .D(n2773));   // coms.v(192[10] 220[6])
    SB_DFF data_in_frame_0___i113 (.Q(data_in_field[112]), .C(CLK_c), .D(n2774));   // coms.v(192[10] 220[6])
    SB_DFF data_out_0___i6 (.Q(\data_out[10] [5]), .C(CLK_c), .D(n2841));   // coms.v(123[10] 164[6])
    SB_CARRY delay_counter_528_add_4_5 (.CI(n4756), .I0(GND_net), .I1(delay_counter[3]), 
            .CO(n4757));
    SB_DFF data_out_0___i21 (.Q(\data_out[18] [4]), .C(CLK_c), .D(n2856));   // coms.v(123[10] 164[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(CLK_c), .D(n2384));   // coms.v(174[10] 182[6])
    SB_LUT4 i14_4_lut_adj_889 (.I0(n23_adj_1935), .I1(n25_adj_1931), .I2(n24_adj_1930), 
            .I3(n26_adj_1927), .O(n1814));   // coms.v(202[14:57])
    defparam i14_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_890 (.I0(data_in_field[139]), .I1(data_in_field[19]), 
            .I2(data_in_field[77]), .I3(GND_net), .O(n5372));   // coms.v(202[14:57])
    defparam i2_3_lut_adj_890.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i134 (.Q(data_in_field[133]), .C(CLK_c), .D(n2795));   // coms.v(192[10] 220[6])
    SB_LUT4 i2_3_lut_adj_891 (.I0(data_in_field[13]), .I1(data_in_field[69]), 
            .I2(data_in_field[110]), .I3(GND_net), .O(n2043));   // coms.v(93[18:87])
    defparam i2_3_lut_adj_891.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_892 (.I0(data_in_field[61]), .I1(data_in_field[140]), 
            .I2(GND_net), .I3(GND_net), .O(n5391));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_892.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_893 (.I0(data_in_field[33]), .I1(data_in_field[92]), 
            .I2(data_in_field[91]), .I3(GND_net), .O(n5403));   // coms.v(86[17:391])
    defparam i2_3_lut_adj_893.LUT_INIT = 16'h9696;
    SB_DFF \FRAME_MATCHER.wait_for_transmission_1803  (.Q(\FRAME_MATCHER.wait_for_transmission ), 
           .C(CLK_c), .D(n6));   // coms.v(192[10] 220[6])
    SB_LUT4 i1_2_lut_adj_894 (.I0(\data_out[10] [4]), .I1(n5409), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3));
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h6666;
    SB_LUT4 delay_counter_528_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(delay_counter[2]), 
            .I3(n4755), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_528_add_4_4 (.CI(n4755), .I0(GND_net), .I1(delay_counter[2]), 
            .CO(n4756));
    SB_LUT4 i2_3_lut_adj_895 (.I0(n5403), .I1(data_in_field[93]), .I2(n1866), 
            .I3(GND_net), .O(n1855));   // coms.v(86[17:391])
    defparam i2_3_lut_adj_895.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_896 (.I0(data_in_field[125]), .I1(data_in_field[35]), 
            .I2(GND_net), .I3(GND_net), .O(n5476));   // coms.v(93[18:87])
    defparam i1_2_lut_adj_896.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_897 (.I0(\data_out[11] [5]), .I1(\data_out[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n5415));
    defparam i1_2_lut_adj_897.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(n2155), .I1(data_in_field[31]), .I2(data_in_field[73]), 
            .I3(data_in_field[137]), .O(n2012));   // coms.v(82[17:399])
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_898 (.I0(data_in_field[91]), .I1(data_in_field[127]), 
            .I2(GND_net), .I3(GND_net), .O(n1908));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h6666;
    SB_LUT4 i2419_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[1] [0]), .I3(data_in_field[8]), .O(n2670));
    defparam i2419_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_0___i20 (.Q(\data_out[18] [3]), .C(CLK_c), .D(n2855));   // coms.v(123[10] 164[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(data_in_field[109]), .I1(data_in_field[45]), 
            .I2(data_in_field[64]), .I3(n5476), .O(n31_adj_1896));   // coms.v(202[14:57])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF delay_counter_528__i4 (.Q(delay_counter[4]), .C(CLK_c), .D(n1[4]));   // coms.v(159[11] 161[5])
    SB_DFF data_in_frame_0___i133 (.Q(data_in_field[132]), .C(CLK_c), .D(n2794));   // coms.v(192[10] 220[6])
    SB_LUT4 i8_3_lut_4_lut (.I0(data_in_field[108]), .I1(data_in_field[106]), 
            .I2(n5560), .I3(data_in_field[2]), .O(n34));   // coms.v(202[14:57])
    defparam i8_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_899 (.I0(data_in_field[93]), .I1(data_in_field[37]), 
            .I2(GND_net), .I3(GND_net), .O(n1955));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h6666;
    SB_LUT4 i1_rep_100_2_lut_3_lut (.I0(data_in_field[109]), .I1(data_in_field[45]), 
            .I2(n2065), .I3(GND_net), .O(n6414));   // coms.v(202[14:57])
    defparam i1_rep_100_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_out[10] [7]), .I1(\data_out[11] [1]), 
            .I2(\data_out[11] [4]), .I3(n5409), .O(n4_adj_4));   // coms.v(81[17:257])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_900 (.I0(n5436), .I1(n1955), .I2(n1948), .I3(GND_net), 
            .O(n5509));   // coms.v(89[18:383])
    defparam i2_3_lut_adj_900.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_901 (.I0(data_in_field[40]), .I1(data_in_field[98]), 
            .I2(data_in_field[100]), .I3(n2101), .O(n6_adj_1917));   // coms.v(202[14:57])
    defparam i1_2_lut_3_lut_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_902 (.I0(data_in_field[40]), .I1(data_in_field[98]), 
            .I2(data_in_field[100]), .I3(data_in_field[23]), .O(n18_adj_1938));   // coms.v(202[14:57])
    defparam i1_2_lut_3_lut_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_903 (.I0(n2080), .I1(n1889), .I2(n2012), .I3(data_in_field[30]), 
            .O(n5491));   // coms.v(82[17:399])
    defparam i3_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_904 (.I0(\data_out[11] [4]), .I1(n5409), .I2(GND_net), 
            .I3(GND_net), .O(n1991));   // coms.v(79[17:447])
    defparam i1_2_lut_adj_904.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_905 (.I0(data_in_field[75]), .I1(data_in_field[90]), 
            .I2(data_in_field[89]), .I3(GND_net), .O(n2065));   // coms.v(82[17:399])
    defparam i1_2_lut_3_lut_adj_905.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5680 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[80]), .I2(data_in_field[88]), .I3(byte_transmit_counter2[1]), 
            .O(n6027));
    defparam byte_transmit_counter2_0__bdd_4_lut_5680.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut (.I0(data_in_field[72]), .I1(data_in_field[16]), 
            .I2(data_in_field[31]), .I3(data_in_field[136]), .O(n6_adj_1939));   // coms.v(83[17:391])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_906 (.I0(data_in_field[50]), .I1(data_in_field[46]), 
            .I2(data_in_field[110]), .I3(GND_net), .O(n5533));   // coms.v(202[14:57])
    defparam i1_2_lut_3_lut_adj_906.LUT_INIT = 16'h9696;
    SB_DFF delay_counter_528__i10 (.Q(delay_counter[10]), .C(CLK_c), .D(n1[10]));   // coms.v(159[11] 161[5])
    SB_DFF data_out_0___i31 (.Q(\data_out[19] [6]), .C(CLK_c), .D(n2866));   // coms.v(123[10] 164[6])
    SB_LUT4 i1_2_lut_adj_907 (.I0(data_in_field[96]), .I1(data_in_field[95]), 
            .I2(GND_net), .I3(GND_net), .O(n5427));   // coms.v(92[18:361])
    defparam i1_2_lut_adj_907.LUT_INIT = 16'h6666;
    SB_DFF data_out_0___i5 (.Q(\data_out[10] [4]), .C(CLK_c), .D(n2840));   // coms.v(123[10] 164[6])
    SB_DFF data_in_frame_0___i130 (.Q(data_in_field[129]), .C(CLK_c), .D(n2791));   // coms.v(192[10] 220[6])
    SB_LUT4 i2418_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[0] [7]), .I3(data_in_field[7]), .O(n2669));
    defparam i2418_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i129 (.Q(data_in_field[128]), .C(CLK_c), .D(n2790));   // coms.v(192[10] 220[6])
    SB_LUT4 i1_2_lut_4_lut_adj_908 (.I0(data_in_field[74]), .I1(data_in_field[78]), 
            .I2(data_in_field[18]), .I3(data_in_field[76]), .O(n1958));   // coms.v(202[14:57])
    defparam i1_2_lut_4_lut_adj_908.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_909 (.I0(data_in_field[97]), .I1(data_in_field[83]), 
            .I2(GND_net), .I3(GND_net), .O(n1886));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_909.LUT_INIT = 16'h6666;
    SB_LUT4 delay_counter_528_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(delay_counter[1]), 
            .I3(n4754), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2417_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[0] [6]), .I3(data_in_field[6]), .O(n2668));
    defparam i2417_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_0___i16 (.Q(\data_out[11] [7]), .C(CLK_c), .D(n2851));   // coms.v(123[10] 164[6])
    SB_DFF data_out_0___i19 (.Q(\data_out[18] [2]), .C(CLK_c), .D(n2854));   // coms.v(123[10] 164[6])
    SB_LUT4 i2_3_lut_adj_910 (.I0(data_in_field[65]), .I1(data_in_field[129]), 
            .I2(data_in_field[69]), .I3(GND_net), .O(n5569));   // coms.v(89[18:383])
    defparam i2_3_lut_adj_910.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_911 (.I0(data_in_field[66]), .I1(data_in_field[79]), 
            .I2(data_in_field[94]), .I3(GND_net), .O(n5545));   // coms.v(202[14:57])
    defparam i2_3_lut_adj_911.LUT_INIT = 16'h9696;
    SB_LUT4 i2416_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[0] [5]), .I3(data_in_field[5]), .O(n2667));
    defparam i2416_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2415_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[0] [4]), .I3(data_in_field[4]), .O(n2666));
    defparam i2415_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_912 (.I0(\data_in[3] [1]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [2]), .O(n26_adj_1940));   // coms.v(197[12:70])
    defparam i10_4_lut_adj_912.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_913 (.I0(data_in_field[38]), .I1(data_in_field[24]), 
            .I2(data_in_field[136]), .I3(data_in_field[39]), .O(n5560));   // coms.v(202[14:57])
    defparam i1_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(CLK_c), .D(n2510));   // coms.v(174[10] 182[6])
    SB_LUT4 i2568_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[19] [5]), .I3(\data_in_frame[19] [5]), .O(n2819));
    defparam i2568_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2561_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[18] [6]), .I3(\data_in_frame[18] [6]), .O(n2812));
    defparam i2561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF delay_counter_528__i8 (.Q(delay_counter[8]), .C(CLK_c), .D(n1[8]));   // coms.v(159[11] 161[5])
    SB_DFF delay_counter_528__i7 (.Q(delay_counter[7]), .C(CLK_c), .D(n1[7]));   // coms.v(159[11] 161[5])
    SB_DFF delay_counter_528__i9 (.Q(delay_counter[9]), .C(CLK_c), .D(n1[9]));   // coms.v(159[11] 161[5])
    SB_DFF delay_counter_528__i3 (.Q(delay_counter[3]), .C(CLK_c), .D(n1[3]));   // coms.v(159[11] 161[5])
    SB_DFF data_out_0___i11 (.Q(\data_out[11] [2]), .C(CLK_c), .D(n2846));   // coms.v(123[10] 164[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(CLK_c), 
           .D(n2821));   // coms.v(192[10] 220[6])
    SB_LUT4 i2557_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[18] [2]), .I3(\data_in_frame[18] [2]), .O(n2808));
    defparam i2557_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2547_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[17] [0]), .I3(data_in_field[136]), .O(n2798));
    defparam i2547_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2548_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[17] [1]), .I3(data_in_field[137]), .O(n2799));
    defparam i2548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n6009_bdd_4_lut (.I0(n6009), .I1(data_in_field[15]), .I2(data_in_field[7]), 
            .I3(byte_transmit_counter2[1]), .O(n6012));
    defparam n6009_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_914 (.I0(data_in_field[94]), .I1(data_in_field[36]), 
            .I2(data_in_field[22]), .I3(GND_net), .O(n5436));   // coms.v(89[18:383])
    defparam i1_2_lut_3_lut_adj_914.LUT_INIT = 16'h9696;
    SB_LUT4 i2551_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[17] [4]), .I3(data_in_field[140]), .O(n2802));
    defparam i2551_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2552_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[17] [5]), .I3(data_in_field[141]), .O(n2803));
    defparam i2552_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_915 (.I0(data_in_field[106]), .I1(n5560), .I2(GND_net), 
            .I3(GND_net), .O(n5412));   // coms.v(89[18:383])
    defparam i1_2_lut_adj_915.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_916 (.I0(data_in_field[122]), .I1(data_in_field[99]), 
            .I2(GND_net), .I3(GND_net), .O(n5375));   // coms.v(82[17:399])
    defparam i1_2_lut_adj_916.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_917 (.I0(data_in_field[97]), .I1(data_in_field[82]), 
            .I2(data_in_field[96]), .I3(GND_net), .O(n1948));   // coms.v(93[18:87])
    defparam i2_3_lut_adj_917.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n2509));   // coms.v(174[10] 182[6])
    SB_LUT4 i1_2_lut_adj_918 (.I0(data_in_field[94]), .I1(data_in_field[116]), 
            .I2(GND_net), .I3(GND_net), .O(n1779));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_918.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut (.I0(data_in_field[60]), .I1(data_in_field[0]), 
            .I2(n2030), .I3(n1917), .O(n5466));   // coms.v(202[14:57])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_919 (.I0(data_in_field[122]), .I1(data_in_field[99]), 
            .I2(data_in_field[86]), .I3(data_in_field[71]), .O(n1889));   // coms.v(82[17:399])
    defparam i2_3_lut_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_920 (.I0(data_in_field[97]), .I1(data_in_field[83]), 
            .I2(n1942), .I3(data_in_field[85]), .O(n5578));   // coms.v(92[18:361])
    defparam i2_3_lut_4_lut_adj_920.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_921 (.I0(data_in_field[81]), .I1(data_in_field[96]), 
            .I2(data_in_field[95]), .I3(GND_net), .O(n1942));   // coms.v(92[18:361])
    defparam i1_2_lut_3_lut_adj_921.LUT_INIT = 16'h9696;
    SB_LUT4 add_1824_2_lut (.I0(n4334), .I1(byte_transmit_counter[0]), .I2(n50_adj_1875), 
            .I3(GND_net), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1824_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_4_lut_adj_922 (.I0(data_in_field[107]), .I1(data_in_field[15]), 
            .I2(data_in_field[121]), .I3(data_in_field[1]), .O(n2080));   // coms.v(202[14:57])
    defparam i2_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_CARRY add_1824_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(n50_adj_1875), 
            .CO(n4703));
    SB_LUT4 i2_3_lut_4_lut_adj_923 (.I0(data_in_field[135]), .I1(data_in_field[92]), 
            .I2(data_in_field[91]), .I3(data_in_field[127]), .O(n5418));   // coms.v(202[14:57])
    defparam i2_3_lut_4_lut_adj_923.LUT_INIT = 16'h6996;
    SB_LUT4 i2134_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[0] [0]), .I3(data_in_field[0]), .O(n2385));
    defparam i2134_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_924 (.I0(data_in_field[129]), .I1(data_in_field[17]), 
            .I2(GND_net), .I3(GND_net), .O(n2155));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut (.I0(byte_transmit_counter2[0]), 
            .I1(\data_in_frame[18] [1]), .I2(\data_in_frame[19] [1]), .I3(byte_transmit_counter2[1]), 
            .O(n6303));
    defparam byte_transmit_counter2_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n6303_bdd_4_lut (.I0(n6303), .I1(data_in_field[137]), .I2(data_in_field[129]), 
            .I3(byte_transmit_counter2[1]), .O(n6306));
    defparam n6303_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2555_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[18] [0]), .I3(\data_in_frame[18] [0]), .O(n2806));
    defparam i2555_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2556_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[18] [1]), .I3(\data_in_frame[18] [1]), .O(n2807));
    defparam i2556_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2559_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[18] [4]), .I3(\data_in_frame[18] [4]), .O(n2810));
    defparam i2559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_925 (.I0(\data_in[3] [6]), .I1(n28_adj_1925), 
            .I2(n22_adj_1924), .I3(\data_in[2] [1]), .O(n30_adj_1941));   // coms.v(197[12:70])
    defparam i14_4_lut_adj_925.LUT_INIT = 16'hfffe;
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(CLK_c), .D(n2508));   // coms.v(174[10] 182[6])
    SB_LUT4 data_in_field_143__I_0_1808_2_lut (.I0(data_in_field[143]), .I1(data_in_field[142]), 
            .I2(GND_net), .I3(GND_net), .O(tx2_transmit_N_1031));   // coms.v(94[18:141])
    defparam data_in_field_143__I_0_1808_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_926 (.I0(data_in_field[86]), .I1(data_in_field[30]), 
            .I2(GND_net), .I3(GND_net), .O(n1917));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(CLK_c), .D(n2507));   // coms.v(174[10] 182[6])
    SB_LUT4 i2545_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[16] [6]), .I3(data_in_field[134]), .O(n2796));
    defparam i2545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(CLK_c), .D(n2506));   // coms.v(174[10] 182[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(CLK_c), .D(n2505));   // coms.v(174[10] 182[6])
    SB_LUT4 i2560_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[18] [5]), .I3(\data_in_frame[18] [5]), .O(n2811));
    defparam i2560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5903 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_in_frame[18] [2]), .I2(\data_in_frame[19] [2]), .I3(byte_transmit_counter2[1]), 
            .O(n6297));
    defparam byte_transmit_counter2_0__bdd_4_lut_5903.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_927 (.I0(data_in_field[29]), .I1(tx2_transmit_N_1031), 
            .I2(data_in_field[85]), .I3(data_in_field[141]), .O(n2030));   // coms.v(202[14:57])
    defparam i3_4_lut_adj_927.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_928 (.I0(data_in_field[60]), .I1(data_in_field[0]), 
            .I2(GND_net), .I3(GND_net), .O(n5590));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_928.LUT_INIT = 16'h6666;
    SB_LUT4 n6297_bdd_4_lut (.I0(n6297), .I1(data_in_field[138]), .I2(data_in_field[130]), 
            .I3(byte_transmit_counter2[1]), .O(n6300));
    defparam n6297_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2541_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[16] [2]), .I3(data_in_field[130]), .O(n2792));
    defparam i2541_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY data_527_add_4_4 (.CI(n4740), .I0(GND_net), .I1(data[2]), 
            .CO(n4741));
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(CLK_c), .D(n2504));   // coms.v(174[10] 182[6])
    SB_DFF data_out_0___i17 (.Q(\data_out[18] [0]), .C(CLK_c), .D(n2852));   // coms.v(123[10] 164[6])
    SB_LUT4 i2414_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[0] [3]), .I3(data_in_field[3]), .O(n2665));
    defparam i2414_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2413_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[0] [2]), .I3(data_in_field[2]), .O(n2664));
    defparam i2413_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_929 (.I0(data_in_field[124]), .I1(data_in_field[102]), 
            .I2(GND_net), .I3(GND_net), .O(n2026));   // coms.v(93[18:87])
    defparam i1_2_lut_adj_929.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_930 (.I0(\data_out[10] [5]), .I1(\data_out[10] [7]), 
            .I2(\data_out[11] [1]), .I3(\data_out[10] [6]), .O(n5440));   // coms.v(81[17:257])
    defparam i1_2_lut_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i2411_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[0] [1]), .I3(data_in_field[1]), .O(n2662));
    defparam i2411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2524_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[14] [1]), .I3(data_in_field[113]), .O(n2775));
    defparam i2524_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_1824_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n4707), .O(tx_transmit_N_568[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1824_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(CLK_c), .D(n2492));   // coms.v(174[10] 182[6])
    SB_DFF tx_transmit_1794 (.Q(tx_transmit), .C(CLK_c), .D(n4813));   // coms.v(123[10] 164[6])
    SB_DFF data_out_0___i18 (.Q(\data_out[18] [1]), .C(CLK_c), .D(n2853));   // coms.v(123[10] 164[6])
    SB_LUT4 i1_2_lut_3_lut_adj_931 (.I0(\data_out[11] [5]), .I1(\data_out[11] [4]), 
            .I2(n5409), .I3(GND_net), .O(n4_adj_5));
    defparam i1_2_lut_3_lut_adj_931.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_932 (.I0(data_in_field[94]), .I1(data_in_field[36]), 
            .I2(GND_net), .I3(GND_net), .O(n2009));   // coms.v(89[18:383])
    defparam i1_2_lut_adj_932.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_933 (.I0(\data_out[11] [4]), .I1(\data_out[11] [7]), 
            .I2(\data_out[11] [5]), .I3(\data_out[11] [6]), .O(n5479));
    defparam i1_2_lut_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_LUT4 i2530_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[14] [7]), .I3(data_in_field[119]), .O(n2781));
    defparam i2530_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2529_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[14] [6]), .I3(data_in_field[118]), .O(n2780));
    defparam i2529_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY delay_counter_528_add_4_3 (.CI(n4754), .I0(GND_net), .I1(delay_counter[1]), 
            .CO(n4755));
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(CLK_c), 
           .D(n2818));   // coms.v(192[10] 220[6])
    SB_LUT4 i2528_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[14] [5]), .I3(data_in_field[117]), .O(n2779));
    defparam i2528_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF byte_transmit_counter__i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
           .D(n2489));   // coms.v(123[10] 164[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(CLK_c), 
           .D(n2820));   // coms.v(192[10] 220[6])
    SB_LUT4 data_527_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(data[1]), 
            .I3(n4739), .O(n69[1])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_528_add_4_2_lut (.I0(GND_net), .I1(n4333), .I2(delay_counter[0]), 
            .I3(GND_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_528_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_528_add_4_2 (.CI(GND_net), .I0(n4333), .I1(delay_counter[0]), 
            .CO(n4754));
    SB_LUT4 data_527_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(data[15]), 
            .I3(n4753), .O(n69[15])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 data_527_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(data[14]), 
            .I3(n4752), .O(n69[14])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY data_527_add_4_16 (.CI(n4752), .I0(GND_net), .I1(data[14]), 
            .CO(n4753));
    SB_LUT4 data_527_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(data[13]), 
            .I3(n4751), .O(n69[13])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY data_527_add_4_15 (.CI(n4751), .I0(GND_net), .I1(data[13]), 
            .CO(n4752));
    SB_LUT4 i1_2_lut_adj_934 (.I0(data_in_field[51]), .I1(data_in_field[9]), 
            .I2(GND_net), .I3(GND_net), .O(n5369));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_935 (.I0(data_in_field[32]), .I1(data_in_field[33]), 
            .I2(data_in_field[54]), .I3(n5369), .O(n2125));   // coms.v(202[14:57])
    defparam i3_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5898 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_in_frame[18] [3]), .I2(\data_in_frame[19] [3]), .I3(byte_transmit_counter2[1]), 
            .O(n6279));
    defparam byte_transmit_counter2_0__bdd_4_lut_5898.LUT_INIT = 16'he4aa;
    SB_CARRY data_527_add_4_3 (.CI(n4739), .I0(GND_net), .I1(data[1]), 
            .CO(n4740));
    SB_LUT4 i2527_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[14] [4]), .I3(data_in_field[116]), .O(n2778));
    defparam i2527_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(CLK_c), 
           .D(n2817));   // coms.v(192[10] 220[6])
    SB_LUT4 i1_2_lut_adj_936 (.I0(data_in_field[38]), .I1(data_in_field[21]), 
            .I2(GND_net), .I3(GND_net), .O(n2062));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_936.LUT_INIT = 16'h6666;
    SB_LUT4 n6279_bdd_4_lut (.I0(n6279), .I1(data_in_field[139]), .I2(data_in_field[131]), 
            .I3(byte_transmit_counter2[1]), .O(n6282));
    defparam n6279_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_937 (.I0(\data_out[11] [7]), .I1(\data_out[11] [5]), 
            .I2(\data_out[11] [6]), .I3(GND_net), .O(n1579));
    defparam i1_2_lut_3_lut_adj_937.LUT_INIT = 16'h9696;
    SB_LUT4 data_527_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(data[12]), 
            .I3(n4750), .O(n69[12])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY data_527_add_4_14 (.CI(n4750), .I0(GND_net), .I1(data[12]), 
            .CO(n4751));
    SB_LUT4 i2_3_lut_adj_938 (.I0(data_in_field[78]), .I1(data_in_field[18]), 
            .I2(data_in_field[76]), .I3(GND_net), .O(n5388));   // coms.v(202[14:57])
    defparam i2_3_lut_adj_938.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5884 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[119]), .I2(data_in_field[127]), .I3(byte_transmit_counter2[1]), 
            .O(n6273));
    defparam byte_transmit_counter2_0__bdd_4_lut_5884.LUT_INIT = 16'he4aa;
    SB_LUT4 i2526_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[14] [3]), .I3(data_in_field[115]), .O(n2777));
    defparam i2526_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2525_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[14] [2]), .I3(data_in_field[114]), .O(n2776));
    defparam i2525_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2531_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[15] [0]), .I3(data_in_field[120]), .O(n2782));
    defparam i2531_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n6027_bdd_4_lut (.I0(n6027), .I1(data_in_field[72]), .I2(data_in_field[64]), 
            .I3(byte_transmit_counter2[1]), .O(n5794));
    defparam n6027_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR byte_transmit_counter2_525_526__i1 (.Q(byte_transmit_counter2[0]), 
            .C(CLK_c), .E(n195), .D(n2[0]), .R(n2325));   // coms.v(212[39:65])
    SB_CARRY add_1824_7 (.CI(n4707), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n4708));
    SB_LUT4 i2553_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[17] [6]), .I3(data_in_field[142]), .O(n2804));
    defparam i2553_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n6273_bdd_4_lut (.I0(n6273), .I1(data_in_field[111]), .I2(data_in_field[103]), 
            .I3(byte_transmit_counter2[1]), .O(n5686));
    defparam n6273_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF byte_transmit_counter__i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
           .D(n2875));   // coms.v(123[10] 164[6])
    SB_LUT4 data_527_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(data[0]), 
            .I3(VCC_net), .O(n69[0])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR byte_transmit_counter2_525_526__i2 (.Q(byte_transmit_counter2[1]), 
            .C(CLK_c), .E(n195), .D(n2[1]), .R(n2325));   // coms.v(212[39:65])
    SB_DFFESR byte_transmit_counter2_525_526__i3 (.Q(byte_transmit_counter2[2]), 
            .C(CLK_c), .E(n195), .D(n2[2]), .R(n2325));   // coms.v(212[39:65])
    SB_LUT4 i2_3_lut_adj_939 (.I0(data_in_field[59]), .I1(data_in_field[123]), 
            .I2(data_in_field[3]), .I3(GND_net), .O(n1979));   // coms.v(83[17:391])
    defparam i2_3_lut_adj_939.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5879 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_in_frame[18] [4]), .I2(\data_in_frame[19] [4]), .I3(byte_transmit_counter2[1]), 
            .O(n6267));
    defparam byte_transmit_counter2_0__bdd_4_lut_5879.LUT_INIT = 16'he4aa;
    SB_LUT4 i2549_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[17] [2]), .I3(data_in_field[138]), .O(n2800));
    defparam i2549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY data_527_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(data[0]), 
            .CO(n4739));
    SB_LUT4 add_1824_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n4706), .O(tx_transmit_N_568[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1824_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n6267_bdd_4_lut (.I0(n6267), .I1(data_in_field[140]), .I2(data_in_field[132]), 
            .I3(byte_transmit_counter2[1]), .O(n6270));
    defparam n6267_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_940 (.I0(data_in_field[138]), .I1(data_in_field[130]), 
            .I2(GND_net), .I3(GND_net), .O(n2056));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut (.I0(byte_transmit_counter2[2]), 
            .I1(n5994), .I2(n5686), .I3(byte_transmit_counter2[3]), .O(n6261));
    defparam byte_transmit_counter2_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter2_525_526_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[4]), .I3(n4738), .O(n2[4])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_525_526_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n6261_bdd_4_lut (.I0(n6261), .I1(n6000), .I2(n6012), .I3(byte_transmit_counter2[3]), 
            .O(n6264));
    defparam n6261_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2536_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[15] [5]), .I3(data_in_field[125]), .O(n2787));
    defparam i2536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut (.I0(data_in_field[41]), .I1(data_in_field[12]), 
            .I2(data_in_field[124]), .I3(data_in_field[102]), .O(n2101));   // coms.v(92[18:361])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_941 (.I0(data_in_field[31]), .I1(data_in_field[136]), 
            .I2(GND_net), .I3(GND_net), .O(n2113));   // coms.v(83[17:391])
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5874 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[22]), .I2(data_in_field[30]), .I3(byte_transmit_counter2[1]), 
            .O(n6255));
    defparam byte_transmit_counter2_0__bdd_4_lut_5874.LUT_INIT = 16'he4aa;
    SB_LUT4 i2535_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[15] [4]), .I3(data_in_field[124]), .O(n2786));
    defparam i2535_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n6255_bdd_4_lut (.I0(n6255), .I1(data_in_field[14]), .I2(data_in_field[6]), 
            .I3(byte_transmit_counter2[1]), .O(n5692));
    defparam n6255_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2534_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[15] [3]), .I3(data_in_field[123]), .O(n2785));
    defparam i2534_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2533_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[15] [2]), .I3(data_in_field[122]), .O(n2784));
    defparam i2533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5675 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[112]), .I2(data_in_field[120]), .I3(byte_transmit_counter2[1]), 
            .O(n6021));
    defparam byte_transmit_counter2_0__bdd_4_lut_5675.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_942 (.I0(data_in_field[72]), .I1(data_in_field[16]), 
            .I2(GND_net), .I3(GND_net), .O(n2089));   // coms.v(83[17:391])
    defparam i1_2_lut_adj_942.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_943 (.I0(data_in_field[50]), .I1(data_in_field[46]), 
            .I2(GND_net), .I3(GND_net), .O(n2077));   // coms.v(93[18:87])
    defparam i1_2_lut_adj_943.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5864 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[54]), .I2(data_in_field[62]), .I3(byte_transmit_counter2[1]), 
            .O(n6249));
    defparam byte_transmit_counter2_0__bdd_4_lut_5864.LUT_INIT = 16'he4aa;
    SB_LUT4 i2532_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[15] [1]), .I3(data_in_field[121]), .O(n2783));
    defparam i2532_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n6249_bdd_4_lut (.I0(n6249), .I1(data_in_field[46]), .I2(data_in_field[38]), 
            .I3(byte_transmit_counter2[1]), .O(n5695));
    defparam n6249_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_944 (.I0(data_in_field[64]), .I1(data_in_field[125]), 
            .I2(data_in_field[35]), .I3(GND_net), .O(n1913));   // coms.v(93[18:87])
    defparam i1_2_lut_3_lut_adj_944.LUT_INIT = 16'h9696;
    SB_LUT4 n6021_bdd_4_lut (.I0(n6021), .I1(data_in_field[104]), .I2(data_in_field[96]), 
            .I3(byte_transmit_counter2[1]), .O(n5797));
    defparam n6021_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5859 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[86]), .I2(data_in_field[94]), .I3(byte_transmit_counter2[1]), 
            .O(n6243));
    defparam byte_transmit_counter2_0__bdd_4_lut_5859.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_945 (.I0(data_in_field[95]), .I1(data_in_field[80]), 
            .I2(data_in_field[138]), .I3(data_in_field[130]), .O(n1835));   // coms.v(202[14:57])
    defparam i1_2_lut_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 n6243_bdd_4_lut (.I0(n6243), .I1(data_in_field[78]), .I2(data_in_field[70]), 
            .I3(byte_transmit_counter2[1]), .O(n5698));
    defparam n6243_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_946 (.I0(data_in_field[77]), .I1(data_in_field[135]), 
            .I2(data_in_field[92]), .I3(n1908), .O(n1973));   // coms.v(202[14:57])
    defparam i1_2_lut_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_947 (.I0(data_in_field[133]), .I1(data_in_field[143]), 
            .I2(data_in_field[38]), .I3(data_in_field[21]), .O(n5378));   // coms.v(202[14:57])
    defparam i2_3_lut_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i2538_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[15] [7]), .I3(data_in_field[127]), .O(n2789));
    defparam i2538_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_948 (.I0(n1958), .I1(n2056), .I2(n1979), .I3(n6_adj_1939), 
            .O(n5506));   // coms.v(83[17:391])
    defparam i4_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5661 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[55]), .I2(data_in_field[63]), .I3(byte_transmit_counter2[1]), 
            .O(n5997));
    defparam byte_transmit_counter2_0__bdd_4_lut_5661.LUT_INIT = 16'he4aa;
    SB_LUT4 i2537_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[15] [6]), .I3(data_in_field[126]), .O(n2788));
    defparam i2537_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n5997_bdd_4_lut (.I0(n5997), .I1(data_in_field[47]), .I2(data_in_field[39]), 
            .I3(byte_transmit_counter2[1]), .O(n6000));
    defparam n5997_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_949 (.I0(data_in_field[98]), .I1(data_in_field[100]), 
            .I2(GND_net), .I3(GND_net), .O(n5394));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5854 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[118]), .I2(data_in_field[126]), .I3(byte_transmit_counter2[1]), 
            .O(n6237));
    defparam byte_transmit_counter2_0__bdd_4_lut_5854.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_950 (.I0(tx_transmit_N_568[4]), .I1(n81_adj_1872), 
            .I2(n15), .I3(tx_transmit_N_568[2]), .O(n2870));   // coms.v(135[5:24])
    defparam i1_2_lut_4_lut_adj_950.LUT_INIT = 16'hcd00;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5670 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[23]), .I2(data_in_field[31]), .I3(byte_transmit_counter2[1]), 
            .O(n6009));
    defparam byte_transmit_counter2_0__bdd_4_lut_5670.LUT_INIT = 16'he4aa;
    SB_LUT4 n6237_bdd_4_lut (.I0(n6237), .I1(data_in_field[110]), .I2(data_in_field[102]), 
            .I3(byte_transmit_counter2[1]), .O(n5701));
    defparam n6237_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_951 (.I0(data_in_field[90]), .I1(data_in_field[89]), 
            .I2(GND_net), .I3(GND_net), .O(n1866));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_5869 (.I0(byte_transmit_counter2[2]), 
            .I1(n5698), .I2(n5701), .I3(byte_transmit_counter2[3]), .O(n6231));
    defparam byte_transmit_counter2_2__bdd_4_lut_5869.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5652 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[87]), .I2(data_in_field[95]), .I3(byte_transmit_counter2[1]), 
            .O(n5991));
    defparam byte_transmit_counter2_0__bdd_4_lut_5652.LUT_INIT = 16'he4aa;
    SB_CARRY add_1824_4 (.CI(n4704), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n4705));
    SB_LUT4 n6231_bdd_4_lut (.I0(n6231), .I1(n5695), .I2(n5692), .I3(byte_transmit_counter2[3]), 
            .O(n6234));
    defparam n6231_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_952 (.I0(data_in_field[109]), .I1(data_in_field[45]), 
            .I2(GND_net), .I3(GND_net), .O(n2149));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_5699 (.I0(byte_transmit_counter2[2]), 
            .I1(n5794), .I2(n5797), .I3(byte_transmit_counter2[3]), .O(n6015));
    defparam byte_transmit_counter2_2__bdd_4_lut_5699.LUT_INIT = 16'he4aa;
    SB_DFFESR byte_transmit_counter2_525_526__i4 (.Q(byte_transmit_counter2[3]), 
            .C(CLK_c), .E(n195), .D(n2[3]), .R(n2325));   // coms.v(212[39:65])
    SB_LUT4 byte_transmit_counter2_525_526_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[3]), .I3(n4737), .O(n2[3])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_525_526_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5849 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_in_frame[18] [5]), .I2(\data_in_frame[19] [5]), .I3(byte_transmit_counter2[1]), 
            .O(n6225));
    defparam byte_transmit_counter2_0__bdd_4_lut_5849.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_953 (.I0(data_in_field[68]), .I1(data_in_field[8]), 
            .I2(GND_net), .I3(GND_net), .O(n2039));   // coms.v(89[18:383])
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 n6225_bdd_4_lut (.I0(n6225), .I1(data_in_field[141]), .I2(data_in_field[133]), 
            .I3(byte_transmit_counter2[1]), .O(n6228));
    defparam n6225_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_954 (.I0(data_in_field[23]), .I1(data_in_field[7]), 
            .I2(data_in_field[53]), .I3(n2039), .O(n5458));   // coms.v(202[14:57])
    defparam i3_4_lut_adj_954.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5839 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[21]), .I2(data_in_field[29]), .I3(byte_transmit_counter2[1]), 
            .O(n6219));
    defparam byte_transmit_counter2_0__bdd_4_lut_5839.LUT_INIT = 16'he4aa;
    SB_LUT4 n5991_bdd_4_lut (.I0(n5991), .I1(data_in_field[79]), .I2(data_in_field[71]), 
            .I3(byte_transmit_counter2[1]), .O(n5994));
    defparam n5991_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n6219_bdd_4_lut (.I0(n6219), .I1(data_in_field[13]), .I2(data_in_field[5]), 
            .I3(byte_transmit_counter2[1]), .O(n5707));
    defparam n6219_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_955 (.I0(data_in_field[105]), .I1(n5458), .I2(GND_net), 
            .I3(GND_net), .O(n1994));   // coms.v(202[14:57])
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut_adj_956 (.I0(n25_adj_1929), .I1(n27_adj_1928), .I2(n26), 
            .I3(n28_adj_1926), .O(n4795));
    defparam i15_4_lut_adj_956.LUT_INIT = 16'h8000;
    SB_LUT4 i9_4_lut_adj_957 (.I0(\data_in[3] [2]), .I1(\data_in[2] [4]), 
            .I2(\data_in[3] [3]), .I3(\data_in[0] [0]), .O(n25_adj_1948));   // coms.v(197[12:70])
    defparam i9_4_lut_adj_957.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_958 (.I0(n25_adj_1948), .I1(n4795), .I2(n30_adj_1941), 
            .I3(n26_adj_1940), .O(n1729));   // coms.v(197[12:70])
    defparam i1_4_lut_adj_958.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_959 (.I0(\data_out[10] [2]), .I1(\data_out[10] [6]), 
            .I2(\data_out[11] [0]), .I3(GND_net), .O(n4_adj_6));
    defparam i1_2_lut_3_lut_adj_959.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_960 (.I0(data_in_field[47]), .I1(data_in_field[61]), 
            .I2(data_in_field[62]), .I3(GND_net), .O(n5551));   // coms.v(82[17:399])
    defparam i1_2_lut_3_lut_adj_960.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_961 (.I0(data_in_field[137]), .I1(data_in_field[25]), 
            .I2(data_in_field[39]), .I3(data_in_field[55]), .O(n5515));   // coms.v(92[18:361])
    defparam i1_2_lut_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_962 (.I0(data_in_field[34]), .I1(data_in_field[139]), 
            .I2(data_in_field[19]), .I3(data_in_field[77]), .O(n2092));   // coms.v(202[14:57])
    defparam i1_2_lut_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out[10] [2]), .I1(\data_out[10] [6]), 
            .I2(\data_out[10] [3]), .I3(GND_net), .O(n7));   // coms.v(85[17:241])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_963 (.I0(\data_out[10] [0]), .I1(\data_out[11] [3]), 
            .I2(\data_out[11] [2]), .I3(n5421), .O(n5400));   // coms.v(85[17:241])
    defparam i1_2_lut_4_lut_adj_963.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_964 (.I0(data_in_field[101]), .I1(data_in_field[13]), 
            .I2(data_in_field[69]), .I3(data_in_field[110]), .O(n6_adj_1918));   // coms.v(93[18:87])
    defparam i1_2_lut_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_965 (.I0(data_in_field[137]), .I1(data_in_field[25]), 
            .I2(data_in_field[39]), .I3(data_in_field[71]), .O(n5542));   // coms.v(92[18:361])
    defparam i1_2_lut_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_966 (.I0(data_in_field[65]), .I1(data_in_field[5]), 
            .I2(n10_adj_1915), .I3(data_in_field[21]), .O(n5521));   // coms.v(86[17:391])
    defparam i5_3_lut_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 i1047_2_lut (.I0(byte_transmit_counter2[2]), .I1(byte_transmit_counter2[3]), 
            .I2(GND_net), .I3(GND_net), .O(n1081));   // coms.v(189[35:57])
    defparam i1047_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5622_4_lut (.I0(byte_transmit_counter2[0]), .I1(byte_transmit_counter2[4]), 
            .I2(n1081), .I3(byte_transmit_counter2[1]), .O(\FRAME_MATCHER.wait_for_transmission_N_909 ));
    defparam i5622_4_lut.LUT_INIT = 16'h373f;
    SB_LUT4 i1_2_lut_3_lut_adj_967 (.I0(data_in_field[65]), .I1(data_in_field[5]), 
            .I2(data_in_field[4]), .I3(GND_net), .O(n2104));   // coms.v(86[17:391])
    defparam i1_2_lut_3_lut_adj_967.LUT_INIT = 16'h9696;
    SB_LUT4 i746_2_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n1253));   // coms.v(39[29:50])
    defparam i746_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i951_2_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n1251));   // coms.v(39[29:50])
    defparam i951_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out[18] [7]), 
            .I1(\data_out[19] [7]), .I2(byte_transmit_counter[0]), .I3(GND_net), 
            .O(n17_adj_1950));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5563_3_lut (.I0(n17_adj_1950), .I1(n1251), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n5827));   // coms.v(39[29:50])
    defparam i5563_3_lut.LUT_INIT = 16'h2323;
    SB_LUT4 i1006_4_lut (.I0(byte_transmit_counter[0]), .I1(\data_out[10] [7]), 
            .I2(byte_transmit_counter[3]), .I3(\data_out[11] [7]), .O(n1249));   // coms.v(39[29:50])
    defparam i1006_4_lut.LUT_INIT = 16'he545;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_4_lut (.I0(n1249), .I1(n5827), 
            .I2(byte_transmit_counter[4]), .I3(n1253), .O(i_Tx_Byte[7]));   // coms.v(39[29:50])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_4_lut.LUT_INIT = 16'hcacf;
    SB_LUT4 i1_2_lut_3_lut_adj_968 (.I0(\data_out[10] [7]), .I1(\data_out[11] [1]), 
            .I2(\data_out[10] [6]), .I3(GND_net), .O(n5448));   // coms.v(81[17:257])
    defparam i1_2_lut_3_lut_adj_968.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5834 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[53]), .I2(data_in_field[61]), .I3(byte_transmit_counter2[1]), 
            .O(n6213));
    defparam byte_transmit_counter2_0__bdd_4_lut_5834.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_969 (.I0(data_in_field[120]), .I1(data_in_field[128]), 
            .I2(data_in_field[98]), .I3(GND_net), .O(n2107));   // coms.v(89[18:383])
    defparam i2_3_lut_adj_969.LUT_INIT = 16'h9696;
    SB_LUT4 n6213_bdd_4_lut (.I0(n6213), .I1(data_in_field[45]), .I2(data_in_field[37]), 
            .I3(byte_transmit_counter2[1]), .O(n5710));
    defparam n6213_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_970 (.I0(n1973), .I1(n1892), .I2(n1942), .I3(n2095), 
            .O(n12_adj_1951));   // coms.v(202[14:57])
    defparam i5_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_971 (.I0(data_in_field[20]), .I1(data_in_field[34]), 
            .I2(data_in_field[132]), .I3(n2143), .O(n5557));   // coms.v(202[14:57])
    defparam i1_2_lut_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5829 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[85]), .I2(data_in_field[93]), .I3(byte_transmit_counter2[1]), 
            .O(n6207));
    defparam byte_transmit_counter2_0__bdd_4_lut_5829.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_972 (.I0(n2107), .I1(n12_adj_1951), .I2(n1994), 
            .I3(data_in_field[37]), .O(n5488));   // coms.v(202[14:57])
    defparam i6_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 n6207_bdd_4_lut (.I0(n6207), .I1(data_in_field[77]), .I2(data_in_field[69]), 
            .I3(byte_transmit_counter2[1]), .O(n5713));
    defparam n6207_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_973 (.I0(data_in_field[48]), .I1(data_in_field[63]), 
            .I2(data_in_field[62]), .I3(data_in_field[90]), .O(n5443));   // coms.v(83[17:391])
    defparam i1_2_lut_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_974 (.I0(data_in_field[48]), .I1(data_in_field[63]), 
            .I2(data_in_field[62]), .I3(n5593), .O(n5430));   // coms.v(83[17:391])
    defparam i1_2_lut_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_975 (.I0(\data_out[11] [3]), .I1(\data_out[11] [2]), 
            .I2(n5421), .I3(GND_net), .O(n135));   // coms.v(79[17:447])
    defparam i1_2_lut_3_lut_adj_975.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5824 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[117]), .I2(data_in_field[125]), .I3(byte_transmit_counter2[1]), 
            .O(n6201));
    defparam byte_transmit_counter2_0__bdd_4_lut_5824.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_976 (.I0(n2000), .I1(n2056), .I2(n2074), 
            .I3(data_in_field[41]), .O(n5527));   // coms.v(202[14:57])
    defparam i2_3_lut_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 i3445_2_lut (.I0(tx2_active), .I1(r_SM_Main_2__N_1770[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3689));
    defparam i3445_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 n6201_bdd_4_lut (.I0(n6201), .I1(data_in_field[109]), .I2(data_in_field[101]), 
            .I3(byte_transmit_counter2[1]), .O(n5716));
    defparam n6201_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15_4_lut_adj_977 (.I0(data_in_field[80]), .I1(data_in_field[48]), 
            .I2(data_in_field[70]), .I3(\data_in[18] [7]), .O(n42));   // coms.v(202[14:57])
    defparam i15_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_5844 (.I0(byte_transmit_counter2[2]), 
            .I1(n5713), .I2(n5716), .I3(byte_transmit_counter2[3]), .O(n6195));
    defparam byte_transmit_counter2_2__bdd_4_lut_5844.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_978 (.I0(\data_out[11] [3]), .I1(\data_out[11] [2]), 
            .I2(\data_out[11] [0]), .I3(GND_net), .O(n5409));   // coms.v(79[17:447])
    defparam i1_2_lut_3_lut_adj_978.LUT_INIT = 16'h9696;
    SB_LUT4 n6195_bdd_4_lut (.I0(n6195), .I1(n5710), .I2(n5707), .I3(byte_transmit_counter2[3]), 
            .O(n6198));
    defparam n6195_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i19_4_lut_adj_979 (.I0(n5506), .I1(n5533), .I2(n6414), .I3(n5542), 
            .O(n46));   // coms.v(202[14:57])
    defparam i19_4_lut_adj_979.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter2_525_526__i5 (.Q(byte_transmit_counter2[4]), 
            .C(CLK_c), .E(n195), .D(n2[4]), .R(n2325));   // coms.v(212[39:65])
    SB_LUT4 add_1824_3_lut (.I0(n4334), .I1(byte_transmit_counter[1]), .I2(GND_net), 
            .I3(n4703), .O(n2869)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1824_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 data_527_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(data[11]), 
            .I3(n4749), .O(n69[11])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY byte_transmit_counter2_525_526_add_4_5 (.CI(n4737), .I0(GND_net), 
            .I1(byte_transmit_counter2[3]), .CO(n4738));
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5819 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[20]), .I2(data_in_field[28]), .I3(byte_transmit_counter2[1]), 
            .O(n6189));
    defparam byte_transmit_counter2_0__bdd_4_lut_5819.LUT_INIT = 16'he4aa;
    SB_LUT4 i17_4_lut (.I0(n2062), .I1(n2125), .I2(data_in_field[126]), 
            .I3(n5436), .O(n44));   // coms.v(202[14:57])
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(data_in_field[12]), .I1(n36), .I2(n5466), .I3(n2026), 
            .O(n45));   // coms.v(202[14:57])
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_525_526_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[2]), .I3(n4736), .O(n2[2])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_525_526_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY data_527_add_4_13 (.CI(n4749), .I0(GND_net), .I1(data[11]), 
            .CO(n4750));
    SB_LUT4 i2_3_lut_4_lut_adj_980 (.I0(data_in_field[131]), .I1(data_in_field[11]), 
            .I2(data_in_field[123]), .I3(data_in_field[67]), .O(n1926));   // coms.v(92[18:361])
    defparam i2_3_lut_4_lut_adj_980.LUT_INIT = 16'h6996;
    SB_LUT4 i9_2_lut_3_lut (.I0(data_in_field[131]), .I1(data_in_field[11]), 
            .I2(n5488), .I3(GND_net), .O(n36));   // coms.v(92[18:361])
    defparam i9_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_981 (.I0(\data_out[11] [3]), .I1(n5479), 
            .I2(\data_out[10] [7]), .I3(GND_net), .O(n7_adj_7));
    defparam i2_2_lut_3_lut_adj_981.LUT_INIT = 16'h9696;
    SB_LUT4 n6189_bdd_4_lut (.I0(n6189), .I1(data_in_field[12]), .I2(data_in_field[4]), 
            .I3(byte_transmit_counter2[1]), .O(n5722));
    defparam n6189_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(CLK_c), 
           .D(n2816));   // coms.v(192[10] 220[6])
    SB_LUT4 i16_4_lut (.I0(n2155), .I1(n2104), .I2(data_in_field[82]), 
            .I3(n2080), .O(n43));   // coms.v(202[14:57])
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_982 (.I0(data_in_field[87]), .I1(data_in_field[128]), 
            .I2(data_in_field[143]), .I3(data_in_field[142]), .O(n5539));   // coms.v(83[17:391])
    defparam i1_2_lut_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5809 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[52]), .I2(data_in_field[60]), .I3(byte_transmit_counter2[1]), 
            .O(n6183));
    defparam byte_transmit_counter2_0__bdd_4_lut_5809.LUT_INIT = 16'he4aa;
    SB_LUT4 i7_3_lut_adj_983 (.I0(data_in_field[107]), .I1(n5515), .I2(data_in_field[121]), 
            .I3(GND_net), .O(n24_adj_1877));   // coms.v(202[14:57])
    defparam i7_3_lut_adj_983.LUT_INIT = 16'h9696;
    SB_LUT4 i13_4_lut_adj_984 (.I0(n5545), .I1(n5578), .I2(n5569), .I3(n18_adj_1938), 
            .O(n30));   // coms.v(202[14:57])
    defparam i13_4_lut_adj_984.LUT_INIT = 16'h6996;
    SB_LUT4 n6183_bdd_4_lut (.I0(n6183), .I1(data_in_field[44]), .I2(data_in_field[36]), 
            .I3(byte_transmit_counter2[1]), .O(n5725));
    defparam n6183_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_985 (.I0(\data_in[19] [7]), .I1(data_in_field[36]), 
            .I2(data_in_field[131]), .I3(data_in_field[141]), .O(n22_adj_1886));   // coms.v(86[17:391])
    defparam i8_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 i2542_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[16] [3]), .I3(data_in_field[131]), .O(n2793));
    defparam i2542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_986 (.I0(n1779), .I1(n1889), .I2(n1948), .I3(data_in_field[108]), 
            .O(n18_adj_1887));   // coms.v(202[14:57])
    defparam i7_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5804 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[84]), .I2(data_in_field[92]), .I3(byte_transmit_counter2[1]), 
            .O(n6177));
    defparam byte_transmit_counter2_0__bdd_4_lut_5804.LUT_INIT = 16'he4aa;
    SB_LUT4 n6177_bdd_4_lut (.I0(n6177), .I1(data_in_field[76]), .I2(data_in_field[68]), 
            .I3(byte_transmit_counter2[1]), .O(n5728));
    defparam n6177_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_987 (.I0(\data_out[11] [3]), .I1(n5479), 
            .I2(\data_out[10] [0]), .I3(\data_out[11] [2]), .O(n5364));
    defparam i2_3_lut_4_lut_adj_987.LUT_INIT = 16'h6996;
    SB_LUT4 i2546_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[16] [7]), .I3(data_in_field[135]), .O(n2797));
    defparam i2546_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5799 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[116]), .I2(data_in_field[124]), .I3(byte_transmit_counter2[1]), 
            .O(n6171));
    defparam byte_transmit_counter2_0__bdd_4_lut_5799.LUT_INIT = 16'he4aa;
    SB_LUT4 n6171_bdd_4_lut (.I0(n6171), .I1(data_in_field[108]), .I2(data_in_field[100]), 
            .I3(byte_transmit_counter2[1]), .O(n5731));
    defparam n6171_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2550_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[17] [3]), .I3(data_in_field[139]), .O(n2801));
    defparam i2550_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut_adj_988 (.I0(n5418), .I1(n5491), .I2(n5443), .I3(n5509), 
            .O(n44_adj_1894));   // coms.v(202[14:57])
    defparam i18_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 i2554_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[17] [7]), .I3(data_in_field[143]), .O(n2805));
    defparam i2554_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2558_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[18] [3]), .I3(\data_in_frame[18] [3]), .O(n2809));
    defparam i2558_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2562_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[18] [7]), .I3(\data_in_frame[18] [7]), .O(n2813));
    defparam i2562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2563_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[19] [0]), .I3(\data_in_frame[19] [0]), .O(n2814));
    defparam i2563_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2564_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[19] [1]), .I3(\data_in_frame[19] [1]), .O(n2815));
    defparam i2564_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2565_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[19] [2]), .I3(\data_in_frame[19] [2]), .O(n2816));
    defparam i2565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter2_2__bdd_4_lut_5814 (.I0(byte_transmit_counter2[2]), 
            .I1(n5728), .I2(n5731), .I3(byte_transmit_counter2[3]), .O(n6165));
    defparam byte_transmit_counter2_2__bdd_4_lut_5814.LUT_INIT = 16'he4aa;
    SB_LUT4 i2566_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[19] [3]), .I3(\data_in_frame[19] [3]), .O(n2817));
    defparam i2566_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_989 (.I0(data_in_field[25]), .I1(data_in_field[120]), 
            .I2(n2089), .I3(n1994), .O(n41));   // coms.v(202[14:57])
    defparam i15_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 i4_3_lut (.I0(n5533), .I1(data_in_field[117]), .I2(n1855), 
            .I3(GND_net), .O(n12_adj_1898));   // coms.v(202[14:57])
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 n6165_bdd_4_lut (.I0(n6165), .I1(n5725), .I2(n5722), .I3(byte_transmit_counter2[3]), 
            .O(n6168));
    defparam n6165_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2569_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[19] [6]), .I3(\data_in_frame[19] [6]), .O(n2820));
    defparam i2569_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2567_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[19] [4]), .I3(\data_in_frame[19] [4]), .O(n2818));
    defparam i2567_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(CLK_c), 
           .D(n2815));   // coms.v(192[10] 220[6])
    SB_LUT4 i1_2_lut_3_lut_adj_990 (.I0(\data_out[10] [1]), .I1(\data_out[10] [3]), 
            .I2(\data_out[11] [3]), .I3(GND_net), .O(n4_adj_8));   // coms.v(79[17:447])
    defparam i1_2_lut_3_lut_adj_990.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out[10] [1]), .I1(\data_out[10] [3]), 
            .I2(\data_out[11] [0]), .I3(n5424), .O(n8_adj_9));   // coms.v(79[17:447])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2570_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[19] [7]), .I3(\data_in_frame[19] [7]), .O(n2821));
    defparam i2570_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2539_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[16] [0]), .I3(data_in_field[128]), .O(n2790));
    defparam i2539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2540_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[16] [1]), .I3(data_in_field[129]), .O(n2791));
    defparam i2540_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2543_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[16] [4]), .I3(data_in_field[132]), .O(n2794));
    defparam i2543_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_991 (.I0(\data_in[19] [6]), .I1(n2026), .I2(n1958), 
            .I3(n5391), .O(n13));   // coms.v(202[14:57])
    defparam i5_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i2544_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[16] [5]), .I3(data_in_field[133]), .O(n2795));
    defparam i2544_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_3_lut (.I0(n5458), .I1(n2155), .I2(data_in_field[73]), 
            .I3(GND_net), .O(n28_adj_1955));   // coms.v(82[17:399])
    defparam i8_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2523_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[14] [0]), .I3(data_in_field[112]), .O(n2774));
    defparam i2523_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2522_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[13] [7]), .I3(data_in_field[111]), .O(n2773));
    defparam i2522_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2521_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[13] [6]), .I3(data_in_field[110]), .O(n2772));
    defparam i2521_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2520_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[13] [5]), .I3(data_in_field[109]), .O(n2771));
    defparam i2520_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2519_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[13] [4]), .I3(data_in_field[108]), .O(n2770));
    defparam i2519_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(CLK_c), 
           .D(n2814));   // coms.v(192[10] 220[6])
    SB_LUT4 i13_4_lut_adj_992 (.I0(n2043), .I1(data_in_field[18]), .I2(data_in_field[107]), 
            .I3(n5372), .O(n33));   // coms.v(82[17:399])
    defparam i13_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5794 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[19]), .I2(data_in_field[27]), .I3(byte_transmit_counter2[1]), 
            .O(n6159));
    defparam byte_transmit_counter2_0__bdd_4_lut_5794.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_adj_993 (.I0(n1814), .I1(n2143), .I2(\data_in[19] [1]), 
            .I3(data_in_field[109]), .O(n32_adj_1901));   // coms.v(82[17:399])
    defparam i12_4_lut_adj_993.LUT_INIT = 16'h6996;
    SB_LUT4 n6159_bdd_4_lut (.I0(n6159), .I1(data_in_field[11]), .I2(data_in_field[3]), 
            .I3(byte_transmit_counter2[1]), .O(n5737));
    defparam n6159_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_994 (.I0(\data_out[10] [1]), .I1(\data_out[10] [3]), 
            .I2(\data_out[10] [5]), .I3(GND_net), .O(n5433));   // coms.v(79[17:447])
    defparam i1_2_lut_3_lut_adj_994.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_995 (.I0(\data_out[10] [0]), .I1(\data_out[10] [4]), 
            .I2(\data_out[11] [6]), .I3(\data_out[11] [7]), .O(n4_adj_10));
    defparam i1_2_lut_3_lut_4_lut_adj_995.LUT_INIT = 16'h6996;
    SB_LUT4 i2518_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[13] [3]), .I3(data_in_field[107]), .O(n2769));
    defparam i2518_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_996 (.I0(n2053), .I1(n2101), .I2(n2134), .I3(data_in_field[50]), 
            .O(n31_adj_1900));   // coms.v(82[17:399])
    defparam i11_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_DFF delay_counter_528__i6 (.Q(delay_counter[6]), .C(CLK_c), .D(n1[6]));   // coms.v(159[11] 161[5])
    SB_LUT4 i2_2_lut_3_lut_adj_997 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter[2]), .I3(GND_net), .O(n1508));   // coms.v(39[29:50])
    defparam i2_2_lut_3_lut_adj_997.LUT_INIT = 16'h0404;
    SB_CARRY byte_transmit_counter2_525_526_add_4_4 (.CI(n4736), .I0(GND_net), 
            .I1(byte_transmit_counter2[2]), .CO(n4737));
    SB_LUT4 i2517_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[13] [2]), .I3(data_in_field[106]), .O(n2768));
    defparam i2517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5784 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[51]), .I2(data_in_field[59]), .I3(byte_transmit_counter2[1]), 
            .O(n6153));
    defparam byte_transmit_counter2_0__bdd_4_lut_5784.LUT_INIT = 16'he4aa;
    SB_LUT4 i15_4_lut_adj_998 (.I0(n5497), .I1(n5548), .I2(n5515), .I3(n5581), 
            .O(n35));   // coms.v(82[17:399])
    defparam i15_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_999 (.I0(n33), .I1(n5378), .I2(n28_adj_1955), 
            .I3(n5430), .O(n37));   // coms.v(82[17:399])
    defparam i17_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 i2516_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[13] [1]), .I3(data_in_field[105]), .O(n2767));
    defparam i2516_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2515_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[13] [0]), .I3(data_in_field[104]), .O(n2766));
    defparam i2515_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1000 (.I0(\data_out[10] [0]), .I1(\data_out[10] [4]), 
            .I2(\data_out[10] [2]), .I3(GND_net), .O(n5424));
    defparam i1_2_lut_3_lut_adj_1000.LUT_INIT = 16'h9696;
    SB_LUT4 i2514_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[12] [7]), .I3(data_in_field[103]), .O(n2765));
    defparam i2514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2513_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[12] [6]), .I3(data_in_field[102]), .O(n2764));
    defparam i2513_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2512_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[12] [5]), .I3(data_in_field[101]), .O(n2763));
    defparam i2512_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2511_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[12] [4]), .I3(data_in_field[100]), .O(n2762));
    defparam i2511_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(CLK_c), 
           .D(n2813));   // coms.v(192[10] 220[6])
    SB_LUT4 i2_2_lut (.I0(data_in_field[57]), .I1(data_in_field[117]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_1957));   // coms.v(92[18:361])
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2510_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[12] [3]), .I3(data_in_field[99]), .O(n2761));
    defparam i2510_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n6015_bdd_4_lut (.I0(n6015), .I1(n5791), .I2(n5788), .I3(byte_transmit_counter2[3]), 
            .O(n6018));
    defparam n6015_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n6153_bdd_4_lut (.I0(n6153), .I1(data_in_field[43]), .I2(data_in_field[35]), 
            .I3(byte_transmit_counter2[1]), .O(n5740));
    defparam n6153_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_3_lut_4_lut_adj_1001 (.I0(data_in_field[88]), .I1(data_in_field[28]), 
            .I2(data_in_field[98]), .I3(data_in_field[121]), .O(n23_adj_1935));   // coms.v(202[14:57])
    defparam i8_3_lut_4_lut_adj_1001.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(CLK_c), 
           .D(n2809));   // coms.v(192[10] 220[6])
    SB_LUT4 i2509_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[12] [2]), .I3(data_in_field[98]), .O(n2760));
    defparam i2509_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2508_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[12] [1]), .I3(data_in_field[97]), .O(n2759));
    defparam i2508_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2507_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[12] [0]), .I3(data_in_field[96]), .O(n2758));
    defparam i2507_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i144 (.Q(data_in_field[143]), .C(CLK_c), .D(n2805));   // coms.v(192[10] 220[6])
    SB_LUT4 byte_transmit_counter2_525_526_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(byte_transmit_counter2[1]), .I3(n4735), .O(n2[1])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_525_526_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5779 (.I0(byte_transmit_counter2[0]), 
            .I1(\data_in_frame[18] [6]), .I2(\data_in_frame[19] [6]), .I3(byte_transmit_counter2[1]), 
            .O(n6147));
    defparam byte_transmit_counter2_0__bdd_4_lut_5779.LUT_INIT = 16'he4aa;
    SB_LUT4 i8_4_lut_adj_1002 (.I0(data_in_field[132]), .I1(data_in_field[109]), 
            .I2(data_in_field[139]), .I3(n5469), .O(n20_adj_1958));   // coms.v(92[18:361])
    defparam i8_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 n6147_bdd_4_lut (.I0(n6147), .I1(data_in_field[142]), .I2(data_in_field[134]), 
            .I3(byte_transmit_counter2[1]), .O(n6150));
    defparam n6147_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i140 (.Q(data_in_field[139]), .C(CLK_c), .D(n2801));   // coms.v(192[10] 220[6])
    SB_LUT4 i6_3_lut (.I0(n5578), .I1(data_in_field[101]), .I2(data_in_field[87]), 
            .I3(GND_net), .O(n18_adj_1904));   // coms.v(92[18:361])
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2506_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[11] [7]), .I3(data_in_field[95]), .O(n2757));
    defparam i2506_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY byte_transmit_counter2_525_526_add_4_3 (.CI(n4735), .I0(GND_net), 
            .I1(byte_transmit_counter2[1]), .CO(n4736));
    SB_LUT4 i7_3_lut_4_lut (.I0(data_in_field[88]), .I1(data_in_field[28]), 
            .I2(data_in_field[26]), .I3(data_in_field[58]), .O(n20_adj_1878));   // coms.v(202[14:57])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i136 (.Q(data_in_field[135]), .C(CLK_c), .D(n2797));   // coms.v(192[10] 220[6])
    SB_CARRY add_1824_6 (.CI(n4706), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n4707));
    SB_LUT4 i2505_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[11] [6]), .I3(data_in_field[94]), .O(n2756));
    defparam i2505_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2504_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[11] [5]), .I3(data_in_field[93]), .O(n2755));
    defparam i2504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i132 (.Q(data_in_field[131]), .C(CLK_c), .D(n2793));   // coms.v(192[10] 220[6])
    SB_LUT4 i2503_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[11] [4]), .I3(data_in_field[92]), .O(n2754));
    defparam i2503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2502_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[11] [3]), .I3(data_in_field[91]), .O(n2753));
    defparam i2502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2501_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[11] [2]), .I3(data_in_field[90]), .O(n2752));
    defparam i2501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1003 (.I0(data_in_field[53]), .I1(n20_adj_1958), 
            .I2(n14_adj_1957), .I3(\data_in[18] [5]), .O(n22_adj_1903));   // coms.v(92[18:361])
    defparam i10_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5774 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[83]), .I2(data_in_field[91]), .I3(byte_transmit_counter2[1]), 
            .O(n6141));
    defparam byte_transmit_counter2_0__bdd_4_lut_5774.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1004 (.I0(tx_transmit_N_568[4]), .I1(n81_adj_1872), 
            .I2(n15), .I3(tx_transmit_N_568[3]), .O(n2871));   // coms.v(135[5:24])
    defparam i1_2_lut_4_lut_adj_1004.LUT_INIT = 16'hcd00;
    SB_LUT4 n6141_bdd_4_lut (.I0(n6141), .I1(data_in_field[75]), .I2(data_in_field[67]), 
            .I3(byte_transmit_counter2[1]), .O(n5743));
    defparam n6141_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter2_525_526_add_4_2_lut (.I0(GND_net), .I1(\FRAME_MATCHER.wait_for_transmission_N_909 ), 
            .I2(byte_transmit_counter2[0]), .I3(GND_net), .O(n2[0])) /* synthesis syn_instantiated=1 */ ;
    defparam byte_transmit_counter2_525_526_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 data_527_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(data[10]), 
            .I3(n4748), .O(n69[10])) /* synthesis syn_instantiated=1 */ ;
    defparam data_527_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1824_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n4705), .O(tx_transmit_N_568[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1824_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2500_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[11] [1]), .I3(data_in_field[89]), .O(n2751));
    defparam i2500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2499_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[11] [0]), .I3(data_in_field[88]), .O(n2750));
    defparam i2499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2498_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[10] [7]), .I3(data_in_field[87]), .O(n2749));
    defparam i2498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2497_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[10] [6]), .I3(data_in_field[86]), .O(n2748));
    defparam i2497_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2496_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[10] [5]), .I3(data_in_field[85]), .O(n2747));
    defparam i2496_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2495_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[10] [4]), .I3(data_in_field[84]), .O(n2746));
    defparam i2495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2494_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[10] [3]), .I3(data_in_field[83]), .O(n2745));
    defparam i2494_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1005 (.I0(\data_out[11] [7]), .I1(\data_out[11] [6]), 
            .I2(\data_out[11] [5]), .I3(\data_out[11] [4]), .O(n5421));   // coms.v(91[18:225])
    defparam i2_3_lut_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i2493_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[10] [2]), .I3(data_in_field[82]), .O(n2744));
    defparam i2493_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1006 (.I0(data_in_field[87]), .I1(data_in_field[2]), 
            .I2(n1973), .I3(n2065), .O(n18_adj_1959));   // coms.v(82[17:399])
    defparam i7_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1007 (.I0(data_in_field[57]), .I1(n5551), .I2(data_in_field[113]), 
            .I3(GND_net), .O(n16));   // coms.v(82[17:399])
    defparam i5_3_lut_adj_1007.LUT_INIT = 16'h9696;
    SB_LUT4 i2492_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[10] [1]), .I3(data_in_field[81]), .O(n2743));
    defparam i2492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2491_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[10] [0]), .I3(data_in_field[80]), .O(n2742));
    defparam i2491_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2490_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[9] [7]), .I3(data_in_field[79]), .O(n2741));
    defparam i2490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2489_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[9] [6]), .I3(data_in_field[78]), .O(n2740));
    defparam i2489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1008 (.I0(n5575), .I1(n18_adj_1959), .I2(\data_in[19] [3]), 
            .I3(data_in_field[43]), .O(n20_adj_1870));   // coms.v(82[17:399])
    defparam i9_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_0__bdd_4_lut_5769 (.I0(byte_transmit_counter2[0]), 
            .I1(data_in_field[115]), .I2(data_in_field[123]), .I3(byte_transmit_counter2[1]), 
            .O(n6135));
    defparam byte_transmit_counter2_0__bdd_4_lut_5769.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(byte_transmit_counter[3]), .I2(n5853), .I3(byte_transmit_counter[2]), 
            .O(n6309));   // coms.v(39[29:50])
    defparam byte_transmit_counter_2__bdd_4_lut_4_lut.LUT_INIT = 16'h77c0;
    SB_LUT4 i5628_2_lut (.I0(\FRAME_MATCHER.wait_for_transmission ), .I1(n3703), 
            .I2(GND_net), .I3(GND_net), .O(n2325));
    defparam i5628_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2_3_lut_4_lut_adj_1009 (.I0(data_in_field[32]), .I1(data_in_field[88]), 
            .I2(data_in_field[58]), .I3(data_in_field[114]), .O(n5575));   // coms.v(83[17:391])
    defparam i2_3_lut_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_1_i31_4_lut (.I0(n6060), .I1(n6306), 
            .I2(byte_transmit_counter2[4]), .I3(n1081), .O(tx2_data[1]));   // coms.v(189[35:57])
    defparam byte_transmit_counter2_4__I_0_Mux_1_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i2_3_lut_4_lut_adj_1010 (.I0(data_in_field[32]), .I1(data_in_field[88]), 
            .I2(n1779), .I3(data_in_field[60]), .O(n5500));   // coms.v(83[17:391])
    defparam i2_3_lut_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_2_i31_4_lut (.I0(n6102), .I1(n6300), 
            .I2(byte_transmit_counter2[4]), .I3(n1081), .O(tx2_data[2]));   // coms.v(189[35:57])
    defparam byte_transmit_counter2_4__I_0_Mux_2_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_3_i31_4_lut (.I0(n6132), .I1(n6282), 
            .I2(byte_transmit_counter2[4]), .I3(n1081), .O(tx2_data[3]));   // coms.v(189[35:57])
    defparam byte_transmit_counter2_4__I_0_Mux_3_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_4_i31_4_lut (.I0(n6168), .I1(n6270), 
            .I2(byte_transmit_counter2[4]), .I3(n1081), .O(tx2_data[4]));   // coms.v(189[35:57])
    defparam byte_transmit_counter2_4__I_0_Mux_4_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_5_i31_4_lut (.I0(n6198), .I1(n6228), 
            .I2(byte_transmit_counter2[4]), .I3(n1081), .O(tx2_data[5]));   // coms.v(189[35:57])
    defparam byte_transmit_counter2_4__I_0_Mux_5_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_6_i31_4_lut (.I0(n6234), .I1(n6150), 
            .I2(byte_transmit_counter2[4]), .I3(n1081), .O(tx2_data[6]));   // coms.v(189[35:57])
    defparam byte_transmit_counter2_4__I_0_Mux_6_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter2_4__I_0_Mux_7_i31_4_lut (.I0(n6264), .I1(n6084), 
            .I2(byte_transmit_counter2[4]), .I3(n1081), .O(tx2_data[7]));   // coms.v(189[35:57])
    defparam byte_transmit_counter2_4__I_0_Mux_7_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i2488_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[9] [5]), .I3(data_in_field[77]), .O(n2739));
    defparam i2488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2487_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[9] [4]), .I3(data_in_field[76]), .O(n2738));
    defparam i2487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2486_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[9] [3]), .I3(data_in_field[75]), .O(n2737));
    defparam i2486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2485_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[9] [2]), .I3(data_in_field[74]), .O(n2736));
    defparam i2485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2484_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[9] [1]), .I3(data_in_field[73]), .O(n2735));
    defparam i2484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2483_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[9] [0]), .I3(data_in_field[72]), .O(n2734));
    defparam i2483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_3_lut_4_lut (.I0(data_in_field[124]), .I1(data_in_field[4]), 
            .I2(data_in_field[101]), .I3(data_in_field[87]), .O(n18));   // coms.v(202[14:57])
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2482_3_lut_4_lut (.I0(n1729), .I1(\FRAME_MATCHER.wait_for_transmission ), 
            .I2(\data_in[8] [7]), .I3(data_in_field[71]), .O(n2733));
    defparam i2482_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i489_3_lut_4_lut (.I0(n3703), .I1(tx2_active), .I2(r_SM_Main_2__N_1770[0]), 
            .I3(\FRAME_MATCHER.wait_for_transmission ), .O(n195));   // coms.v(209[14] 219[8])
    defparam i489_3_lut_4_lut.LUT_INIT = 16'h0355;
    uart_tx tx (.GND_net(GND_net), .r_SM_Main({r_SM_Main}), .r_Clock_Count({Open_1, 
            Open_2, Open_3, Open_4, Open_5, Open_6, Open_7, \r_Clock_Count[1] , 
            Open_8}), .n2388(n2388), .VCC_net(VCC_net), .\r_Clock_Count[8] (\r_Clock_Count[8] ), 
            .CLK_N_keep(CLK_c), .n2418(n2418), .\r_Clock_Count[6] (\r_Clock_Count[6] ), 
            .tx_o(tx_o), .n321(n321), .\r_Clock_Count[0] (\r_Clock_Count[0] ), 
            .\tx_data[0]_N_keep (tx_data[0]), .n1519(n1519), .n2826(n2826), 
            .\r_Tx_Data[3] (\r_Tx_Data[3] ), .n2827(n2827), .\r_Tx_Data[4] (\r_Tx_Data[4] ), 
            .n2447(n2447), .\r_SM_Main_2__N_1770[0] (tx_transmit), .\r_Tx_Data[1] (\r_Tx_Data[1] ), 
            .\r_Tx_Data[2] (\r_Tx_Data[2] ), .tx_enable(tx_enable), .n2825(n2825), 
            .n2824(n2824), .n2830(n2830), .\r_Tx_Data[7] (\r_Tx_Data[7] ), 
            .n2829(n2829), .\r_Tx_Data[6] (\r_Tx_Data[6] ), .n2478(n2478), 
            .tx_active(tx_active), .n2476(n2476), .n2828(n2828), .\r_Tx_Data[5] (\r_Tx_Data[5] ), 
            .\r_Clock_Count[3] (\r_Clock_Count[3] ), .\r_Clock_Count[4] (\r_Clock_Count[4] ), 
            .n2467(n2467), .n2470(n2470), .n313(n313), .n315(n315), 
            .n317(n317), .n11(n11), .n782(n782), .n318(n318), .n5111(n5111), 
            .n4155(n4155), .n320(n320), .n5818(n5818), .n5(n5)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1 */ ;   // coms.v(41[11:71])
    uart_tx_U0 tx2 (.n2450(n2450), .VCC_net(VCC_net), .r_Bit_Index({Open_9, 
            Open_10, \r_Bit_Index[0] }), .CLK_c(CLK_c), .r_SM_Main({\r_SM_Main[2]_adj_11 , 
            Open_11, Open_12}), .GND_net(GND_net), .\r_SM_Main[1] (\r_SM_Main[1]_adj_12 ), 
            .n4544(n4544), .n2486(n2486), .tx2_active(tx2_active), .n313(n313_adj_13), 
            .\r_Clock_Count[8] (\r_Clock_Count[8]_adj_14 ), .\r_SM_Main_2__N_1770[0] (r_SM_Main_2__N_1770[0]), 
            .tx2_o(tx2_o), .n4(n4_adj_15), .n2208(n2208), .n2339(n2339), 
            .tx2_data({tx2_data}), .n2415(n2415), .tx2_enable(tx2_enable)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(190[11:78])
    uart_rx rx (.\r_Bit_Index[0] (\r_Bit_Index[0]_adj_16 ), .GND_net(GND_net), 
            .VCC_net(VCC_net), .CLK_c(CLK_c), .n1757(n1757), .n2836(n2836), 
            .rx_data({rx_data}), .r_SM_Main({r_SM_Main_adj_22}), .\r_SM_Main_2__N_1824[2] (\r_SM_Main_2__N_1824[2] ), 
            .n2837(n2837), .n2834(n2834), .n2833(n2833), .n1764(n1764), 
            .n4(n4_adj_20), .n5089(n5089), .rx_data_ready(rx_data_ready), 
            .n1760(n1760), .n4_adj_1(n4_adj_21), .n2822(n2822), .r_Rx_Data(r_Rx_Data), 
            .rx_i(rx_i), .n3636(n3636), .n5355(n5355), .n2381(n2381), 
            .n2380(n2380), .n2455(n2455)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // coms.v(169[11:45])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (GND_net, r_SM_Main, r_Clock_Count, n2388, VCC_net, 
            \r_Clock_Count[8] , CLK_N_keep, n2418, \r_Clock_Count[6] , 
            tx_o, n321, \r_Clock_Count[0] , \tx_data[0]_N_keep , n1519, 
            n2826, \r_Tx_Data[3] , n2827, \r_Tx_Data[4] , n2447, \r_SM_Main_2__N_1770[0] , 
            \r_Tx_Data[1] , \r_Tx_Data[2] , tx_enable, n2825, n2824, 
            n2830, \r_Tx_Data[7] , n2829, \r_Tx_Data[6] , n2478, tx_active, 
            n2476, n2828, \r_Tx_Data[5] , \r_Clock_Count[3] , \r_Clock_Count[4] , 
            n2467, n2470, n313, n315, n317, n11, n782, n318, 
            n5111, n4155, n320, n5818, n5) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1 */ ;
    input GND_net;
    output [2:0]r_SM_Main;
    output [8:0]r_Clock_Count;
    input n2388;
    input VCC_net;
    output \r_Clock_Count[8] ;
    input CLK_N_keep;
    input n2418;
    output \r_Clock_Count[6] ;
    output tx_o;
    output n321;
    output \r_Clock_Count[0] ;
    input \tx_data[0]_N_keep ;
    output n1519;
    input n2826;
    output \r_Tx_Data[3] ;
    input n2827;
    output \r_Tx_Data[4] ;
    input n2447;
    input \r_SM_Main_2__N_1770[0] ;
    output \r_Tx_Data[1] ;
    output \r_Tx_Data[2] ;
    output tx_enable;
    input n2825;
    input n2824;
    input n2830;
    output \r_Tx_Data[7] ;
    input n2829;
    output \r_Tx_Data[6] ;
    input n2478;
    output tx_active;
    input n2476;
    input n2828;
    output \r_Tx_Data[5] ;
    output \r_Clock_Count[3] ;
    output \r_Clock_Count[4] ;
    input n2467;
    input n2470;
    output n313;
    output n315;
    output n317;
    input n11;
    output n782;
    output n318;
    input n5111;
    output n4155;
    output n320;
    output n5818;
    output n5;
    
    
    wire n6054, n6288;
    wire [2:0]r_Bit_Index;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(33[16:27])
    
    wire o_Tx_Serial_N_1798, n12, n4764, n4765, n3120;
    wire [8:0]r_Clock_Count_c;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    
    wire n15, n10, n5883;
    wire [7:0]r_Tx_Data;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(34[16:25])
    
    wire n2479, n5812, n14, n2880, n6051;
    wire [2:0]r_SM_Main_2__N_1767;
    
    wire n5153, n5885, n2483, n5821, n5095, n5117;
    wire [2:0]n307;
    
    wire n40, n2247, n2356, n3631, n5195, n5357, n5629, n10_adj_1868, 
        n14_adj_1869, n3644, n2177, n6285, n4771, n5884, n4770, 
        n4769, n4768, n4767, n5627, n4766;
    
    SB_LUT4 i367827_i1_3_lut (.I0(n6054), .I1(n6288), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_1798));
    defparam i367827_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26_3_lut (.I0(o_Tx_Serial_N_1798), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n12));
    defparam i26_3_lut.LUT_INIT = 16'h1c1c;
    SB_CARRY add_59_3 (.CI(n4764), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n4765));
    SB_LUT4 i33_3_lut (.I0(r_SM_Main[2]), .I1(n3120), .I2(r_Clock_Count_c[2]), 
            .I3(GND_net), .O(n15));
    defparam i33_3_lut.LUT_INIT = 16'haeae;
    SB_DFFE r_Clock_Count__i8 (.Q(\r_Clock_Count[8] ), .C(CLK_N_keep), .E(VCC_net), 
            .D(n2388));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(\r_Clock_Count[6] ), .C(CLK_N_keep), .D(n2418));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i25_3_lut (.I0(n12), .I1(tx_o), .I2(r_SM_Main[2]), .I3(GND_net), 
            .O(n10));
    defparam i25_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 add_59_2_lut (.I0(GND_net), .I1(\r_Clock_Count[0] ), .I2(GND_net), 
            .I3(VCC_net), .O(n321)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(\r_Clock_Count[0] ), .I1(GND_net), 
            .CO(n4764));
    SB_LUT4 i2845_4_lut (.I0(\tx_data[0]_N_keep ), .I1(n5883), .I2(r_Tx_Data[0]), 
            .I3(n1519), .O(n2479));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(34[16:25])
    defparam i2845_4_lut.LUT_INIT = 16'hcac0;
    SB_DFF r_Tx_Data_i3 (.Q(\r_Tx_Data[3] ), .C(CLK_N_keep), .D(n2826));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i4 (.Q(\r_Tx_Data[4] ), .C(CLK_N_keep), .D(n2827));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Clock_Count__i0 (.Q(\r_Clock_Count[0] ), .C(CLK_N_keep), .E(VCC_net), 
            .D(n2447));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i28_4_lut (.I0(\r_SM_Main_2__N_1770[0] ), .I1(n5812), .I2(r_SM_Main[1]), 
            .I3(r_Bit_Index[0]), .O(n14));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    defparam i28_4_lut.LUT_INIT = 16'hca0a;
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count_c[7]), .C(CLK_N_keep), .D(n2880));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 n6051_bdd_4_lut (.I0(n6051), .I1(\r_Tx_Data[1] ), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n6054));
    defparam n6051_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n14), .I2(r_SM_Main_2__N_1767[1]), 
            .I3(r_SM_Main[0]), .O(n5153));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    defparam i1_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_5889 (.I0(r_Bit_Index[0]), .I1(\r_Tx_Data[2] ), 
            .I2(\r_Tx_Data[3] ), .I3(r_Bit_Index[1]), .O(n6051));
    defparam r_Bit_Index_0__bdd_4_lut_5889.LUT_INIT = 16'he4aa;
    SB_LUT4 i2880_3_lut (.I0(r_Clock_Count_c[2]), .I1(n5885), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n2483));
    defparam i2880_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(tx_enable));
    defparam i8_1_lut.LUT_INIT = 16'h5555;
    SB_DFF r_Tx_Data_i2 (.Q(\r_Tx_Data[2] ), .C(CLK_N_keep), .D(n2825));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i1 (.Q(\r_Tx_Data[1] ), .C(CLK_N_keep), .D(n2824));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i13_4_lut (.I0(r_Clock_Count_c[5]), .I1(n5821), .I2(r_SM_Main[2]), 
            .I3(r_Clock_Count_c[2]), .O(n5095));
    defparam i13_4_lut.LUT_INIT = 16'ha0ac;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_N_keep), .D(n5117));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i15_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(33[16:27])
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n40));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2105_4_lut (.I0(n2247), .I1(r_SM_Main[1]), .I2(r_Bit_Index[0]), 
            .I3(n40), .O(n2356));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2105_4_lut.LUT_INIT = 16'ha222;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_1767[1]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n2247));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i3227_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n307[2]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(33[16:27])
    defparam i3227_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i3388_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(GND_net), 
            .I3(GND_net), .O(n3631));
    defparam i3388_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_N_keep), .D(n5195));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i7 (.Q(\r_Tx_Data[7] ), .C(CLK_N_keep), .D(n2830));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_N_keep), .E(n2247), 
            .D(n307[2]), .R(n2356));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_N_keep), .E(n2247), 
            .D(n307[1]), .R(n2356));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count_c[5]), .C(CLK_N_keep), .D(n5095));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i6 (.Q(\r_Tx_Data[6] ), .C(CLK_N_keep), .D(n2829));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count_c[2]), .C(CLK_N_keep), .D(n2483));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_N_keep), .D(n5153));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_N_keep), .D(n2479));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_N_keep), .D(n2478));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(CLK_N_keep), .D(n10));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_N_keep), .E(VCC_net), 
            .D(n2476));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Data_i5 (.Q(\r_Tx_Data[5] ), .C(CLK_N_keep), .D(n2828));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_N_keep), .D(n5357));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i5283_3_lut_4_lut (.I0(r_Clock_Count[1]), .I1(\r_Clock_Count[0] ), 
            .I2(\r_Clock_Count[3] ), .I3(r_Clock_Count_c[7]), .O(n5629));
    defparam i5283_3_lut_4_lut.LUT_INIT = 16'hfff8;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_1770[0] ), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n1519));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i2_2_lut (.I0(\r_Clock_Count[8] ), .I1(\r_Clock_Count[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_1868));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(r_Clock_Count_c[2]), .I1(r_Clock_Count_c[7]), 
            .I2(\r_Clock_Count[4] ), .I3(\r_Clock_Count[6] ), .O(n14_adj_1869));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n3644), .I1(n14_adj_1869), .I2(n10_adj_1868), 
            .I3(r_Clock_Count_c[5]), .O(r_SM_Main_2__N_1767[1]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_804 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_1767[1]), .O(n2177));
    defparam i2_4_lut_adj_804.LUT_INIT = 16'h1101;
    SB_LUT4 i12_3_lut (.I0(n2177), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n5117));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 i5592_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_1770[0] ), 
            .I2(n3631), .I3(\tx_data[0]_N_keep ), .O(n5883));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i5592_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_DFF r_Clock_Count__i4 (.Q(\r_Clock_Count[4] ), .C(CLK_N_keep), .D(n2467));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(\r_Clock_Count[3] ), .C(CLK_N_keep), .D(n2470));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(\r_Tx_Data[6] ), 
            .I2(\r_Tx_Data[7] ), .I3(r_Bit_Index[1]), .O(n6285));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n6285_bdd_4_lut (.I0(n6285), .I1(\r_Tx_Data[5] ), .I2(\r_Tx_Data[4] ), 
            .I3(r_Bit_Index[1]), .O(n6288));
    defparam n6285_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(\r_Clock_Count[8] ), .I2(GND_net), 
            .I3(n4771), .O(n313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_59_9_lut (.I0(n15), .I1(r_Clock_Count_c[7]), .I2(GND_net), 
            .I3(n4770), .O(n5884)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_9 (.CI(n4770), .I0(r_Clock_Count_c[7]), .I1(GND_net), 
            .CO(n4771));
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(\r_Clock_Count[6] ), .I2(GND_net), 
            .I3(n4769), .O(n315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_8 (.CI(n4769), .I0(\r_Clock_Count[6] ), .I1(GND_net), 
            .CO(n4770));
    SB_LUT4 add_59_7_lut (.I0(n3120), .I1(r_Clock_Count_c[5]), .I2(GND_net), 
            .I3(n4768), .O(n5821)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_7 (.CI(n4768), .I0(r_Clock_Count_c[5]), .I1(GND_net), 
            .CO(n4769));
    SB_LUT4 add_59_6_lut (.I0(GND_net), .I1(\r_Clock_Count[4] ), .I2(GND_net), 
            .I3(n4767), .O(n317)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_6 (.CI(n4767), .I0(\r_Clock_Count[4] ), .I1(GND_net), 
            .CO(n4768));
    SB_LUT4 i2874_3_lut (.I0(r_Clock_Count_c[7]), .I1(n5884), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n2880));
    defparam i2874_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3401_2_lut (.I0(r_Clock_Count[1]), .I1(\r_Clock_Count[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n3644));
    defparam i3401_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5281_4_lut (.I0(r_Clock_Count_c[5]), .I1(\r_Clock_Count[8] ), 
            .I2(\r_Clock_Count[6] ), .I3(\r_Clock_Count[4] ), .O(n5627));
    defparam i5281_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_805 (.I0(n5629), .I1(r_SM_Main[2]), .I2(n5627), 
            .I3(n11), .O(n3120));
    defparam i2_4_lut_adj_805.LUT_INIT = 16'h0100;
    SB_LUT4 i1_3_lut (.I0(r_SM_Main[2]), .I1(r_Clock_Count_c[2]), .I2(n3120), 
            .I3(GND_net), .O(n782));
    defparam i1_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(\r_Clock_Count[3] ), .I2(GND_net), 
            .I3(n4766), .O(n318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n4766), .I0(\r_Clock_Count[3] ), .I1(GND_net), 
            .CO(n4767));
    SB_LUT4 add_59_4_lut (.I0(n15), .I1(r_Clock_Count_c[2]), .I2(GND_net), 
            .I3(n4765), .O(n5885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'h8228;
    SB_DFFE r_Tx_Done_44 (.Q(n4155), .C(CLK_N_keep), .E(VCC_net), .D(n5111));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_4 (.CI(n4765), .I0(r_Clock_Count_c[2]), .I1(GND_net), 
            .CO(n4766));
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n4764), .O(n320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5566_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_1767[1]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n5818));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    defparam i5566_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_1767[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n5357));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i1_3_lut_4_lut_adj_806 (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_1767[1]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n5195));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    defparam i1_3_lut_4_lut_adj_806.LUT_INIT = 16'h0078;
    SB_LUT4 i16_3_lut_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_1767[1]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_1770[0] ), .O(n5));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    defparam i16_3_lut_4_lut_4_lut.LUT_INIT = 16'h8580;
    SB_LUT4 i5604_2_lut_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_SM_Main_2__N_1767[1]), .I3(GND_net), .O(n5812));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    defparam i5604_2_lut_3_lut.LUT_INIT = 16'h8080;
    
endmodule
//
// Verilog Description of module uart_tx_U0
//

module uart_tx_U0 (n2450, VCC_net, r_Bit_Index, CLK_c, r_SM_Main, 
            GND_net, \r_SM_Main[1] , n4544, n2486, tx2_active, n313, 
            \r_Clock_Count[8] , \r_SM_Main_2__N_1770[0] , tx2_o, n4, 
            n2208, n2339, tx2_data, n2415, tx2_enable) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n2450;
    input VCC_net;
    output [2:0]r_Bit_Index;
    input CLK_c;
    output [2:0]r_SM_Main;
    input GND_net;
    output \r_SM_Main[1] ;
    output n4544;
    input n2486;
    output tx2_active;
    output n313;
    output \r_Clock_Count[8] ;
    input \r_SM_Main_2__N_1770[0] ;
    output tx2_o;
    output n4;
    output n2208;
    output n2339;
    input [7:0]tx2_data;
    input n2415;
    output tx2_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [8:0]r_Clock_Count;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    
    wire n5824, n5061, n2444;
    wire [2:0]r_SM_Main_c;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    wire [2:0]r_SM_Main_2__N_1767;
    
    wire n6314;
    wire [8:0]n312;
    
    wire n2427, n2441, n2424, n2431;
    wire [2:0]r_Bit_Index_c;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(33[16:27])
    wire [2:0]n307;
    
    wire n4786, n5847, n4785, n1136, n14, n5189, n4784;
    wire [7:0]r_Tx_Data;   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(34[16:25])
    
    wire n6045, n2434, n5203, n2438, n4783, n10, n1624, n6048, 
        n6006, o_Tx_Serial_N_1798, n12, n31, n5631, n9, n78, n4782, 
        n4781, n4780, n5816, n4779, n6003, n14_adj_1867;
    
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .E(VCC_net), 
            .D(n2450));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i18_3_lut (.I0(r_Clock_Count[0]), .I1(n5824), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n5061));
    defparam i18_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(VCC_net), 
            .D(n2444));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_c[0]), .I2(\r_SM_Main[1] ), 
            .I3(r_SM_Main_2__N_1767[1]), .O(n6314));
    defparam i3_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i1_4_lut (.I0(n4544), .I1(r_Clock_Count[6]), .I2(n312[6]), 
            .I3(r_SM_Main[2]), .O(n2427));
    defparam i1_4_lut.LUT_INIT = 16'h88a0;
    SB_DFFE r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(VCC_net), 
            .D(n2441));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx2_active), .C(CLK_c), .D(n2486));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_4_lut_adj_795 (.I0(n4544), .I1(r_Clock_Count[7]), .I2(n312[7]), 
            .I3(r_SM_Main[2]), .O(n2424));
    defparam i1_4_lut_adj_795.LUT_INIT = 16'h88a0;
    SB_LUT4 i1_4_lut_adj_796 (.I0(n4544), .I1(r_Clock_Count[5]), .I2(n312[5]), 
            .I3(r_SM_Main[2]), .O(n2431));
    defparam i1_4_lut_adj_796.LUT_INIT = 16'h88a0;
    SB_LUT4 i615_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(98[36:51])
    defparam i615_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(\r_Clock_Count[8] ), .I2(GND_net), 
            .I3(n4786), .O(n313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5567_2_lut (.I0(r_SM_Main_2__N_1767[1]), .I1(r_Bit_Index[0]), 
            .I2(GND_net), .I3(GND_net), .O(n5847));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(33[16:27])
    defparam i5567_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n4785), .O(n312[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28_4_lut (.I0(\r_SM_Main_2__N_1770[0] ), .I1(n5847), .I2(\r_SM_Main[1] ), 
            .I3(n1136), .O(n14));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(33[16:27])
    defparam i28_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut_adj_797 (.I0(r_SM_Main[2]), .I1(n14), .I2(r_SM_Main_2__N_1767[1]), 
            .I3(r_SM_Main_c[0]), .O(n5189));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(33[16:27])
    defparam i1_4_lut_adj_797.LUT_INIT = 16'h0544;
    SB_CARRY add_59_9 (.CI(n4785), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n4786));
    SB_LUT4 i622_3_lut (.I0(r_Bit_Index_c[2]), .I1(r_Bit_Index_c[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n307[2]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(98[36:51])
    defparam i622_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n4784), .O(n312[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index_c[1]), .O(n6045));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_798 (.I0(n4544), .I1(r_Clock_Count[4]), .I2(n312[4]), 
            .I3(r_SM_Main[2]), .O(n2434));
    defparam i1_4_lut_adj_798.LUT_INIT = 16'h88a0;
    SB_CARRY add_59_8 (.CI(n4784), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n4785));
    SB_DFF r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(CLK_c), .D(n5203));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(VCC_net), 
            .D(n2438));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n4783), .O(n312[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF o_Tx_Serial_45 (.Q(tx2_o), .C(CLK_c), .D(n10));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main_c[0]), .I1(\r_SM_Main_2__N_1770[0] ), 
            .I2(\r_SM_Main[1] ), .I3(r_SM_Main[2]), .O(n1624));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 n6045_bdd_4_lut (.I0(n6045), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index_c[1]), .O(n6048));
    defparam n6045_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5614_4_lut_4_lut (.I0(r_SM_Main_c[0]), .I1(\r_SM_Main_2__N_1770[0] ), 
            .I2(\r_SM_Main[1] ), .I3(r_SM_Main_2__N_1767[1]), .O(n4));
    defparam i5614_4_lut_4_lut.LUT_INIT = 16'ha404;
    SB_LUT4 i367224_i1_3_lut (.I0(n6048), .I1(n6006), .I2(r_Bit_Index_c[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_1798));
    defparam i367224_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26_3_lut (.I0(r_SM_Main_c[0]), .I1(o_Tx_Serial_N_1798), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n12));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    defparam i26_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i25_3_lut (.I0(n12), .I1(tx2_o), .I2(r_SM_Main[2]), .I3(GND_net), 
            .O(n10));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    defparam i25_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i5285_4_lut (.I0(r_Clock_Count[7]), .I1(\r_Clock_Count[8] ), 
            .I2(n31), .I3(r_Clock_Count[6]), .O(n5631));
    defparam i5285_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_799 (.I0(r_Clock_Count[3]), .I1(\r_SM_Main[1] ), 
            .I2(r_Clock_Count[4]), .I3(r_SM_Main_c[0]), .O(n9));
    defparam i3_4_lut_adj_799.LUT_INIT = 16'h0504;
    SB_LUT4 i1_4_lut_adj_800 (.I0(r_SM_Main[2]), .I1(n78), .I2(n9), .I3(n5631), 
            .O(n4544));
    defparam i1_4_lut_adj_800.LUT_INIT = 16'haaba;
    SB_CARRY add_59_7 (.CI(n4783), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n4784));
    SB_DFFE r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(VCC_net), 
            .D(n2434));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_4_lut_adj_801 (.I0(n4544), .I1(r_Clock_Count[3]), .I2(n312[3]), 
            .I3(r_SM_Main[2]), .O(n2438));
    defparam i1_4_lut_adj_801.LUT_INIT = 16'h88a0;
    SB_LUT4 i1_4_lut_adj_802 (.I0(n4544), .I1(r_Clock_Count[2]), .I2(n312[2]), 
            .I3(r_SM_Main[2]), .O(n2441));
    defparam i1_4_lut_adj_802.LUT_INIT = 16'h88a0;
    SB_DFFE r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(VCC_net), 
            .D(n2431));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n4782), .O(n312[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .D(n2424));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_6 (.CI(n4782), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n4783));
    SB_DFFE r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(VCC_net), 
            .D(n2427));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n6314));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n4781), .O(n312[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n4781), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n4782));
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n4780), .O(n312[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_4 (.CI(n4780), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n4781));
    SB_LUT4 add_59_3_lut (.I0(n4544), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n4779), .O(n5816)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'h8228;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(CLK_c), .E(n2208), 
            .D(n307[2]), .R(n2339));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_3 (.CI(n4779), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n4780));
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(CLK_c), .D(n5189));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_2_lut (.I0(n4544), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n5824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'h8228;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(CLK_c), .E(n2208), 
            .D(n307[1]), .R(n2339));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n4779));
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n1624), .D(tx2_data[0]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_4_lut_adj_803 (.I0(r_SM_Main[2]), .I1(\r_SM_Main[1] ), .I2(r_SM_Main_2__N_1767[1]), 
            .I3(r_SM_Main_c[0]), .O(n5203));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(31[16:25])
    defparam i1_4_lut_adj_803.LUT_INIT = 16'h1444;
    SB_LUT4 i4294_3_lut (.I0(r_Clock_Count[1]), .I1(n5816), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n2444));
    defparam i4294_3_lut.LUT_INIT = 16'hacac;
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .D(n5061));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_5690 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index_c[1]), .O(n6003));
    defparam r_Bit_Index_0__bdd_4_lut_5690.LUT_INIT = 16'he4aa;
    SB_LUT4 n6003_bdd_4_lut (.I0(n6003), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index_c[1]), .O(n6006));
    defparam n6003_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i895_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1136));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(96[21:36])
    defparam i895_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i85_2_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(GND_net), .O(n78));
    defparam i85_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(32[16:29])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut (.I0(\r_Clock_Count[8] ), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[3]), 
            .I3(r_Clock_Count[6]), .O(n14_adj_1867));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n31), .I1(n14_adj_1867), .I2(n78), .I3(r_Clock_Count[4]), 
            .O(r_SM_Main_2__N_1767[1]));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main_2__N_1767[1]), .I1(r_SM_Main_c[0]), 
            .I2(\r_SM_Main[1] ), .I3(r_SM_Main[2]), .O(n2208));
    defparam i2_4_lut.LUT_INIT = 16'h0023;
    SB_LUT4 i2088_4_lut (.I0(n2208), .I1(r_Bit_Index[0]), .I2(\r_SM_Main[1] ), 
            .I3(n1136), .O(n2339));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    defparam i2088_4_lut.LUT_INIT = 16'h8a0a;
    SB_DFF r_Clock_Count__i8 (.Q(\r_Clock_Count[8] ), .C(CLK_c), .D(n2415));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n1624), .D(tx2_data[1]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n1624), .D(tx2_data[2]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n1624), .D(tx2_data[3]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n1624), .D(tx2_data[4]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n1624), .D(tx2_data[5]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n1624), .D(tx2_data[6]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n1624), .D(tx2_data[7]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(40[10] 143[8])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx2_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx2_enable));   // roboy_fpga_code/roboy_fpga_code/uart/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (\r_Bit_Index[0] , GND_net, VCC_net, CLK_c, n1757, 
            n2836, rx_data, r_SM_Main, \r_SM_Main_2__N_1824[2] , n2837, 
            n2834, n2833, n1764, n4, n5089, rx_data_ready, n1760, 
            n4_adj_1, n2822, r_Rx_Data, rx_i, n3636, n5355, n2381, 
            n2380, n2455) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output \r_Bit_Index[0] ;
    input GND_net;
    input VCC_net;
    input CLK_c;
    output n1757;
    input n2836;
    output [7:0]rx_data;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_1824[2] ;
    input n2837;
    input n2834;
    input n2833;
    output n1764;
    output n4;
    input n5089;
    output rx_data_ready;
    output n1760;
    output n4_adj_1;
    input n2822;
    output r_Rx_Data;
    input rx_i;
    output n3636;
    input n5355;
    input n2381;
    input n2380;
    input n2455;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]r_Bit_Index;   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(33[17:28])
    wire [2:0]n326;
    
    wire n2453, n1706;
    wire [7:0]r_Clock_Count;   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(32[17:30])
    
    wire n5860, n359, n4284, n5855, n2502, n2881, n5069, n6294, 
        n5613, n2879, n2878, n5361, n17, n1724, n5817, n36, 
        n2877, n2876;
    wire [2:0]r_SM_Main_2__N_1821;
    
    wire n5857, n75, n3589, n5815, n5856, n3850, n6291, n5858, 
        r_Rx_Data_R, n5859, n4778, n5854, n4777, n2259, n2367, 
        n4776, n4775, n4774, n5823, n5822, n4773, n4772, n8, 
        n5633;
    
    SB_LUT4 i593_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(102[36:51])
    defparam i593_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .E(VCC_net), 
            .D(n2453));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[2]), .I1(n1706), .I2(r_Bit_Index[1]), 
            .I3(GND_net), .O(n1757));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(52[7] 143[14])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n2836));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 i4017_3_lut (.I0(r_Clock_Count[1]), .I1(n5860), .I2(n359), 
            .I3(GND_net), .O(n4284));
    defparam i4017_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3997_3_lut (.I0(r_Clock_Count[0]), .I1(n5855), .I2(n359), 
            .I3(GND_net), .O(n2502));
    defparam i3997_3_lut.LUT_INIT = 16'hacac;
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .D(n2881));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .D(n5069));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 i5636_2_lut (.I0(r_SM_Main[2]), .I1(n6294), .I2(GND_net), 
            .I3(GND_net), .O(n5613));
    defparam i5636_2_lut.LUT_INIT = 16'h1111;
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .D(n2879));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .D(n2878));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5361));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(36[17:26])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5574_4_lut (.I0(r_SM_Main[0]), .I1(n17), .I2(n5361), .I3(n1724), 
            .O(n5817));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(36[17:26])
    defparam i5574_4_lut.LUT_INIT = 16'h55d5;
    SB_LUT4 i16_4_lut (.I0(r_SM_Main[2]), .I1(n5817), .I2(\r_SM_Main_2__N_1824[2] ), 
            .I3(r_SM_Main[1]), .O(n36));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(36[17:26])
    defparam i16_4_lut.LUT_INIT = 16'hafbb;
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .D(n2877));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n2837));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n2834));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n2833));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .D(n2876));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(r_SM_Main_2__N_1821[1]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut_adj_791 (.I0(n1706), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n1764));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_791.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_1824[2] ), .O(n1706));
    defparam i2_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 equal_27_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(97[17:39])
    defparam equal_27_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .E(VCC_net), .D(n5089));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_2_lut_adj_792 (.I0(\r_Bit_Index[0] ), .I1(n1706), .I2(GND_net), 
            .I3(GND_net), .O(n1760));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_792.LUT_INIT = 16'heeee;
    SB_LUT4 equal_26_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(97[17:39])
    defparam equal_26_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n2822));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 i4005_3_lut (.I0(r_Clock_Count[4]), .I1(n5857), .I2(n359), 
            .I3(GND_net), .O(n2877));
    defparam i4005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i90_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_1824[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n75));
    defparam i90_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5560_2_lut (.I0(r_Rx_Data), .I1(n3589), .I2(GND_net), .I3(GND_net), 
            .O(n5815));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(36[17:26])
    defparam i5560_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n5815), .I2(n75), .I3(r_SM_Main[1]), 
            .O(r_SM_Main_2__N_1821[1]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(36[17:26])
    defparam i1_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i4001_3_lut (.I0(r_Clock_Count[3]), .I1(n5856), .I2(n359), 
            .I3(GND_net), .O(n2876));
    defparam i4001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut (.I0(\r_SM_Main_2__N_1824[2] ), .I1(n3850), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n6291));
    defparam r_SM_Main_0__bdd_4_lut_4_lut.LUT_INIT = 16'haf70;
    SB_LUT4 i4009_3_lut (.I0(r_Clock_Count[5]), .I1(n5858), .I2(n359), 
            .I3(GND_net), .O(n2878));
    defparam i4009_3_lut.LUT_INIT = 16'hacac;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n5613));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(rx_i));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(41[10] 45[8])
    SB_LUT4 add_62_9_lut (.I0(n36), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n4778), .O(n5859)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(n36), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n4777), .O(n5854)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'h8228;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n2259), 
            .D(n326[2]), .R(n2367));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_CARRY add_62_8 (.CI(n4777), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n4778));
    SB_LUT4 i3393_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n3636));
    defparam i3393_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3992_3_lut (.I0(r_Clock_Count[6]), .I1(n5854), .I2(n359), 
            .I3(GND_net), .O(n2879));
    defparam i3992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_62_7_lut (.I0(n36), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n4776), .O(n5858)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_7 (.CI(n4776), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n4777));
    SB_LUT4 add_62_6_lut (.I0(n36), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n4775), .O(n5857)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n4775), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n4776));
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .D(n2502));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_5_lut (.I0(n36), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n4774), .O(n5856)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'h8228;
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .D(n4284));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_CARRY add_62_5 (.CI(n4774), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n4775));
    SB_LUT4 n6291_bdd_4_lut (.I0(n6291), .I1(n5823), .I2(r_Rx_Data), .I3(r_SM_Main[1]), 
            .O(n6294));
    defparam n6291_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n5355));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_4_lut (.I0(n36), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n4773), .O(n5822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'h8228;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n2381));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n2380));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_CARRY add_62_4 (.CI(n4773), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n4774));
    SB_LUT4 add_62_3_lut (.I0(n36), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n4772), .O(n5860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_3 (.CI(n4772), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n4773));
    SB_LUT4 add_62_2_lut (.I0(n36), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n5855)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n4772));
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n2259), 
            .D(n326[1]), .R(n2367));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 i11_3_lut (.I0(n5822), .I1(r_Clock_Count[2]), .I2(n359), .I3(GND_net), 
            .O(n5069));
    defparam i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_793 (.I0(r_Rx_Data), .I1(r_SM_Main[2]), .I2(n3589), 
            .I3(r_SM_Main[1]), .O(n359));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(36[17:26])
    defparam i1_4_lut_adj_793.LUT_INIT = 16'hccec;
    SB_LUT4 i4013_3_lut (.I0(r_Clock_Count[7]), .I1(n5859), .I2(n359), 
            .I3(GND_net), .O(n2881));
    defparam i4013_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut (.I0(r_Clock_Count[0]), .I1(n1724), .I2(r_Clock_Count[1]), 
            .I3(r_Rx_Data), .O(n17));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_4_lut_adj_794 (.I0(r_Clock_Count[0]), .I1(n1724), .I2(r_Clock_Count[1]), 
            .I3(r_SM_Main[0]), .O(n3589));
    defparam i1_2_lut_4_lut_adj_794.LUT_INIT = 16'h0200;
    SB_LUT4 i3_3_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[4]), .I2(r_Clock_Count[3]), 
            .I3(GND_net), .O(n8));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5277_4_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[2]), .I2(n8), 
            .I3(r_Clock_Count[5]), .O(n1724));
    defparam i5277_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[1]), .I1(n1724), .I2(r_Clock_Count[0]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_1824[2] ));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(32[17:30])
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i2116_2_lut_3_lut (.I0(n3850), .I1(r_SM_Main[1]), .I2(n2259), 
            .I3(GND_net), .O(n2367));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(52[7] 143[14])
    defparam i2116_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i2202_3_lut_4_lut (.I0(n3850), .I1(r_SM_Main[1]), .I2(\r_Bit_Index[0] ), 
            .I3(n5633), .O(n2453));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(52[7] 143[14])
    defparam i2202_3_lut_4_lut.LUT_INIT = 16'hf004;
    SB_LUT4 i600_2_lut_3_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n326[2]));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(102[36:51])
    defparam i600_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n3850));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(102[36:51])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1824[2] ), .O(n2259));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i5287_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_1824[2] ), .O(n5633));
    defparam i5287_3_lut_4_lut.LUT_INIT = 16'heefe;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n2455));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(49[10] 144[8])
    SB_LUT4 i5570_2_lut_3_lut (.I0(n1724), .I1(r_Clock_Count[0]), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n5823));   // roboy_fpga_code/roboy_fpga_code/uart/uart_rx.v(36[17:26])
    defparam i5570_2_lut_3_lut.LUT_INIT = 16'h0404;
    
endmodule
