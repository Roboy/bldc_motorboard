// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Aug 26 2019 01:17:31

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    inout PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    inout PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    inout PIN_1;
    output LED;
    input CLK;

    wire N__37951;
    wire N__37950;
    wire N__37949;
    wire N__37942;
    wire N__37941;
    wire N__37940;
    wire N__37933;
    wire N__37932;
    wire N__37931;
    wire N__37924;
    wire N__37923;
    wire N__37922;
    wire N__37915;
    wire N__37914;
    wire N__37913;
    wire N__37906;
    wire N__37905;
    wire N__37904;
    wire N__37887;
    wire N__37884;
    wire N__37881;
    wire N__37880;
    wire N__37877;
    wire N__37874;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37857;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37808;
    wire N__37805;
    wire N__37802;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37764;
    wire N__37761;
    wire N__37758;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37745;
    wire N__37740;
    wire N__37737;
    wire N__37736;
    wire N__37735;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37727;
    wire N__37726;
    wire N__37721;
    wire N__37718;
    wire N__37717;
    wire N__37716;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37708;
    wire N__37707;
    wire N__37706;
    wire N__37705;
    wire N__37704;
    wire N__37703;
    wire N__37702;
    wire N__37699;
    wire N__37696;
    wire N__37693;
    wire N__37686;
    wire N__37681;
    wire N__37676;
    wire N__37673;
    wire N__37666;
    wire N__37663;
    wire N__37658;
    wire N__37641;
    wire N__37638;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37623;
    wire N__37622;
    wire N__37621;
    wire N__37620;
    wire N__37619;
    wire N__37618;
    wire N__37617;
    wire N__37616;
    wire N__37615;
    wire N__37614;
    wire N__37613;
    wire N__37612;
    wire N__37611;
    wire N__37610;
    wire N__37609;
    wire N__37608;
    wire N__37607;
    wire N__37606;
    wire N__37605;
    wire N__37604;
    wire N__37603;
    wire N__37602;
    wire N__37601;
    wire N__37600;
    wire N__37599;
    wire N__37598;
    wire N__37597;
    wire N__37596;
    wire N__37595;
    wire N__37594;
    wire N__37593;
    wire N__37592;
    wire N__37591;
    wire N__37590;
    wire N__37589;
    wire N__37588;
    wire N__37587;
    wire N__37586;
    wire N__37585;
    wire N__37584;
    wire N__37583;
    wire N__37582;
    wire N__37581;
    wire N__37580;
    wire N__37579;
    wire N__37578;
    wire N__37577;
    wire N__37576;
    wire N__37575;
    wire N__37574;
    wire N__37573;
    wire N__37572;
    wire N__37571;
    wire N__37570;
    wire N__37569;
    wire N__37568;
    wire N__37567;
    wire N__37566;
    wire N__37565;
    wire N__37564;
    wire N__37563;
    wire N__37562;
    wire N__37561;
    wire N__37560;
    wire N__37559;
    wire N__37558;
    wire N__37557;
    wire N__37556;
    wire N__37555;
    wire N__37554;
    wire N__37553;
    wire N__37552;
    wire N__37551;
    wire N__37550;
    wire N__37549;
    wire N__37548;
    wire N__37547;
    wire N__37546;
    wire N__37545;
    wire N__37544;
    wire N__37543;
    wire N__37542;
    wire N__37541;
    wire N__37540;
    wire N__37539;
    wire N__37538;
    wire N__37537;
    wire N__37536;
    wire N__37535;
    wire N__37534;
    wire N__37533;
    wire N__37532;
    wire N__37531;
    wire N__37530;
    wire N__37529;
    wire N__37528;
    wire N__37527;
    wire N__37526;
    wire N__37525;
    wire N__37524;
    wire N__37523;
    wire N__37522;
    wire N__37521;
    wire N__37520;
    wire N__37519;
    wire N__37518;
    wire N__37517;
    wire N__37516;
    wire N__37515;
    wire N__37514;
    wire N__37513;
    wire N__37512;
    wire N__37511;
    wire N__37510;
    wire N__37509;
    wire N__37508;
    wire N__37507;
    wire N__37506;
    wire N__37505;
    wire N__37504;
    wire N__37503;
    wire N__37502;
    wire N__37501;
    wire N__37500;
    wire N__37499;
    wire N__37498;
    wire N__37497;
    wire N__37496;
    wire N__37495;
    wire N__37494;
    wire N__37493;
    wire N__37492;
    wire N__37491;
    wire N__37490;
    wire N__37489;
    wire N__37488;
    wire N__37487;
    wire N__37486;
    wire N__37485;
    wire N__37484;
    wire N__37483;
    wire N__37482;
    wire N__37481;
    wire N__37480;
    wire N__37479;
    wire N__37478;
    wire N__37477;
    wire N__37476;
    wire N__37475;
    wire N__37474;
    wire N__37473;
    wire N__37472;
    wire N__37471;
    wire N__37470;
    wire N__37469;
    wire N__37468;
    wire N__37467;
    wire N__37466;
    wire N__37465;
    wire N__37464;
    wire N__37463;
    wire N__37462;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37089;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37047;
    wire N__37044;
    wire N__37041;
    wire N__37038;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37026;
    wire N__37023;
    wire N__37020;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36987;
    wire N__36984;
    wire N__36981;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36969;
    wire N__36966;
    wire N__36965;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36954;
    wire N__36949;
    wire N__36946;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36924;
    wire N__36921;
    wire N__36912;
    wire N__36911;
    wire N__36910;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36902;
    wire N__36901;
    wire N__36900;
    wire N__36899;
    wire N__36898;
    wire N__36897;
    wire N__36896;
    wire N__36895;
    wire N__36894;
    wire N__36893;
    wire N__36892;
    wire N__36887;
    wire N__36884;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36855;
    wire N__36852;
    wire N__36849;
    wire N__36842;
    wire N__36837;
    wire N__36832;
    wire N__36829;
    wire N__36828;
    wire N__36827;
    wire N__36826;
    wire N__36825;
    wire N__36814;
    wire N__36811;
    wire N__36806;
    wire N__36801;
    wire N__36792;
    wire N__36791;
    wire N__36790;
    wire N__36789;
    wire N__36788;
    wire N__36787;
    wire N__36786;
    wire N__36785;
    wire N__36784;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36772;
    wire N__36771;
    wire N__36770;
    wire N__36769;
    wire N__36768;
    wire N__36763;
    wire N__36756;
    wire N__36753;
    wire N__36752;
    wire N__36749;
    wire N__36748;
    wire N__36745;
    wire N__36742;
    wire N__36733;
    wire N__36732;
    wire N__36731;
    wire N__36724;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36708;
    wire N__36703;
    wire N__36696;
    wire N__36687;
    wire N__36684;
    wire N__36683;
    wire N__36682;
    wire N__36681;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36667;
    wire N__36666;
    wire N__36663;
    wire N__36654;
    wire N__36649;
    wire N__36642;
    wire N__36641;
    wire N__36640;
    wire N__36639;
    wire N__36636;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36615;
    wire N__36614;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36600;
    wire N__36591;
    wire N__36588;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36570;
    wire N__36567;
    wire N__36566;
    wire N__36565;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36555;
    wire N__36554;
    wire N__36551;
    wire N__36550;
    wire N__36547;
    wire N__36542;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36526;
    wire N__36519;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36508;
    wire N__36507;
    wire N__36506;
    wire N__36501;
    wire N__36500;
    wire N__36499;
    wire N__36496;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36458;
    wire N__36455;
    wire N__36450;
    wire N__36441;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36430;
    wire N__36427;
    wire N__36424;
    wire N__36421;
    wire N__36414;
    wire N__36413;
    wire N__36412;
    wire N__36409;
    wire N__36408;
    wire N__36403;
    wire N__36400;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36392;
    wire N__36391;
    wire N__36390;
    wire N__36387;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36371;
    wire N__36368;
    wire N__36357;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36276;
    wire N__36275;
    wire N__36272;
    wire N__36269;
    wire N__36264;
    wire N__36261;
    wire N__36260;
    wire N__36257;
    wire N__36252;
    wire N__36249;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36230;
    wire N__36225;
    wire N__36222;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36210;
    wire N__36207;
    wire N__36204;
    wire N__36201;
    wire N__36198;
    wire N__36195;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36176;
    wire N__36175;
    wire N__36174;
    wire N__36173;
    wire N__36170;
    wire N__36169;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36150;
    wire N__36147;
    wire N__36140;
    wire N__36135;
    wire N__36132;
    wire N__36125;
    wire N__36120;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36112;
    wire N__36111;
    wire N__36110;
    wire N__36109;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36097;
    wire N__36094;
    wire N__36089;
    wire N__36082;
    wire N__36075;
    wire N__36074;
    wire N__36073;
    wire N__36072;
    wire N__36071;
    wire N__36070;
    wire N__36069;
    wire N__36068;
    wire N__36065;
    wire N__36064;
    wire N__36063;
    wire N__36062;
    wire N__36059;
    wire N__36058;
    wire N__36057;
    wire N__36056;
    wire N__36055;
    wire N__36054;
    wire N__36053;
    wire N__36052;
    wire N__36049;
    wire N__36048;
    wire N__36047;
    wire N__36046;
    wire N__36045;
    wire N__36044;
    wire N__36043;
    wire N__36040;
    wire N__36035;
    wire N__36032;
    wire N__36025;
    wire N__36024;
    wire N__36023;
    wire N__36022;
    wire N__36021;
    wire N__36020;
    wire N__36019;
    wire N__36016;
    wire N__36015;
    wire N__36014;
    wire N__36011;
    wire N__36008;
    wire N__36001;
    wire N__36000;
    wire N__35999;
    wire N__35992;
    wire N__35987;
    wire N__35984;
    wire N__35983;
    wire N__35982;
    wire N__35981;
    wire N__35980;
    wire N__35979;
    wire N__35978;
    wire N__35977;
    wire N__35976;
    wire N__35975;
    wire N__35974;
    wire N__35971;
    wire N__35966;
    wire N__35965;
    wire N__35964;
    wire N__35963;
    wire N__35962;
    wire N__35957;
    wire N__35948;
    wire N__35945;
    wire N__35944;
    wire N__35943;
    wire N__35942;
    wire N__35941;
    wire N__35940;
    wire N__35939;
    wire N__35936;
    wire N__35935;
    wire N__35934;
    wire N__35933;
    wire N__35932;
    wire N__35931;
    wire N__35930;
    wire N__35929;
    wire N__35928;
    wire N__35927;
    wire N__35926;
    wire N__35925;
    wire N__35924;
    wire N__35923;
    wire N__35920;
    wire N__35919;
    wire N__35918;
    wire N__35911;
    wire N__35908;
    wire N__35907;
    wire N__35906;
    wire N__35905;
    wire N__35904;
    wire N__35903;
    wire N__35902;
    wire N__35901;
    wire N__35900;
    wire N__35899;
    wire N__35894;
    wire N__35887;
    wire N__35884;
    wire N__35881;
    wire N__35880;
    wire N__35879;
    wire N__35878;
    wire N__35877;
    wire N__35876;
    wire N__35869;
    wire N__35862;
    wire N__35857;
    wire N__35854;
    wire N__35853;
    wire N__35850;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35836;
    wire N__35831;
    wire N__35830;
    wire N__35829;
    wire N__35828;
    wire N__35827;
    wire N__35826;
    wire N__35825;
    wire N__35824;
    wire N__35823;
    wire N__35822;
    wire N__35821;
    wire N__35820;
    wire N__35819;
    wire N__35818;
    wire N__35817;
    wire N__35816;
    wire N__35813;
    wire N__35812;
    wire N__35809;
    wire N__35802;
    wire N__35797;
    wire N__35792;
    wire N__35789;
    wire N__35782;
    wire N__35775;
    wire N__35766;
    wire N__35761;
    wire N__35760;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35720;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35704;
    wire N__35699;
    wire N__35694;
    wire N__35693;
    wire N__35690;
    wire N__35689;
    wire N__35688;
    wire N__35687;
    wire N__35686;
    wire N__35685;
    wire N__35684;
    wire N__35683;
    wire N__35682;
    wire N__35681;
    wire N__35674;
    wire N__35671;
    wire N__35668;
    wire N__35659;
    wire N__35654;
    wire N__35651;
    wire N__35642;
    wire N__35641;
    wire N__35640;
    wire N__35637;
    wire N__35636;
    wire N__35635;
    wire N__35634;
    wire N__35633;
    wire N__35632;
    wire N__35631;
    wire N__35630;
    wire N__35629;
    wire N__35628;
    wire N__35623;
    wire N__35616;
    wire N__35607;
    wire N__35604;
    wire N__35601;
    wire N__35594;
    wire N__35591;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35575;
    wire N__35570;
    wire N__35559;
    wire N__35558;
    wire N__35557;
    wire N__35550;
    wire N__35547;
    wire N__35536;
    wire N__35533;
    wire N__35524;
    wire N__35519;
    wire N__35518;
    wire N__35517;
    wire N__35516;
    wire N__35515;
    wire N__35512;
    wire N__35511;
    wire N__35510;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35502;
    wire N__35501;
    wire N__35500;
    wire N__35499;
    wire N__35496;
    wire N__35489;
    wire N__35486;
    wire N__35479;
    wire N__35478;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35466;
    wire N__35457;
    wire N__35454;
    wire N__35451;
    wire N__35450;
    wire N__35449;
    wire N__35448;
    wire N__35443;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35405;
    wire N__35402;
    wire N__35401;
    wire N__35398;
    wire N__35385;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35373;
    wire N__35368;
    wire N__35363;
    wire N__35358;
    wire N__35353;
    wire N__35350;
    wire N__35349;
    wire N__35348;
    wire N__35347;
    wire N__35346;
    wire N__35345;
    wire N__35344;
    wire N__35343;
    wire N__35342;
    wire N__35339;
    wire N__35330;
    wire N__35325;
    wire N__35322;
    wire N__35311;
    wire N__35306;
    wire N__35303;
    wire N__35296;
    wire N__35289;
    wire N__35284;
    wire N__35279;
    wire N__35270;
    wire N__35267;
    wire N__35262;
    wire N__35261;
    wire N__35260;
    wire N__35259;
    wire N__35258;
    wire N__35257;
    wire N__35256;
    wire N__35255;
    wire N__35252;
    wire N__35245;
    wire N__35242;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35220;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35196;
    wire N__35185;
    wire N__35178;
    wire N__35175;
    wire N__35170;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35145;
    wire N__35132;
    wire N__35129;
    wire N__35124;
    wire N__35103;
    wire N__35100;
    wire N__35099;
    wire N__35096;
    wire N__35093;
    wire N__35090;
    wire N__35087;
    wire N__35086;
    wire N__35081;
    wire N__35078;
    wire N__35073;
    wire N__35070;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35052;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35040;
    wire N__35039;
    wire N__35038;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35018;
    wire N__35015;
    wire N__35014;
    wire N__35013;
    wire N__35012;
    wire N__35009;
    wire N__35008;
    wire N__35007;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34993;
    wire N__34988;
    wire N__34983;
    wire N__34974;
    wire N__34971;
    wire N__34970;
    wire N__34969;
    wire N__34968;
    wire N__34963;
    wire N__34962;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34945;
    wire N__34940;
    wire N__34937;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34835;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34812;
    wire N__34809;
    wire N__34808;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34706;
    wire N__34705;
    wire N__34702;
    wire N__34697;
    wire N__34696;
    wire N__34695;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34683;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34671;
    wire N__34668;
    wire N__34659;
    wire N__34658;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34650;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34642;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34626;
    wire N__34621;
    wire N__34618;
    wire N__34613;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34554;
    wire N__34551;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34532;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34521;
    wire N__34520;
    wire N__34519;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34500;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34478;
    wire N__34477;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34461;
    wire N__34458;
    wire N__34457;
    wire N__34454;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34444;
    wire N__34439;
    wire N__34436;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34419;
    wire N__34412;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34402;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34382;
    wire N__34381;
    wire N__34380;
    wire N__34379;
    wire N__34376;
    wire N__34375;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34342;
    wire N__34339;
    wire N__34332;
    wire N__34331;
    wire N__34330;
    wire N__34329;
    wire N__34328;
    wire N__34327;
    wire N__34326;
    wire N__34325;
    wire N__34324;
    wire N__34323;
    wire N__34322;
    wire N__34321;
    wire N__34320;
    wire N__34319;
    wire N__34316;
    wire N__34309;
    wire N__34304;
    wire N__34303;
    wire N__34302;
    wire N__34301;
    wire N__34296;
    wire N__34291;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34279;
    wire N__34278;
    wire N__34271;
    wire N__34270;
    wire N__34269;
    wire N__34262;
    wire N__34257;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34226;
    wire N__34223;
    wire N__34212;
    wire N__34211;
    wire N__34208;
    wire N__34207;
    wire N__34206;
    wire N__34205;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34197;
    wire N__34188;
    wire N__34187;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34173;
    wire N__34172;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34155;
    wire N__34148;
    wire N__34145;
    wire N__34134;
    wire N__34133;
    wire N__34132;
    wire N__34131;
    wire N__34130;
    wire N__34123;
    wire N__34118;
    wire N__34117;
    wire N__34116;
    wire N__34115;
    wire N__34114;
    wire N__34109;
    wire N__34108;
    wire N__34105;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34083;
    wire N__34080;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34072;
    wire N__34071;
    wire N__34070;
    wire N__34069;
    wire N__34068;
    wire N__34067;
    wire N__34066;
    wire N__34061;
    wire N__34060;
    wire N__34059;
    wire N__34058;
    wire N__34057;
    wire N__34050;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34036;
    wire N__34031;
    wire N__34026;
    wire N__34023;
    wire N__34018;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34003;
    wire N__34000;
    wire N__33997;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33971;
    wire N__33968;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33951;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33894;
    wire N__33893;
    wire N__33892;
    wire N__33889;
    wire N__33888;
    wire N__33885;
    wire N__33884;
    wire N__33883;
    wire N__33878;
    wire N__33873;
    wire N__33870;
    wire N__33869;
    wire N__33868;
    wire N__33865;
    wire N__33862;
    wire N__33859;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33843;
    wire N__33834;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33798;
    wire N__33795;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33782;
    wire N__33781;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33740;
    wire N__33739;
    wire N__33738;
    wire N__33737;
    wire N__33736;
    wire N__33733;
    wire N__33724;
    wire N__33723;
    wire N__33722;
    wire N__33719;
    wire N__33714;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33701;
    wire N__33698;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33675;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33665;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33657;
    wire N__33656;
    wire N__33655;
    wire N__33652;
    wire N__33647;
    wire N__33640;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33611;
    wire N__33610;
    wire N__33609;
    wire N__33606;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33572;
    wire N__33571;
    wire N__33570;
    wire N__33563;
    wire N__33558;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33544;
    wire N__33541;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33524;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33491;
    wire N__33490;
    wire N__33489;
    wire N__33488;
    wire N__33483;
    wire N__33476;
    wire N__33471;
    wire N__33468;
    wire N__33467;
    wire N__33466;
    wire N__33461;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33438;
    wire N__33437;
    wire N__33436;
    wire N__33433;
    wire N__33432;
    wire N__33429;
    wire N__33422;
    wire N__33417;
    wire N__33416;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33363;
    wire N__33360;
    wire N__33357;
    wire N__33356;
    wire N__33351;
    wire N__33348;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33332;
    wire N__33329;
    wire N__33326;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33312;
    wire N__33309;
    wire N__33306;
    wire N__33303;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33291;
    wire N__33290;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33275;
    wire N__33274;
    wire N__33273;
    wire N__33272;
    wire N__33271;
    wire N__33270;
    wire N__33269;
    wire N__33268;
    wire N__33267;
    wire N__33264;
    wire N__33263;
    wire N__33262;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33254;
    wire N__33253;
    wire N__33252;
    wire N__33251;
    wire N__33250;
    wire N__33247;
    wire N__33246;
    wire N__33245;
    wire N__33244;
    wire N__33243;
    wire N__33242;
    wire N__33241;
    wire N__33240;
    wire N__33239;
    wire N__33238;
    wire N__33235;
    wire N__33234;
    wire N__33233;
    wire N__33232;
    wire N__33231;
    wire N__33230;
    wire N__33229;
    wire N__33228;
    wire N__33227;
    wire N__33220;
    wire N__33219;
    wire N__33218;
    wire N__33217;
    wire N__33212;
    wire N__33203;
    wire N__33198;
    wire N__33191;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33176;
    wire N__33175;
    wire N__33174;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33166;
    wire N__33165;
    wire N__33164;
    wire N__33163;
    wire N__33160;
    wire N__33159;
    wire N__33158;
    wire N__33157;
    wire N__33156;
    wire N__33155;
    wire N__33154;
    wire N__33153;
    wire N__33144;
    wire N__33139;
    wire N__33138;
    wire N__33137;
    wire N__33136;
    wire N__33135;
    wire N__33132;
    wire N__33131;
    wire N__33130;
    wire N__33129;
    wire N__33126;
    wire N__33125;
    wire N__33124;
    wire N__33123;
    wire N__33122;
    wire N__33121;
    wire N__33120;
    wire N__33119;
    wire N__33118;
    wire N__33117;
    wire N__33112;
    wire N__33109;
    wire N__33108;
    wire N__33107;
    wire N__33106;
    wire N__33105;
    wire N__33104;
    wire N__33103;
    wire N__33102;
    wire N__33099;
    wire N__33098;
    wire N__33097;
    wire N__33096;
    wire N__33095;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33087;
    wire N__33086;
    wire N__33085;
    wire N__33084;
    wire N__33083;
    wire N__33082;
    wire N__33081;
    wire N__33078;
    wire N__33077;
    wire N__33076;
    wire N__33075;
    wire N__33074;
    wire N__33071;
    wire N__33070;
    wire N__33069;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33055;
    wire N__33050;
    wire N__33047;
    wire N__33038;
    wire N__33027;
    wire N__33026;
    wire N__33015;
    wire N__33010;
    wire N__33007;
    wire N__33006;
    wire N__33005;
    wire N__33000;
    wire N__32995;
    wire N__32994;
    wire N__32993;
    wire N__32992;
    wire N__32991;
    wire N__32990;
    wire N__32989;
    wire N__32988;
    wire N__32987;
    wire N__32986;
    wire N__32985;
    wire N__32984;
    wire N__32983;
    wire N__32982;
    wire N__32979;
    wire N__32978;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32970;
    wire N__32969;
    wire N__32958;
    wire N__32953;
    wire N__32944;
    wire N__32935;
    wire N__32932;
    wire N__32925;
    wire N__32920;
    wire N__32917;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32905;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32881;
    wire N__32878;
    wire N__32875;
    wire N__32870;
    wire N__32869;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32861;
    wire N__32860;
    wire N__32853;
    wire N__32848;
    wire N__32847;
    wire N__32846;
    wire N__32843;
    wire N__32840;
    wire N__32839;
    wire N__32838;
    wire N__32835;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32813;
    wire N__32808;
    wire N__32807;
    wire N__32806;
    wire N__32805;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32784;
    wire N__32781;
    wire N__32780;
    wire N__32779;
    wire N__32778;
    wire N__32777;
    wire N__32774;
    wire N__32773;
    wire N__32770;
    wire N__32769;
    wire N__32768;
    wire N__32767;
    wire N__32764;
    wire N__32763;
    wire N__32762;
    wire N__32761;
    wire N__32760;
    wire N__32759;
    wire N__32758;
    wire N__32757;
    wire N__32756;
    wire N__32747;
    wire N__32744;
    wire N__32739;
    wire N__32734;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32718;
    wire N__32709;
    wire N__32706;
    wire N__32705;
    wire N__32704;
    wire N__32695;
    wire N__32690;
    wire N__32681;
    wire N__32676;
    wire N__32671;
    wire N__32666;
    wire N__32661;
    wire N__32656;
    wire N__32649;
    wire N__32644;
    wire N__32643;
    wire N__32640;
    wire N__32639;
    wire N__32638;
    wire N__32637;
    wire N__32632;
    wire N__32623;
    wire N__32614;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32591;
    wire N__32590;
    wire N__32589;
    wire N__32588;
    wire N__32587;
    wire N__32582;
    wire N__32575;
    wire N__32572;
    wire N__32563;
    wire N__32554;
    wire N__32549;
    wire N__32542;
    wire N__32531;
    wire N__32528;
    wire N__32521;
    wire N__32516;
    wire N__32505;
    wire N__32502;
    wire N__32497;
    wire N__32494;
    wire N__32485;
    wire N__32480;
    wire N__32475;
    wire N__32474;
    wire N__32469;
    wire N__32462;
    wire N__32459;
    wire N__32454;
    wire N__32449;
    wire N__32444;
    wire N__32439;
    wire N__32438;
    wire N__32437;
    wire N__32434;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32380;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32372;
    wire N__32363;
    wire N__32354;
    wire N__32351;
    wire N__32348;
    wire N__32343;
    wire N__32340;
    wire N__32333;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32321;
    wire N__32304;
    wire N__32303;
    wire N__32300;
    wire N__32297;
    wire N__32296;
    wire N__32295;
    wire N__32294;
    wire N__32293;
    wire N__32292;
    wire N__32291;
    wire N__32290;
    wire N__32289;
    wire N__32288;
    wire N__32287;
    wire N__32286;
    wire N__32285;
    wire N__32284;
    wire N__32283;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32268;
    wire N__32265;
    wire N__32258;
    wire N__32251;
    wire N__32246;
    wire N__32245;
    wire N__32244;
    wire N__32243;
    wire N__32242;
    wire N__32241;
    wire N__32240;
    wire N__32239;
    wire N__32238;
    wire N__32237;
    wire N__32236;
    wire N__32235;
    wire N__32234;
    wire N__32233;
    wire N__32232;
    wire N__32231;
    wire N__32230;
    wire N__32229;
    wire N__32228;
    wire N__32227;
    wire N__32226;
    wire N__32223;
    wire N__32222;
    wire N__32221;
    wire N__32220;
    wire N__32219;
    wire N__32218;
    wire N__32217;
    wire N__32216;
    wire N__32213;
    wire N__32212;
    wire N__32211;
    wire N__32208;
    wire N__32207;
    wire N__32206;
    wire N__32205;
    wire N__32204;
    wire N__32203;
    wire N__32202;
    wire N__32201;
    wire N__32184;
    wire N__32179;
    wire N__32174;
    wire N__32173;
    wire N__32172;
    wire N__32171;
    wire N__32170;
    wire N__32169;
    wire N__32166;
    wire N__32165;
    wire N__32164;
    wire N__32163;
    wire N__32162;
    wire N__32161;
    wire N__32160;
    wire N__32157;
    wire N__32148;
    wire N__32145;
    wire N__32144;
    wire N__32143;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32135;
    wire N__32134;
    wire N__32133;
    wire N__32132;
    wire N__32131;
    wire N__32130;
    wire N__32129;
    wire N__32128;
    wire N__32127;
    wire N__32126;
    wire N__32125;
    wire N__32124;
    wire N__32123;
    wire N__32122;
    wire N__32117;
    wire N__32112;
    wire N__32111;
    wire N__32106;
    wire N__32101;
    wire N__32100;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32092;
    wire N__32091;
    wire N__32090;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32086;
    wire N__32085;
    wire N__32084;
    wire N__32077;
    wire N__32076;
    wire N__32073;
    wire N__32072;
    wire N__32071;
    wire N__32070;
    wire N__32069;
    wire N__32068;
    wire N__32067;
    wire N__32066;
    wire N__32065;
    wire N__32064;
    wire N__32063;
    wire N__32060;
    wire N__32059;
    wire N__32058;
    wire N__32057;
    wire N__32056;
    wire N__32055;
    wire N__32054;
    wire N__32053;
    wire N__32052;
    wire N__32049;
    wire N__32044;
    wire N__32039;
    wire N__32030;
    wire N__32025;
    wire N__32024;
    wire N__32021;
    wire N__32016;
    wire N__32011;
    wire N__32008;
    wire N__32007;
    wire N__32006;
    wire N__32005;
    wire N__32004;
    wire N__32001;
    wire N__32000;
    wire N__31999;
    wire N__31998;
    wire N__31997;
    wire N__31996;
    wire N__31995;
    wire N__31994;
    wire N__31991;
    wire N__31986;
    wire N__31975;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31958;
    wire N__31953;
    wire N__31948;
    wire N__31945;
    wire N__31944;
    wire N__31943;
    wire N__31942;
    wire N__31941;
    wire N__31940;
    wire N__31939;
    wire N__31938;
    wire N__31937;
    wire N__31936;
    wire N__31933;
    wire N__31932;
    wire N__31931;
    wire N__31930;
    wire N__31927;
    wire N__31924;
    wire N__31919;
    wire N__31916;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31901;
    wire N__31896;
    wire N__31893;
    wire N__31888;
    wire N__31887;
    wire N__31884;
    wire N__31883;
    wire N__31882;
    wire N__31877;
    wire N__31868;
    wire N__31863;
    wire N__31854;
    wire N__31851;
    wire N__31850;
    wire N__31849;
    wire N__31848;
    wire N__31847;
    wire N__31846;
    wire N__31845;
    wire N__31840;
    wire N__31835;
    wire N__31830;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31804;
    wire N__31795;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31772;
    wire N__31769;
    wire N__31762;
    wire N__31751;
    wire N__31746;
    wire N__31741;
    wire N__31734;
    wire N__31721;
    wire N__31716;
    wire N__31715;
    wire N__31714;
    wire N__31713;
    wire N__31712;
    wire N__31711;
    wire N__31710;
    wire N__31709;
    wire N__31708;
    wire N__31707;
    wire N__31706;
    wire N__31705;
    wire N__31704;
    wire N__31701;
    wire N__31700;
    wire N__31699;
    wire N__31694;
    wire N__31689;
    wire N__31680;
    wire N__31671;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31651;
    wire N__31646;
    wire N__31641;
    wire N__31632;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31606;
    wire N__31595;
    wire N__31592;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31551;
    wire N__31548;
    wire N__31541;
    wire N__31530;
    wire N__31521;
    wire N__31512;
    wire N__31509;
    wire N__31498;
    wire N__31493;
    wire N__31482;
    wire N__31479;
    wire N__31468;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31436;
    wire N__31433;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31416;
    wire N__31413;
    wire N__31412;
    wire N__31411;
    wire N__31408;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31368;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31357;
    wire N__31354;
    wire N__31351;
    wire N__31348;
    wire N__31341;
    wire N__31338;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31326;
    wire N__31323;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31311;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31298;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31281;
    wire N__31278;
    wire N__31277;
    wire N__31276;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31210;
    wire N__31205;
    wire N__31202;
    wire N__31197;
    wire N__31194;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31184;
    wire N__31183;
    wire N__31178;
    wire N__31175;
    wire N__31170;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31144;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31130;
    wire N__31127;
    wire N__31126;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31114;
    wire N__31111;
    wire N__31104;
    wire N__31103;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31089;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31045;
    wire N__31040;
    wire N__31037;
    wire N__31032;
    wire N__31031;
    wire N__31028;
    wire N__31027;
    wire N__31024;
    wire N__31019;
    wire N__31014;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31001;
    wire N__31000;
    wire N__30997;
    wire N__30994;
    wire N__30993;
    wire N__30990;
    wire N__30985;
    wire N__30982;
    wire N__30975;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30967;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30936;
    wire N__30935;
    wire N__30934;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30917;
    wire N__30912;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30896;
    wire N__30893;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30882;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30858;
    wire N__30855;
    wire N__30846;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30833;
    wire N__30830;
    wire N__30829;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30780;
    wire N__30779;
    wire N__30776;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30735;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30695;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30629;
    wire N__30628;
    wire N__30625;
    wire N__30620;
    wire N__30615;
    wire N__30614;
    wire N__30611;
    wire N__30608;
    wire N__30607;
    wire N__30606;
    wire N__30605;
    wire N__30600;
    wire N__30597;
    wire N__30594;
    wire N__30593;
    wire N__30590;
    wire N__30585;
    wire N__30580;
    wire N__30573;
    wire N__30570;
    wire N__30569;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30561;
    wire N__30560;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30534;
    wire N__30531;
    wire N__30530;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30522;
    wire N__30519;
    wire N__30518;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30498;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30453;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30439;
    wire N__30434;
    wire N__30431;
    wire N__30428;
    wire N__30423;
    wire N__30420;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30390;
    wire N__30387;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30341;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30308;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30291;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30280;
    wire N__30277;
    wire N__30274;
    wire N__30271;
    wire N__30264;
    wire N__30261;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30230;
    wire N__30225;
    wire N__30220;
    wire N__30217;
    wire N__30210;
    wire N__30209;
    wire N__30208;
    wire N__30207;
    wire N__30206;
    wire N__30205;
    wire N__30204;
    wire N__30201;
    wire N__30200;
    wire N__30199;
    wire N__30198;
    wire N__30195;
    wire N__30194;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30186;
    wire N__30185;
    wire N__30184;
    wire N__30181;
    wire N__30180;
    wire N__30177;
    wire N__30176;
    wire N__30175;
    wire N__30174;
    wire N__30173;
    wire N__30172;
    wire N__30171;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30154;
    wire N__30153;
    wire N__30150;
    wire N__30149;
    wire N__30148;
    wire N__30147;
    wire N__30146;
    wire N__30145;
    wire N__30144;
    wire N__30141;
    wire N__30136;
    wire N__30133;
    wire N__30132;
    wire N__30129;
    wire N__30128;
    wire N__30127;
    wire N__30126;
    wire N__30125;
    wire N__30122;
    wire N__30121;
    wire N__30114;
    wire N__30113;
    wire N__30112;
    wire N__30111;
    wire N__30110;
    wire N__30109;
    wire N__30106;
    wire N__30105;
    wire N__30102;
    wire N__30101;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30093;
    wire N__30090;
    wire N__30089;
    wire N__30086;
    wire N__30081;
    wire N__30074;
    wire N__30071;
    wire N__30070;
    wire N__30069;
    wire N__30066;
    wire N__30065;
    wire N__30062;
    wire N__30061;
    wire N__30060;
    wire N__30059;
    wire N__30056;
    wire N__30055;
    wire N__30054;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30040;
    wire N__30035;
    wire N__30030;
    wire N__30029;
    wire N__30026;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30018;
    wire N__30017;
    wire N__30016;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29999;
    wire N__29994;
    wire N__29989;
    wire N__29986;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29971;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29949;
    wire N__29948;
    wire N__29947;
    wire N__29944;
    wire N__29943;
    wire N__29940;
    wire N__29939;
    wire N__29938;
    wire N__29935;
    wire N__29930;
    wire N__29929;
    wire N__29926;
    wire N__29925;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29911;
    wire N__29908;
    wire N__29897;
    wire N__29892;
    wire N__29883;
    wire N__29878;
    wire N__29875;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29857;
    wire N__29854;
    wire N__29847;
    wire N__29842;
    wire N__29839;
    wire N__29828;
    wire N__29827;
    wire N__29826;
    wire N__29825;
    wire N__29824;
    wire N__29823;
    wire N__29818;
    wire N__29813;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29803;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29792;
    wire N__29787;
    wire N__29786;
    wire N__29783;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29765;
    wire N__29752;
    wire N__29745;
    wire N__29742;
    wire N__29735;
    wire N__29732;
    wire N__29723;
    wire N__29718;
    wire N__29713;
    wire N__29710;
    wire N__29703;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29675;
    wire N__29668;
    wire N__29661;
    wire N__29646;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29612;
    wire N__29609;
    wire N__29608;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29558;
    wire N__29555;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29514;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29484;
    wire N__29483;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29469;
    wire N__29460;
    wire N__29459;
    wire N__29458;
    wire N__29455;
    wire N__29450;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29412;
    wire N__29409;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29354;
    wire N__29349;
    wire N__29346;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29334;
    wire N__29333;
    wire N__29328;
    wire N__29327;
    wire N__29326;
    wire N__29325;
    wire N__29322;
    wire N__29321;
    wire N__29318;
    wire N__29317;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29286;
    wire N__29283;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29268;
    wire N__29265;
    wire N__29264;
    wire N__29261;
    wire N__29258;
    wire N__29253;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29239;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29204;
    wire N__29203;
    wire N__29202;
    wire N__29201;
    wire N__29200;
    wire N__29199;
    wire N__29198;
    wire N__29193;
    wire N__29190;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29175;
    wire N__29174;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29138;
    wire N__29135;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29117;
    wire N__29116;
    wire N__29115;
    wire N__29114;
    wire N__29113;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29101;
    wire N__29098;
    wire N__29093;
    wire N__29092;
    wire N__29091;
    wire N__29090;
    wire N__29089;
    wire N__29088;
    wire N__29087;
    wire N__29082;
    wire N__29079;
    wire N__29074;
    wire N__29071;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29045;
    wire N__29042;
    wire N__29025;
    wire N__29022;
    wire N__29021;
    wire N__29018;
    wire N__29017;
    wire N__29016;
    wire N__29015;
    wire N__29012;
    wire N__29011;
    wire N__29010;
    wire N__29009;
    wire N__29006;
    wire N__29005;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28993;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28979;
    wire N__28978;
    wire N__28977;
    wire N__28976;
    wire N__28975;
    wire N__28974;
    wire N__28973;
    wire N__28970;
    wire N__28969;
    wire N__28968;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28958;
    wire N__28957;
    wire N__28956;
    wire N__28949;
    wire N__28946;
    wire N__28937;
    wire N__28934;
    wire N__28925;
    wire N__28922;
    wire N__28917;
    wire N__28910;
    wire N__28907;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28883;
    wire N__28880;
    wire N__28877;
    wire N__28872;
    wire N__28869;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28857;
    wire N__28854;
    wire N__28851;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28841;
    wire N__28840;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28817;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28800;
    wire N__28799;
    wire N__28796;
    wire N__28793;
    wire N__28790;
    wire N__28787;
    wire N__28782;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28745;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28697;
    wire N__28692;
    wire N__28689;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28677;
    wire N__28674;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28647;
    wire N__28644;
    wire N__28641;
    wire N__28640;
    wire N__28639;
    wire N__28638;
    wire N__28637;
    wire N__28636;
    wire N__28629;
    wire N__28622;
    wire N__28617;
    wire N__28614;
    wire N__28613;
    wire N__28610;
    wire N__28609;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28598;
    wire N__28597;
    wire N__28594;
    wire N__28587;
    wire N__28584;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28567;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28533;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28518;
    wire N__28517;
    wire N__28514;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28496;
    wire N__28495;
    wire N__28490;
    wire N__28487;
    wire N__28486;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28478;
    wire N__28477;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28461;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28433;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28402;
    wire N__28395;
    wire N__28392;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28368;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28349;
    wire N__28348;
    wire N__28345;
    wire N__28340;
    wire N__28339;
    wire N__28338;
    wire N__28333;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28311;
    wire N__28310;
    wire N__28307;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28299;
    wire N__28296;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28281;
    wire N__28278;
    wire N__28277;
    wire N__28274;
    wire N__28271;
    wire N__28270;
    wire N__28267;
    wire N__28264;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28239;
    wire N__28238;
    wire N__28235;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28204;
    wire N__28197;
    wire N__28196;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28169;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28157;
    wire N__28152;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28130;
    wire N__28127;
    wire N__28126;
    wire N__28123;
    wire N__28122;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28100;
    wire N__28097;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28082;
    wire N__28079;
    wire N__28074;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28045;
    wire N__28044;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28032;
    wire N__28029;
    wire N__28020;
    wire N__28017;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28005;
    wire N__28002;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27987;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27960;
    wire N__27957;
    wire N__27954;
    wire N__27953;
    wire N__27952;
    wire N__27951;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27941;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27923;
    wire N__27916;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27861;
    wire N__27858;
    wire N__27857;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27819;
    wire N__27816;
    wire N__27815;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27795;
    wire N__27792;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27755;
    wire N__27754;
    wire N__27753;
    wire N__27750;
    wire N__27749;
    wire N__27748;
    wire N__27747;
    wire N__27746;
    wire N__27745;
    wire N__27744;
    wire N__27743;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27721;
    wire N__27720;
    wire N__27719;
    wire N__27718;
    wire N__27717;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27703;
    wire N__27702;
    wire N__27691;
    wire N__27688;
    wire N__27687;
    wire N__27686;
    wire N__27685;
    wire N__27684;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27667;
    wire N__27666;
    wire N__27665;
    wire N__27664;
    wire N__27663;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27648;
    wire N__27647;
    wire N__27646;
    wire N__27641;
    wire N__27636;
    wire N__27635;
    wire N__27634;
    wire N__27633;
    wire N__27632;
    wire N__27629;
    wire N__27624;
    wire N__27621;
    wire N__27614;
    wire N__27613;
    wire N__27612;
    wire N__27609;
    wire N__27608;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27574;
    wire N__27569;
    wire N__27568;
    wire N__27565;
    wire N__27558;
    wire N__27557;
    wire N__27554;
    wire N__27547;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27517;
    wire N__27514;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27490;
    wire N__27487;
    wire N__27482;
    wire N__27477;
    wire N__27470;
    wire N__27465;
    wire N__27444;
    wire N__27443;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27327;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27286;
    wire N__27285;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27271;
    wire N__27268;
    wire N__27261;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27243;
    wire N__27242;
    wire N__27241;
    wire N__27238;
    wire N__27235;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27181;
    wire N__27176;
    wire N__27173;
    wire N__27168;
    wire N__27165;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27157;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27145;
    wire N__27138;
    wire N__27137;
    wire N__27134;
    wire N__27133;
    wire N__27132;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27120;
    wire N__27115;
    wire N__27112;
    wire N__27109;
    wire N__27104;
    wire N__27099;
    wire N__27098;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27071;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27053;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27007;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26991;
    wire N__26990;
    wire N__26987;
    wire N__26986;
    wire N__26983;
    wire N__26982;
    wire N__26979;
    wire N__26974;
    wire N__26971;
    wire N__26964;
    wire N__26961;
    wire N__26960;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26952;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26937;
    wire N__26934;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26918;
    wire N__26917;
    wire N__26914;
    wire N__26909;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26890;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26878;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26866;
    wire N__26859;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26829;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26814;
    wire N__26805;
    wire N__26802;
    wire N__26801;
    wire N__26800;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26766;
    wire N__26763;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26700;
    wire N__26697;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26676;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26649;
    wire N__26646;
    wire N__26645;
    wire N__26644;
    wire N__26643;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26613;
    wire N__26612;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26600;
    wire N__26595;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26579;
    wire N__26576;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26561;
    wire N__26558;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26538;
    wire N__26537;
    wire N__26534;
    wire N__26533;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26495;
    wire N__26494;
    wire N__26493;
    wire N__26490;
    wire N__26485;
    wire N__26482;
    wire N__26475;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26460;
    wire N__26459;
    wire N__26458;
    wire N__26457;
    wire N__26456;
    wire N__26451;
    wire N__26446;
    wire N__26443;
    wire N__26436;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26424;
    wire N__26421;
    wire N__26418;
    wire N__26417;
    wire N__26414;
    wire N__26413;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26400;
    wire N__26391;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26353;
    wire N__26350;
    wire N__26347;
    wire N__26344;
    wire N__26337;
    wire N__26334;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26322;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26307;
    wire N__26304;
    wire N__26303;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26277;
    wire N__26274;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26262;
    wire N__26259;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26235;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26217;
    wire N__26214;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26195;
    wire N__26192;
    wire N__26187;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26162;
    wire N__26159;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26123;
    wire N__26120;
    wire N__26117;
    wire N__26112;
    wire N__26111;
    wire N__26106;
    wire N__26103;
    wire N__26100;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26085;
    wire N__26082;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26067;
    wire N__26064;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26025;
    wire N__26022;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26007;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25995;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25984;
    wire N__25983;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25962;
    wire N__25959;
    wire N__25950;
    wire N__25947;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25936;
    wire N__25935;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25921;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25905;
    wire N__25902;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25894;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25869;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25821;
    wire N__25818;
    wire N__25813;
    wire N__25810;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25794;
    wire N__25793;
    wire N__25790;
    wire N__25789;
    wire N__25788;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25776;
    wire N__25773;
    wire N__25764;
    wire N__25761;
    wire N__25760;
    wire N__25757;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25716;
    wire N__25715;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25695;
    wire N__25692;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25674;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25662;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25647;
    wire N__25644;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25629;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25599;
    wire N__25596;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25584;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25572;
    wire N__25569;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25555;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25543;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25531;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25500;
    wire N__25497;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25463;
    wire N__25462;
    wire N__25459;
    wire N__25456;
    wire N__25455;
    wire N__25454;
    wire N__25451;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25430;
    wire N__25427;
    wire N__25422;
    wire N__25413;
    wire N__25410;
    wire N__25409;
    wire N__25408;
    wire N__25407;
    wire N__25406;
    wire N__25405;
    wire N__25404;
    wire N__25403;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25392;
    wire N__25391;
    wire N__25390;
    wire N__25387;
    wire N__25386;
    wire N__25383;
    wire N__25382;
    wire N__25381;
    wire N__25376;
    wire N__25373;
    wire N__25372;
    wire N__25369;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25316;
    wire N__25307;
    wire N__25306;
    wire N__25305;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25269;
    wire N__25260;
    wire N__25259;
    wire N__25258;
    wire N__25257;
    wire N__25256;
    wire N__25253;
    wire N__25252;
    wire N__25249;
    wire N__25248;
    wire N__25247;
    wire N__25244;
    wire N__25239;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25190;
    wire N__25185;
    wire N__25182;
    wire N__25173;
    wire N__25170;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25148;
    wire N__25145;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25134;
    wire N__25131;
    wire N__25126;
    wire N__25123;
    wire N__25118;
    wire N__25113;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25105;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25045;
    wire N__25044;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25026;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25018;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25006;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24983;
    wire N__24982;
    wire N__24979;
    wire N__24974;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24959;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24890;
    wire N__24887;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24870;
    wire N__24869;
    wire N__24868;
    wire N__24865;
    wire N__24862;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24819;
    wire N__24816;
    wire N__24807;
    wire N__24806;
    wire N__24803;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24782;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24750;
    wire N__24747;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24605;
    wire N__24604;
    wire N__24603;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24569;
    wire N__24566;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24529;
    wire N__24528;
    wire N__24527;
    wire N__24522;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24369;
    wire N__24366;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24345;
    wire N__24344;
    wire N__24339;
    wire N__24336;
    wire N__24331;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24317;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24264;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24210;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24180;
    wire N__24177;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24134;
    wire N__24131;
    wire N__24128;
    wire N__24123;
    wire N__24120;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24099;
    wire N__24098;
    wire N__24097;
    wire N__24096;
    wire N__24093;
    wire N__24086;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24068;
    wire N__24067;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24055;
    wire N__24052;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24038;
    wire N__24037;
    wire N__24034;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23985;
    wire N__23984;
    wire N__23981;
    wire N__23980;
    wire N__23979;
    wire N__23978;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23930;
    wire N__23929;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23917;
    wire N__23910;
    wire N__23907;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23890;
    wire N__23885;
    wire N__23882;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23835;
    wire N__23832;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23817;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23780;
    wire N__23779;
    wire N__23778;
    wire N__23775;
    wire N__23768;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23677;
    wire N__23676;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23662;
    wire N__23655;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23622;
    wire N__23619;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23562;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23550;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23535;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23510;
    wire N__23509;
    wire N__23506;
    wire N__23501;
    wire N__23496;
    wire N__23493;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23457;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23414;
    wire N__23413;
    wire N__23410;
    wire N__23405;
    wire N__23400;
    wire N__23397;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23354;
    wire N__23353;
    wire N__23350;
    wire N__23345;
    wire N__23340;
    wire N__23339;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23310;
    wire N__23307;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23299;
    wire N__23298;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23284;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23238;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23227;
    wire N__23222;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23181;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23157;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23116;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23048;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23025;
    wire N__23022;
    wire N__23021;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22986;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22967;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22916;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22896;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22813;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22801;
    wire N__22794;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22674;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22650;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22642;
    wire N__22639;
    wire N__22638;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22608;
    wire N__22605;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22593;
    wire N__22590;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22575;
    wire N__22574;
    wire N__22571;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22531;
    wire N__22530;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22515;
    wire N__22506;
    wire N__22503;
    wire N__22502;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22485;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22464;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22439;
    wire N__22438;
    wire N__22435;
    wire N__22430;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22415;
    wire N__22414;
    wire N__22411;
    wire N__22406;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22364;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22350;
    wire N__22347;
    wire N__22346;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22328;
    wire N__22317;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22309;
    wire N__22304;
    wire N__22301;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22278;
    wire N__22275;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22228;
    wire N__22223;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22206;
    wire N__22203;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22189;
    wire N__22188;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22170;
    wire N__22167;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22092;
    wire N__22091;
    wire N__22088;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22077;
    wire N__22074;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22056;
    wire N__22055;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22027;
    wire N__22020;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22006;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21984;
    wire N__21983;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21975;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21945;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21914;
    wire N__21911;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21896;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21881;
    wire N__21876;
    wire N__21873;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21853;
    wire N__21848;
    wire N__21845;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21809;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21798;
    wire N__21797;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21771;
    wire N__21770;
    wire N__21769;
    wire N__21766;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21698;
    wire N__21697;
    wire N__21694;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21669;
    wire N__21666;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21624;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21597;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21585;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21573;
    wire N__21572;
    wire N__21569;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21543;
    wire N__21540;
    wire N__21539;
    wire N__21538;
    wire N__21537;
    wire N__21534;
    wire N__21529;
    wire N__21528;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21513;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21413;
    wire N__21412;
    wire N__21409;
    wire N__21404;
    wire N__21399;
    wire N__21396;
    wire N__21395;
    wire N__21392;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21361;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21308;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21241;
    wire N__21236;
    wire N__21233;
    wire N__21228;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21211;
    wire N__21210;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21195;
    wire N__21192;
    wire N__21183;
    wire N__21180;
    wire N__21179;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21164;
    wire N__21161;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21128;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21101;
    wire N__21100;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21088;
    wire N__21081;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21056;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21033;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21003;
    wire N__21002;
    wire N__21001;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20978;
    wire N__20977;
    wire N__20968;
    wire N__20963;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20951;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20943;
    wire N__20940;
    wire N__20935;
    wire N__20932;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20892;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20858;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20847;
    wire N__20844;
    wire N__20843;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20825;
    wire N__20818;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20780;
    wire N__20777;
    wire N__20770;
    wire N__20767;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20741;
    wire N__20740;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20714;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20702;
    wire N__20697;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20657;
    wire N__20654;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20626;
    wire N__20619;
    wire N__20616;
    wire N__20615;
    wire N__20614;
    wire N__20613;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20593;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20559;
    wire N__20556;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20544;
    wire N__20543;
    wire N__20542;
    wire N__20541;
    wire N__20538;
    wire N__20533;
    wire N__20530;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20499;
    wire N__20496;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20417;
    wire N__20416;
    wire N__20413;
    wire N__20412;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20404;
    wire N__20403;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20364;
    wire N__20363;
    wire N__20362;
    wire N__20361;
    wire N__20360;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20349;
    wire N__20346;
    wire N__20345;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20330;
    wire N__20327;
    wire N__20320;
    wire N__20317;
    wire N__20316;
    wire N__20313;
    wire N__20304;
    wire N__20301;
    wire N__20300;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20265;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20236;
    wire N__20235;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20201;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20164;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20150;
    wire N__20147;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20129;
    wire N__20124;
    wire N__20123;
    wire N__20122;
    wire N__20119;
    wire N__20118;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20102;
    wire N__20097;
    wire N__20094;
    wire N__20093;
    wire N__20092;
    wire N__20089;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20073;
    wire N__20070;
    wire N__20067;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20045;
    wire N__20044;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20033;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20015;
    wire N__20004;
    wire N__20001;
    wire N__20000;
    wire N__19999;
    wire N__19998;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19990;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19969;
    wire N__19956;
    wire N__19953;
    wire N__19952;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19898;
    wire N__19897;
    wire N__19894;
    wire N__19889;
    wire N__19884;
    wire N__19881;
    wire N__19880;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19869;
    wire N__19864;
    wire N__19861;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19818;
    wire N__19815;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19791;
    wire N__19790;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19731;
    wire N__19730;
    wire N__19729;
    wire N__19726;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19688;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19671;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19641;
    wire N__19640;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19617;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19602;
    wire N__19593;
    wire N__19590;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19575;
    wire N__19572;
    wire N__19567;
    wire N__19564;
    wire N__19557;
    wire N__19554;
    wire N__19553;
    wire N__19550;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19533;
    wire N__19530;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19503;
    wire N__19500;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19486;
    wire N__19481;
    wire N__19478;
    wire N__19473;
    wire N__19470;
    wire N__19469;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19450;
    wire N__19443;
    wire N__19440;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19406;
    wire N__19405;
    wire N__19402;
    wire N__19397;
    wire N__19392;
    wire N__19389;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19377;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19337;
    wire N__19336;
    wire N__19333;
    wire N__19328;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19294;
    wire N__19289;
    wire N__19286;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19274;
    wire N__19273;
    wire N__19270;
    wire N__19265;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19235;
    wire N__19234;
    wire N__19233;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19219;
    wire N__19212;
    wire N__19209;
    wire N__19208;
    wire N__19207;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19192;
    wire N__19191;
    wire N__19190;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19171;
    wire N__19164;
    wire N__19163;
    wire N__19160;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19136;
    wire N__19133;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19106;
    wire N__19105;
    wire N__19102;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19084;
    wire N__19077;
    wire N__19074;
    wire N__19071;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19043;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19026;
    wire N__19023;
    wire N__19022;
    wire N__19021;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire N__18990;
    wire N__18987;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18977;
    wire N__18976;
    wire N__18973;
    wire N__18968;
    wire N__18963;
    wire N__18962;
    wire N__18959;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18945;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18930;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18914;
    wire N__18911;
    wire N__18910;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18898;
    wire N__18895;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18881;
    wire N__18878;
    wire N__18877;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18855;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18841;
    wire N__18836;
    wire N__18833;
    wire N__18828;
    wire N__18825;
    wire N__18824;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18813;
    wire N__18812;
    wire N__18809;
    wire N__18804;
    wire N__18799;
    wire N__18792;
    wire N__18791;
    wire N__18790;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18763;
    wire N__18758;
    wire N__18755;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18726;
    wire N__18719;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18695;
    wire N__18694;
    wire N__18691;
    wire N__18686;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18671;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18654;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18646;
    wire N__18641;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18624;
    wire N__18621;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18609;
    wire N__18606;
    wire N__18605;
    wire N__18602;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18578;
    wire N__18577;
    wire N__18574;
    wire N__18573;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18552;
    wire N__18547;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18509;
    wire N__18508;
    wire N__18505;
    wire N__18500;
    wire N__18495;
    wire N__18492;
    wire N__18489;
    wire N__18488;
    wire N__18487;
    wire N__18484;
    wire N__18479;
    wire N__18474;
    wire N__18471;
    wire N__18470;
    wire N__18467;
    wire N__18466;
    wire N__18465;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18441;
    wire N__18432;
    wire N__18431;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18403;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18381;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18358;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18346;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18329;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18312;
    wire N__18309;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18290;
    wire N__18287;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18262;
    wire N__18259;
    wire N__18252;
    wire N__18249;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18237;
    wire N__18236;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18212;
    wire N__18211;
    wire N__18208;
    wire N__18203;
    wire N__18198;
    wire N__18195;
    wire N__18194;
    wire N__18193;
    wire N__18190;
    wire N__18187;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18171;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18152;
    wire N__18151;
    wire N__18150;
    wire N__18147;
    wire N__18140;
    wire N__18135;
    wire N__18134;
    wire N__18133;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18121;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18105;
    wire N__18104;
    wire N__18101;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18089;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18039;
    wire N__18036;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18024;
    wire N__18023;
    wire N__18022;
    wire N__18019;
    wire N__18018;
    wire N__18017;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18007;
    wire N__18006;
    wire N__18005;
    wire N__18004;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17996;
    wire N__17993;
    wire N__17992;
    wire N__17987;
    wire N__17984;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17967;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17953;
    wire N__17946;
    wire N__17931;
    wire N__17928;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17914;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17898;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17880;
    wire N__17877;
    wire N__17874;
    wire N__17871;
    wire N__17870;
    wire N__17869;
    wire N__17866;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17851;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17837;
    wire N__17836;
    wire N__17833;
    wire N__17828;
    wire N__17825;
    wire N__17820;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17805;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17783;
    wire N__17782;
    wire N__17779;
    wire N__17774;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17760;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17748;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17730;
    wire N__17727;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17709;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17697;
    wire N__17696;
    wire N__17695;
    wire N__17692;
    wire N__17691;
    wire N__17690;
    wire N__17689;
    wire N__17688;
    wire N__17685;
    wire N__17684;
    wire N__17683;
    wire N__17680;
    wire N__17675;
    wire N__17670;
    wire N__17667;
    wire N__17660;
    wire N__17655;
    wire N__17646;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17638;
    wire N__17637;
    wire N__17636;
    wire N__17635;
    wire N__17634;
    wire N__17631;
    wire N__17630;
    wire N__17627;
    wire N__17622;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17589;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17577;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17566;
    wire N__17565;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17551;
    wire N__17544;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17517;
    wire N__17514;
    wire N__17511;
    wire N__17508;
    wire N__17505;
    wire N__17504;
    wire N__17501;
    wire N__17500;
    wire N__17499;
    wire N__17496;
    wire N__17493;
    wire N__17488;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17445;
    wire N__17442;
    wire N__17441;
    wire N__17440;
    wire N__17439;
    wire N__17436;
    wire N__17435;
    wire N__17432;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17418;
    wire N__17409;
    wire N__17406;
    wire N__17403;
    wire N__17400;
    wire N__17397;
    wire N__17394;
    wire N__17391;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17379;
    wire N__17376;
    wire N__17373;
    wire N__17372;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17355;
    wire N__17354;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17322;
    wire N__17319;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17311;
    wire N__17310;
    wire N__17309;
    wire N__17304;
    wire N__17301;
    wire N__17296;
    wire N__17289;
    wire N__17286;
    wire N__17285;
    wire N__17284;
    wire N__17283;
    wire N__17280;
    wire N__17277;
    wire N__17274;
    wire N__17273;
    wire N__17270;
    wire N__17265;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17248;
    wire N__17241;
    wire N__17238;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17223;
    wire N__17220;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17212;
    wire N__17211;
    wire N__17210;
    wire N__17209;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17187;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17166;
    wire N__17163;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17155;
    wire N__17154;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17140;
    wire N__17133;
    wire N__17130;
    wire N__17127;
    wire N__17126;
    wire N__17125;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17113;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17087;
    wire N__17086;
    wire N__17085;
    wire N__17082;
    wire N__17079;
    wire N__17076;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17058;
    wire N__17055;
    wire N__17052;
    wire N__17049;
    wire N__17046;
    wire N__17043;
    wire N__17040;
    wire N__17037;
    wire N__17034;
    wire N__17031;
    wire N__17028;
    wire N__17027;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17010;
    wire N__17007;
    wire N__17002;
    wire N__16999;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16971;
    wire N__16968;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16950;
    wire N__16947;
    wire N__16944;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16890;
    wire N__16887;
    wire N__16882;
    wire N__16879;
    wire N__16872;
    wire N__16869;
    wire N__16868;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16839;
    wire N__16836;
    wire N__16835;
    wire N__16830;
    wire N__16827;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16813;
    wire N__16812;
    wire N__16809;
    wire N__16806;
    wire N__16801;
    wire N__16794;
    wire N__16791;
    wire N__16790;
    wire N__16789;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16776;
    wire N__16771;
    wire N__16768;
    wire N__16767;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16752;
    wire N__16743;
    wire N__16740;
    wire N__16737;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16713;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16695;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16680;
    wire N__16677;
    wire N__16674;
    wire N__16671;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16646;
    wire N__16645;
    wire N__16642;
    wire N__16641;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16599;
    wire N__16598;
    wire N__16595;
    wire N__16594;
    wire N__16591;
    wire N__16588;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16575;
    wire N__16566;
    wire N__16565;
    wire N__16562;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16512;
    wire N__16511;
    wire N__16510;
    wire N__16507;
    wire N__16502;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16490;
    wire N__16489;
    wire N__16488;
    wire N__16485;
    wire N__16478;
    wire N__16473;
    wire N__16470;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16446;
    wire N__16445;
    wire N__16444;
    wire N__16439;
    wire N__16436;
    wire N__16431;
    wire N__16430;
    wire N__16427;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16416;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16399;
    wire N__16392;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16371;
    wire N__16368;
    wire N__16363;
    wire N__16362;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16335;
    wire N__16332;
    wire N__16331;
    wire N__16330;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16318;
    wire N__16311;
    wire N__16308;
    wire N__16307;
    wire N__16306;
    wire N__16305;
    wire N__16298;
    wire N__16297;
    wire N__16296;
    wire N__16295;
    wire N__16294;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16286;
    wire N__16277;
    wire N__16274;
    wire N__16269;
    wire N__16266;
    wire N__16263;
    wire N__16260;
    wire N__16251;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16235;
    wire N__16230;
    wire N__16227;
    wire N__16224;
    wire N__16223;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16212;
    wire N__16211;
    wire N__16210;
    wire N__16209;
    wire N__16208;
    wire N__16203;
    wire N__16194;
    wire N__16189;
    wire N__16184;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16172;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16110;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16095;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16085;
    wire N__16080;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16032;
    wire N__16029;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16017;
    wire N__16014;
    wire N__16011;
    wire N__16010;
    wire N__16009;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15983;
    wire N__15982;
    wire N__15981;
    wire N__15978;
    wire N__15975;
    wire N__15968;
    wire N__15963;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15945;
    wire N__15944;
    wire N__15943;
    wire N__15940;
    wire N__15935;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15921;
    wire N__15918;
    wire N__15915;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15907;
    wire N__15902;
    wire N__15899;
    wire N__15894;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15879;
    wire N__15876;
    wire N__15873;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15843;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15822;
    wire N__15819;
    wire N__15816;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15808;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15792;
    wire N__15791;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15762;
    wire N__15759;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15747;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15736;
    wire N__15735;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15719;
    wire N__15714;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15702;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15676;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15664;
    wire N__15657;
    wire N__15654;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15623;
    wire N__15620;
    wire N__15617;
    wire N__15612;
    wire N__15611;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15599;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15552;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15544;
    wire N__15541;
    wire N__15540;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15530;
    wire N__15525;
    wire N__15516;
    wire N__15513;
    wire N__15512;
    wire N__15509;
    wire N__15508;
    wire N__15505;
    wire N__15502;
    wire N__15499;
    wire N__15494;
    wire N__15493;
    wire N__15492;
    wire N__15489;
    wire N__15486;
    wire N__15481;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15458;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15441;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15426;
    wire N__15417;
    wire N__15414;
    wire N__15413;
    wire N__15412;
    wire N__15411;
    wire N__15406;
    wire N__15401;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15360;
    wire N__15359;
    wire N__15354;
    wire N__15351;
    wire N__15348;
    wire N__15345;
    wire N__15342;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15330;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15314;
    wire N__15313;
    wire N__15310;
    wire N__15305;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15290;
    wire N__15289;
    wire N__15286;
    wire N__15281;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15266;
    wire N__15265;
    wire N__15262;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15249;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15233;
    wire N__15230;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15213;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15177;
    wire N__15174;
    wire N__15173;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15148;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15123;
    wire N__15122;
    wire N__15121;
    wire N__15120;
    wire N__15111;
    wire N__15110;
    wire N__15109;
    wire N__15108;
    wire N__15107;
    wire N__15104;
    wire N__15095;
    wire N__15090;
    wire N__15087;
    wire N__15084;
    wire N__15081;
    wire N__15078;
    wire N__15075;
    wire N__15072;
    wire N__15069;
    wire N__15068;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15051;
    wire N__15050;
    wire N__15049;
    wire N__15046;
    wire N__15041;
    wire N__15036;
    wire N__15035;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15018;
    wire N__15015;
    wire N__15014;
    wire N__15013;
    wire N__15012;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14996;
    wire N__14995;
    wire N__14994;
    wire N__14993;
    wire N__14992;
    wire N__14991;
    wire N__14988;
    wire N__14985;
    wire N__14982;
    wire N__14975;
    wire N__14972;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14954;
    wire N__14953;
    wire N__14952;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14946;
    wire N__14943;
    wire N__14938;
    wire N__14931;
    wire N__14922;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14905;
    wire N__14898;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14829;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14807;
    wire N__14806;
    wire N__14803;
    wire N__14798;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14775;
    wire N__14774;
    wire N__14773;
    wire N__14770;
    wire N__14765;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14753;
    wire N__14750;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14733;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14714;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14694;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14682;
    wire N__14679;
    wire N__14674;
    wire N__14667;
    wire N__14664;
    wire N__14661;
    wire N__14658;
    wire N__14655;
    wire N__14652;
    wire N__14649;
    wire N__14646;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14598;
    wire N__14595;
    wire N__14594;
    wire N__14591;
    wire N__14590;
    wire N__14587;
    wire N__14586;
    wire N__14583;
    wire N__14576;
    wire N__14571;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14529;
    wire N__14526;
    wire N__14521;
    wire N__14518;
    wire N__14511;
    wire N__14508;
    wire N__14505;
    wire N__14502;
    wire N__14499;
    wire N__14496;
    wire N__14493;
    wire N__14490;
    wire N__14487;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14475;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14465;
    wire N__14464;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire N__14436;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14421;
    wire N__14418;
    wire N__14415;
    wire N__14414;
    wire N__14411;
    wire N__14410;
    wire N__14409;
    wire N__14406;
    wire N__14403;
    wire N__14398;
    wire N__14391;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14367;
    wire N__14366;
    wire N__14365;
    wire N__14364;
    wire N__14361;
    wire N__14358;
    wire N__14355;
    wire N__14352;
    wire N__14349;
    wire N__14340;
    wire N__14337;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14321;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14301;
    wire N__14298;
    wire N__14297;
    wire N__14294;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14277;
    wire N__14274;
    wire N__14273;
    wire N__14272;
    wire N__14271;
    wire N__14268;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14247;
    wire N__14246;
    wire N__14243;
    wire N__14242;
    wire N__14239;
    wire N__14234;
    wire N__14229;
    wire N__14226;
    wire N__14225;
    wire N__14222;
    wire N__14221;
    wire N__14220;
    wire N__14219;
    wire N__14218;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14207;
    wire N__14206;
    wire N__14205;
    wire N__14200;
    wire N__14195;
    wire N__14190;
    wire N__14187;
    wire N__14182;
    wire N__14179;
    wire N__14174;
    wire N__14171;
    wire N__14168;
    wire N__14157;
    wire N__14154;
    wire N__14151;
    wire N__14148;
    wire N__14145;
    wire N__14142;
    wire N__14139;
    wire N__14136;
    wire N__14133;
    wire N__14132;
    wire N__14129;
    wire N__14128;
    wire N__14127;
    wire N__14126;
    wire N__14125;
    wire N__14124;
    wire N__14123;
    wire N__14120;
    wire N__14119;
    wire N__14116;
    wire N__14115;
    wire N__14114;
    wire N__14113;
    wire N__14112;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14104;
    wire N__14101;
    wire N__14100;
    wire N__14099;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14078;
    wire N__14071;
    wire N__14064;
    wire N__14061;
    wire N__14056;
    wire N__14049;
    wire N__14044;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14017;
    wire N__14016;
    wire N__14013;
    wire N__14012;
    wire N__14011;
    wire N__14008;
    wire N__14007;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13992;
    wire N__13989;
    wire N__13982;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13964;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13929;
    wire N__13928;
    wire N__13927;
    wire N__13922;
    wire N__13919;
    wire N__13918;
    wire N__13915;
    wire N__13914;
    wire N__13913;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13895;
    wire N__13890;
    wire N__13881;
    wire N__13880;
    wire N__13879;
    wire N__13878;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13863;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13833;
    wire N__13830;
    wire N__13827;
    wire N__13824;
    wire N__13821;
    wire N__13818;
    wire N__13815;
    wire N__13812;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13802;
    wire N__13799;
    wire N__13798;
    wire N__13797;
    wire N__13796;
    wire N__13793;
    wire N__13790;
    wire N__13789;
    wire N__13788;
    wire N__13787;
    wire N__13784;
    wire N__13779;
    wire N__13774;
    wire N__13767;
    wire N__13766;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13744;
    wire N__13737;
    wire N__13736;
    wire N__13733;
    wire N__13732;
    wire N__13729;
    wire N__13728;
    wire N__13727;
    wire N__13724;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13707;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13664;
    wire N__13663;
    wire N__13660;
    wire N__13659;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13646;
    wire N__13645;
    wire N__13644;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13630;
    wire N__13627;
    wire N__13624;
    wire N__13619;
    wire N__13616;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13592;
    wire N__13591;
    wire N__13588;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13569;
    wire N__13566;
    wire N__13563;
    wire N__13560;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13548;
    wire N__13545;
    wire N__13542;
    wire N__13539;
    wire N__13536;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13524;
    wire N__13521;
    wire N__13518;
    wire N__13515;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13494;
    wire N__13491;
    wire N__13488;
    wire N__13485;
    wire N__13482;
    wire N__13481;
    wire N__13478;
    wire N__13477;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13461;
    wire N__13458;
    wire N__13455;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13434;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13398;
    wire N__13395;
    wire N__13392;
    wire N__13389;
    wire N__13388;
    wire N__13387;
    wire N__13384;
    wire N__13381;
    wire N__13378;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13353;
    wire N__13350;
    wire N__13347;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13307;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13269;
    wire N__13266;
    wire N__13263;
    wire N__13260;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13252;
    wire N__13249;
    wire N__13244;
    wire N__13239;
    wire N__13236;
    wire N__13233;
    wire N__13230;
    wire N__13227;
    wire N__13224;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13209;
    wire N__13206;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13175;
    wire N__13174;
    wire N__13171;
    wire N__13166;
    wire N__13161;
    wire N__13160;
    wire N__13159;
    wire N__13156;
    wire N__13151;
    wire N__13146;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13136;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13126;
    wire N__13119;
    wire N__13118;
    wire N__13117;
    wire N__13116;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13083;
    wire N__13080;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13070;
    wire N__13069;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13057;
    wire N__13050;
    wire N__13049;
    wire N__13048;
    wire N__13047;
    wire N__13042;
    wire N__13037;
    wire N__13032;
    wire N__13031;
    wire N__13030;
    wire N__13027;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13009;
    wire N__13002;
    wire N__13001;
    wire N__12998;
    wire N__12995;
    wire N__12990;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12978;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12966;
    wire N__12965;
    wire N__12964;
    wire N__12963;
    wire N__12962;
    wire N__12961;
    wire N__12960;
    wire N__12959;
    wire N__12958;
    wire N__12953;
    wire N__12950;
    wire N__12947;
    wire N__12938;
    wire N__12935;
    wire N__12930;
    wire N__12921;
    wire N__12920;
    wire N__12917;
    wire N__12916;
    wire N__12913;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12901;
    wire N__12894;
    wire N__12893;
    wire N__12892;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12884;
    wire N__12883;
    wire N__12882;
    wire N__12881;
    wire N__12878;
    wire N__12877;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12858;
    wire N__12853;
    wire N__12850;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12816;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12793;
    wire N__12788;
    wire N__12783;
    wire N__12782;
    wire N__12781;
    wire N__12778;
    wire N__12775;
    wire N__12772;
    wire N__12765;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12750;
    wire N__12747;
    wire N__12746;
    wire N__12745;
    wire N__12742;
    wire N__12737;
    wire N__12732;
    wire N__12731;
    wire N__12730;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12722;
    wire N__12717;
    wire N__12710;
    wire N__12705;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12682;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12651;
    wire N__12648;
    wire N__12645;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12623;
    wire N__12622;
    wire N__12619;
    wire N__12614;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12582;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12546;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12522;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12450;
    wire N__12447;
    wire N__12444;
    wire N__12441;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12273;
    wire N__12270;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12258;
    wire N__12255;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12231;
    wire N__12228;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire \c0.n6111_cascade_ ;
    wire \c0.n5758_cascade_ ;
    wire \c0.n5761 ;
    wire \c0.data_in_frame_18_1 ;
    wire \c0.data_in_frame_19_1 ;
    wire \c0.n6303_cascade_ ;
    wire \c0.n6057_cascade_ ;
    wire \c0.n6306 ;
    wire \c0.n6060_cascade_ ;
    wire \c0.n6087 ;
    wire \c0.n5770 ;
    wire \c0.n5788_cascade_ ;
    wire \c0.n6027_cascade_ ;
    wire \c0.n5794_cascade_ ;
    wire \c0.n6015 ;
    wire \c0.n6072_cascade_ ;
    wire \c0.n6018 ;
    wire \c0.tx2.r_Tx_Data_1 ;
    wire \c0.tx2.r_Tx_Data_0 ;
    wire \c0.tx2.n6048_cascade_ ;
    wire \c0.tx2.o_Tx_Serial_N_1798_cascade_ ;
    wire bfn_1_29_0_;
    wire \c0.tx2.n4779 ;
    wire \c0.tx2.n4780 ;
    wire \c0.tx2.n318 ;
    wire \c0.tx2.n4781 ;
    wire \c0.tx2.n317 ;
    wire \c0.tx2.n4782 ;
    wire \c0.tx2.n4783 ;
    wire \c0.tx2.n4784 ;
    wire \c0.tx2.n4785 ;
    wire \c0.tx2.n4786 ;
    wire bfn_1_30_0_;
    wire n313_adj_1997;
    wire \c0.n6135_cascade_ ;
    wire \c0.n5746_cascade_ ;
    wire \c0.n6153_cascade_ ;
    wire \c0.n5740_cascade_ ;
    wire \c0.n6129 ;
    wire \c0.n6063 ;
    wire \c0.n5776 ;
    wire \c0.n6099 ;
    wire \c0.tx2.n6006 ;
    wire \c0.n5375_cascade_ ;
    wire \c0.n5755 ;
    wire \c0.n6075_cascade_ ;
    wire \c0.n5773 ;
    wire \c0.n5454_cascade_ ;
    wire \c0.n27_cascade_ ;
    wire \c0.n47 ;
    wire \c0.n52_cascade_ ;
    wire \c0.n31 ;
    wire \c0.n32 ;
    wire \c0.n24_adj_1879_cascade_ ;
    wire \c0.n6102 ;
    wire \c0.tx2.r_Tx_Data_2 ;
    wire \c0.tx2.n6045 ;
    wire \c0.data_in_frame_18_2 ;
    wire \c0.n6297_cascade_ ;
    wire \c0.n6300 ;
    wire \c0.data_in_frame_18_3 ;
    wire \c0.n6279_cascade_ ;
    wire \c0.n6282_cascade_ ;
    wire \c0.n6132 ;
    wire \c0.tx2.r_Tx_Data_3 ;
    wire \c0.n6069 ;
    wire \c0.n6249_cascade_ ;
    wire \c0.n28 ;
    wire \c0.n3703_cascade_ ;
    wire \c0.n6117 ;
    wire \c0.n5536_cascade_ ;
    wire \c0.n5570_cascade_ ;
    wire \c0.n27_adj_1910 ;
    wire \c0.n3689_cascade_ ;
    wire \c0.tx2.n12 ;
    wire \c0.n3689 ;
    wire \c0.n3703 ;
    wire \c0.tx2.r_Bit_Index_2 ;
    wire \c0.tx2.n1136 ;
    wire n4_adj_1973_cascade_;
    wire tx2_active;
    wire \c0.r_SM_Main_2_N_1770_0 ;
    wire tx2_o;
    wire tx2_enable;
    wire \c0.tx2.r_Clock_Count_4 ;
    wire r_SM_Main_1_adj_1993;
    wire \c0.tx2.r_SM_Main_2_N_1767_1_cascade_ ;
    wire \c0.tx2.n315 ;
    wire \c0.tx2.n5824 ;
    wire \c0.tx2.n5816 ;
    wire \c0.tx2.n314 ;
    wire \c0.tx2.n319 ;
    wire \c0.tx2.r_Clock_Count_2 ;
    wire \c0.tx2.r_Clock_Count_0 ;
    wire \c0.tx2.r_Clock_Count_1 ;
    wire \c0.tx2.n316 ;
    wire \c0.tx2.r_Clock_Count_5 ;
    wire \c0.tx2.r_Clock_Count_3 ;
    wire \c0.tx2.n14_adj_1867 ;
    wire \c0.rx.r_Rx_Data_R ;
    wire \c0.tx2.r_Clock_Count_7 ;
    wire r_Clock_Count_8_adj_1994;
    wire \c0.tx2.r_Clock_Count_6 ;
    wire \c0.tx2.n31 ;
    wire \c0.tx2.n9 ;
    wire \c0.tx2.n5631_cascade_ ;
    wire \c0.tx2.n78 ;
    wire n4544;
    wire \c0.n6159_cascade_ ;
    wire \c0.n5737 ;
    wire \c0.n5743 ;
    wire \c0.n6141 ;
    wire \c0.n6123_cascade_ ;
    wire \c0.n5752 ;
    wire data_in_14_7;
    wire \c0.n24_adj_1877 ;
    wire \c0.data_in_frame_19_2 ;
    wire \c0.n5381 ;
    wire \c0.n5381_cascade_ ;
    wire data_in_13_7;
    wire \c0.n2009 ;
    wire data_in_16_6;
    wire \c0.n1942_cascade_ ;
    wire \c0.n18_adj_1938 ;
    wire \c0.n5578_cascade_ ;
    wire \c0.n30 ;
    wire \c0.n5488_cascade_ ;
    wire \c0.n36_cascade_ ;
    wire \c0.n45 ;
    wire \c0.n12 ;
    wire \c0.n5488 ;
    wire \c0.n5489 ;
    wire \c0.n1886 ;
    wire \c0.n1942 ;
    wire \c0.n12_adj_1951 ;
    wire data_in_14_2;
    wire \c0.n5536 ;
    wire \c0.n5586 ;
    wire \c0.data_in_frame_19_3 ;
    wire \c0.n22_adj_1876 ;
    wire \c0.data_in_field_49 ;
    wire \c0.n5991_cascade_ ;
    wire \c0.n6105 ;
    wire \c0.data_in_frame_18_5 ;
    wire \c0.n6225_cascade_ ;
    wire \c0.n6228_cascade_ ;
    wire \c0.tx2.r_Tx_Data_5 ;
    wire \c0.n6267_cascade_ ;
    wire \c0.n6270_cascade_ ;
    wire \c0.tx2.r_Tx_Data_4 ;
    wire \c0.n6081 ;
    wire \c0.n6084 ;
    wire \c0.n5695 ;
    wire \c0.n6234_cascade_ ;
    wire \c0.n1081 ;
    wire \c0.tx2.n1624 ;
    wire \c0.tx2.r_Tx_Data_7 ;
    wire \c0.tx2.r_Tx_Data_6 ;
    wire \c0.tx2.r_Bit_Index_1 ;
    wire \c0.tx2.n6003 ;
    wire \c0.FRAME_MATCHER_wait_for_transmission_N_909 ;
    wire bfn_3_26_0_;
    wire \c0.n4735 ;
    wire \c0.n4736 ;
    wire \c0.n4737 ;
    wire \c0.n4738 ;
    wire \c0.byte_transmit_counter2_4 ;
    wire \c0.n195 ;
    wire \c0.n2325 ;
    wire r_SM_Main_2_adj_1992;
    wire \c0.tx2.n14 ;
    wire \c0.tx2.r_SM_Main_0 ;
    wire n2208;
    wire n2339;
    wire r_Bit_Index_0_adj_1995;
    wire \c0.tx2.r_SM_Main_2_N_1767_1 ;
    wire \c0.tx2.n5847 ;
    wire \c0.rx.n3589 ;
    wire \c0.rx.n3589_cascade_ ;
    wire \c0.rx.n17_cascade_ ;
    wire \c0.rx.n5817 ;
    wire data_in_15_3;
    wire \c0.data_in_field_59 ;
    wire \c0.data_in_field_123 ;
    wire data_in_7_3;
    wire \c0.data_in_field_11 ;
    wire data_in_8_3;
    wire \c0.data_in_field_67 ;
    wire data_in_10_3;
    wire \c0.n5412_cascade_ ;
    wire \c0.n16_adj_1880 ;
    wire \c0.n22_adj_1881_cascade_ ;
    wire \c0.n24_adj_1884 ;
    wire \c0.data_in_field_81 ;
    wire \c0.n5551 ;
    wire \c0.n5551_cascade_ ;
    wire \c0.n1892 ;
    wire \c0.n20 ;
    wire \c0.n19_cascade_ ;
    wire \c0.n5578 ;
    wire \c0.n6177_cascade_ ;
    wire \c0.n5728_cascade_ ;
    wire \c0.n16_adj_1873_cascade_ ;
    wire \c0.n24 ;
    wire \c0.n5725 ;
    wire \c0.n6165 ;
    wire \c0.n6168 ;
    wire \c0.n20_adj_1878 ;
    wire data_in_7_2;
    wire \c0.data_in_field_58 ;
    wire \c0.data_in_frame_19_6 ;
    wire \c0.n6147_cascade_ ;
    wire \c0.n6150 ;
    wire \c0.data_in_frame_19_4 ;
    wire \c0.data_in_field_14 ;
    wire \c0.n6255_cascade_ ;
    wire \c0.n5692 ;
    wire \c0.data_in_field_119 ;
    wire \c0.n6273_cascade_ ;
    wire \c0.data_in_field_111 ;
    wire \c0.n5994 ;
    wire \c0.n5686_cascade_ ;
    wire \c0.n6261_cascade_ ;
    wire \c0.n6264 ;
    wire data_in_18_3;
    wire \c0.data_in_field_104 ;
    wire \c0.n6021_cascade_ ;
    wire \c0.n5797 ;
    wire bfn_4_27_0_;
    wire \c0.rx.n5860 ;
    wire \c0.rx.n4772 ;
    wire \c0.rx.n4773 ;
    wire \c0.rx.n5856 ;
    wire \c0.rx.n4774 ;
    wire \c0.rx.n4775 ;
    wire \c0.rx.n4776 ;
    wire \c0.rx.n4777 ;
    wire \c0.rx.n36 ;
    wire \c0.rx.n4778 ;
    wire \c0.rx.n5361 ;
    wire \c0.rx.n5858 ;
    wire \c0.rx.n5854 ;
    wire \c0.rx.r_Clock_Count_3 ;
    wire \c0.rx.r_Clock_Count_6 ;
    wire \c0.rx.r_Clock_Count_5 ;
    wire \c0.rx.n8_cascade_ ;
    wire \c0.rx.n1724 ;
    wire \c0.rx.n1724_cascade_ ;
    wire \c0.rx.r_Clock_Count_1 ;
    wire \c0.rx.n5855 ;
    wire \c0.rx.r_Clock_Count_0 ;
    wire \c0.rx.n5857 ;
    wire \c0.rx.r_Clock_Count_4 ;
    wire tx_enable;
    wire data_in_16_3;
    wire rx_data_3;
    wire data_in_18_1;
    wire \c0.n6009_cascade_ ;
    wire \c0.n6012 ;
    wire \c0.data_in_field_15 ;
    wire \c0.data_in_field_8 ;
    wire \c0.n2039 ;
    wire \c0.n2039_cascade_ ;
    wire \c0.data_in_field_23 ;
    wire \c0.data_in_field_138 ;
    wire \c0.data_in_field_130 ;
    wire \c0.n6213 ;
    wire \c0.data_in_field_73 ;
    wire \c0.n14_adj_1957_cascade_ ;
    wire \c0.data_in_field_53 ;
    wire \c0.n22_adj_1903_cascade_ ;
    wire \c0.n18_adj_1904 ;
    wire \c0.n20_adj_1905 ;
    wire \c0.n5589_cascade_ ;
    wire \c0.n29 ;
    wire \c0.n5458 ;
    wire \c0.n1994 ;
    wire \c0.n5557 ;
    wire \c0.n17_cascade_ ;
    wire \c0.n5574 ;
    wire \c0.n5572 ;
    wire data_in_8_7;
    wire data_in_17_1;
    wire \c0.n1973 ;
    wire data_in_19_3;
    wire \c0.n18_adj_1959_cascade_ ;
    wire \c0.n16 ;
    wire \c0.n20_adj_1870_cascade_ ;
    wire \c0.n5577 ;
    wire \c0.n2101_cascade_ ;
    wire \c0.n6_adj_1917_cascade_ ;
    wire \c0.data_in_field_68 ;
    wire \c0.n5512 ;
    wire \c0.n5512_cascade_ ;
    wire \c0.n22 ;
    wire \c0.n2155 ;
    wire \c0.n2155_cascade_ ;
    wire \c0.n43 ;
    wire \c0.n2026 ;
    wire data_in_16_1;
    wire \c0.n2080 ;
    wire \c0.n2012 ;
    wire data_in_19_6;
    wire \c0.data_in_frame_19_0 ;
    wire \c0.data_in_field_17 ;
    wire \c0.n6093_cascade_ ;
    wire \c0.n5767 ;
    wire data_in_16_2;
    wire data_in_18_6;
    wire \c0.data_in_frame_18_6 ;
    wire \c0.data_in_frame_18_7 ;
    wire data_in_7_1;
    wire n1764_cascade_;
    wire rx_data_5;
    wire rx_data_6;
    wire \c0.rx.n5822 ;
    wire \c0.rx.r_Clock_Count_2 ;
    wire n4_adj_1980;
    wire n4_adj_1980_cascade_;
    wire rx_data_4;
    wire n2198_cascade_;
    wire \c0.rx.n359 ;
    wire \c0.rx.n5859 ;
    wire \c0.rx.r_Clock_Count_7 ;
    wire \c0.rx.n5823 ;
    wire \c0.rx.n6294_cascade_ ;
    wire r_SM_Main_2_adj_1989;
    wire \c0.rx.n75_cascade_ ;
    wire \c0.rx.n5815 ;
    wire data_in_1_3;
    wire data_in_6_3;
    wire data_in_12_3;
    wire data_in_2_7;
    wire \c0.data_in_field_131 ;
    wire data_in_1_1;
    wire \c0.data_in_field_7 ;
    wire data_in_0_1;
    wire \c0.n2104 ;
    wire \c0.n1835 ;
    wire \c0.n2104_cascade_ ;
    wire data_in_8_1;
    wire \c0.n20_adj_1958 ;
    wire \c0.n31_adj_1896_cascade_ ;
    wire \c0.n41 ;
    wire \c0.data_in_field_6 ;
    wire \c0.n10_adj_1915 ;
    wire \c0.n1913 ;
    wire \c0.data_in_field_64 ;
    wire data_in_8_2;
    wire data_in_5_3;
    wire \c0.n6183 ;
    wire \c0.n2062_cascade_ ;
    wire \c0.n44 ;
    wire \c0.data_in_field_134 ;
    wire \c0.n5503 ;
    wire \c0.n2095 ;
    wire \c0.n16_adj_1871 ;
    wire data_in_11_3;
    wire \c0.n2021 ;
    wire \c0.data_in_field_10 ;
    wire \c0.n2021_cascade_ ;
    wire \c0.data_in_field_41 ;
    wire \c0.n2074_cascade_ ;
    wire \c0.n2000 ;
    wire \c0.data_in_field_26 ;
    wire \c0.data_in_field_135 ;
    wire \c0.n1908 ;
    wire \c0.data_in_field_99 ;
    wire \c0.data_in_field_65 ;
    wire \c0.data_in_field_129 ;
    wire \c0.n5569 ;
    wire \c0.n5569_cascade_ ;
    wire \c0.data_in_field_114 ;
    wire \c0.n20_adj_1882 ;
    wire \c0.n5388 ;
    wire \c0.n5418 ;
    wire \c0.n5491 ;
    wire \c0.n44_adj_1894 ;
    wire \c0.data_in_field_112 ;
    wire \c0.data_in_field_30 ;
    wire \c0.data_in_field_125 ;
    wire \c0.n1889 ;
    wire \c0.data_in_field_76 ;
    wire \c0.data_in_frame_18_4 ;
    wire \c0.n6243_cascade_ ;
    wire \c0.n5698_cascade_ ;
    wire \c0.n6231 ;
    wire \c0.n6237 ;
    wire \c0.data_in_field_102 ;
    wire \c0.n5701 ;
    wire data_in_10_6;
    wire \c0.data_in_field_86 ;
    wire data_in_10_1;
    wire data_in_9_1;
    wire data_in_12_6;
    wire n1764;
    wire rx_data_7;
    wire data_in_15_6;
    wire r_SM_Main_0_adj_1991;
    wire r_SM_Main_2_N_1824_2;
    wire \c0.rx.n6291 ;
    wire \c0.rx.n5633 ;
    wire n3636;
    wire \c0.rx.n3850 ;
    wire r_SM_Main_1_adj_1990;
    wire \c0.rx.n3850_cascade_ ;
    wire \c0.rx.n2259 ;
    wire \c0.rx.n2367 ;
    wire data_in_2_5;
    wire \c0.n26 ;
    wire \c0.n27_adj_1928 ;
    wire \c0.n28_adj_1926_cascade_ ;
    wire \c0.n25_adj_1929 ;
    wire data_in_2_1;
    wire data_in_1_0;
    wire data_in_0_6;
    wire data_in_3_7;
    wire data_in_1_6;
    wire data_in_1_7;
    wire data_in_0_7;
    wire \c0.n30_adj_1941 ;
    wire \c0.n4795 ;
    wire \c0.n26_adj_1940 ;
    wire \c0.n1729_cascade_ ;
    wire \c0.data_in_field_35 ;
    wire \c0.data_in_field_9 ;
    wire \c0.data_in_field_54 ;
    wire \c0.n5369_cascade_ ;
    wire data_in_0_3;
    wire data_in_9_3;
    wire \c0.data_in_field_3 ;
    wire \c0.n2125 ;
    wire \c0.data_in_field_27 ;
    wire \c0.n5469 ;
    wire \c0.data_in_field_83 ;
    wire \c0.n5454 ;
    wire \c0.n5469_cascade_ ;
    wire \c0.n6_adj_1923 ;
    wire \c0.n5548_cascade_ ;
    wire data_in_0_4;
    wire data_in_7_5;
    wire \c0.data_in_field_33 ;
    wire \c0.data_in_field_140 ;
    wire data_in_12_7;
    wire \c0.data_in_field_126 ;
    wire \c0.data_in_field_118 ;
    wire \c0.data_in_field_51 ;
    wire data_in_16_5;
    wire \c0.data_in_field_52 ;
    wire \c0.data_in_field_103 ;
    wire \c0.n2152 ;
    wire \c0.data_in_field_43 ;
    wire \c0.n2152_cascade_ ;
    wire \c0.n5397 ;
    wire data_in_11_6;
    wire \c0.data_in_field_75 ;
    wire data_in_17_6;
    wire \c0.data_in_field_142 ;
    wire \c0.tx2_transmit_N_1031_cascade_ ;
    wire \c0.data_in_field_29 ;
    wire \c0.n2030 ;
    wire \c0.n2030_cascade_ ;
    wire data_in_15_2;
    wire \c0.data_in_field_22 ;
    wire \c0.n5436 ;
    wire \c0.n5436_cascade_ ;
    wire \c0.n5509 ;
    wire \c0.data_in_field_78 ;
    wire \c0.n5509_cascade_ ;
    wire \c0.data_in_field_92 ;
    wire \c0.data_in_field_36 ;
    wire \c0.data_in_field_82 ;
    wire \c0.n1948 ;
    wire data_in_15_1;
    wire data_in_14_1;
    wire \c0.data_in_field_127 ;
    wire n4;
    wire data_in_13_1;
    wire \c0.data_in_field_105 ;
    wire \c0.n18_adj_1887 ;
    wire \c0.n20_adj_1888 ;
    wire data_in_12_1;
    wire \c0.data_in_field_97 ;
    wire \c0.data_in_frame_19_5 ;
    wire data_in_14_6;
    wire data_in_19_7;
    wire \c0.data_in_frame_19_7 ;
    wire data_in_19_5;
    wire data_in_14_0;
    wire data_in_13_0;
    wire data_in_18_4;
    wire \c0.tx.n40_cascade_ ;
    wire n1760;
    wire \c0.tx.n2247 ;
    wire \c0.tx.n2356 ;
    wire \c0.rx.r_Bit_Index_2 ;
    wire \c0.rx.r_Bit_Index_1 ;
    wire \c0.rx.n1706 ;
    wire n1757_cascade_;
    wire rx_data_0;
    wire r_Bit_Index_0;
    wire r_Rx_Data;
    wire n1757;
    wire data_in_3_6;
    wire data_in_0_5;
    wire \c0.n22_adj_1924 ;
    wire \c0.data_in_field_141 ;
    wire \c0.n5527 ;
    wire \c0.n5394_cascade_ ;
    wire \c0.n1926 ;
    wire \c0.n19_adj_1889 ;
    wire \c0.n22_adj_1886 ;
    wire \c0.n5590 ;
    wire \c0.n40_cascade_ ;
    wire \c0.n45_adj_1892 ;
    wire \c0.data_in_field_132 ;
    wire \c0.n1969 ;
    wire \c0.n5403 ;
    wire data_in_19_4;
    wire \c0.data_in_field_115 ;
    wire \c0.n1855_cascade_ ;
    wire \c0.n1917 ;
    wire \c0.data_in_field_34 ;
    wire \c0.n2092 ;
    wire data_in_17_3;
    wire data_in_2_3;
    wire data_in_6_7;
    wire data_in_6_5;
    wire \c0.n25_adj_1948 ;
    wire \c0.data_in_field_94 ;
    wire \c0.data_in_field_66 ;
    wire \c0.data_in_field_79 ;
    wire \c0.n5545 ;
    wire \c0.n46 ;
    wire \c0.data_in_field_95 ;
    wire \c0.data_in_field_96 ;
    wire data_in_15_5;
    wire \c0.n6414 ;
    wire \c0.n5563 ;
    wire data_in_11_1;
    wire \c0.data_in_field_45 ;
    wire \c0.n2065 ;
    wire \c0.n18 ;
    wire \c0.n2149_cascade_ ;
    wire \c0.n21 ;
    wire data_in_3_2;
    wire \c0.n1955 ;
    wire data_in_4_2;
    wire data_in_18_5;
    wire data_in_17_5;
    wire bfn_9_23_0_;
    wire \c0.n4754 ;
    wire \c0.n4755 ;
    wire \c0.n4756 ;
    wire \c0.n4757 ;
    wire \c0.n4758 ;
    wire \c0.n4759 ;
    wire \c0.n4760 ;
    wire \c0.n4761 ;
    wire bfn_9_24_0_;
    wire \c0.n4762 ;
    wire \c0.n4763 ;
    wire \c0.delay_counter_1 ;
    wire \c0.delay_counter_5 ;
    wire \c0.data_in_field_116 ;
    wire \c0.data_in_field_124 ;
    wire \c0.n6171_cascade_ ;
    wire \c0.n5731 ;
    wire \c0.data_in_field_4 ;
    wire \c0.data_in_field_12 ;
    wire \c0.n5722 ;
    wire \c0.tx.n3631_cascade_ ;
    wire \c0.data_in_field_20 ;
    wire \c0.n6189 ;
    wire \c0.tx.n5812_cascade_ ;
    wire \c0.tx.n14_cascade_ ;
    wire r_Tx_Data_7;
    wire r_Tx_Data_6;
    wire bfn_9_27_0_;
    wire \c0.tx.n4764 ;
    wire \c0.tx.n4765 ;
    wire \c0.tx.n4766 ;
    wire \c0.tx.n4767 ;
    wire \c0.tx.n4768 ;
    wire \c0.tx.n4769 ;
    wire \c0.tx.n4770 ;
    wire \c0.tx.n4771 ;
    wire bfn_9_28_0_;
    wire \c0.tx.n5885 ;
    wire \c0.tx.n15 ;
    wire \c0.tx.n5884 ;
    wire data_in_4_3;
    wire data_in_3_3;
    wire data_in_2_2;
    wire data_in_1_2;
    wire \c0.data_in_field_80 ;
    wire \c0.n42_cascade_ ;
    wire \c0.n48 ;
    wire data_in_19_0;
    wire data_in_15_7;
    wire data_in_16_7;
    wire \c0.n25 ;
    wire \c0.n23 ;
    wire \c0.n22_adj_1890 ;
    wire \c0.data_in_field_61 ;
    wire data_in_3_1;
    wire data_in_0_0;
    wire \c0.data_in_field_0 ;
    wire \c0.data_in_field_117 ;
    wire \c0.n1855 ;
    wire \c0.n13 ;
    wire \c0.n12_adj_1898_cascade_ ;
    wire \c0.n47_adj_1897 ;
    wire \c0.n48_adj_1895 ;
    wire \c0.n5567_cascade_ ;
    wire \c0.n49 ;
    wire \c0.n6219 ;
    wire \c0.data_in_field_5 ;
    wire \c0.n1979 ;
    wire \c0.n1958 ;
    wire \c0.n2056 ;
    wire \c0.n5506 ;
    wire \c0.n5575 ;
    wire \c0.n5506_cascade_ ;
    wire \c0.n5539 ;
    wire \c0.n1779 ;
    wire \c0.data_in_field_60 ;
    wire \c0.n5500 ;
    wire \c0.data_in_field_19 ;
    wire \c0.data_in_field_139 ;
    wire data_in_5_5;
    wire data_in_6_1;
    wire data_in_5_1;
    wire data_in_4_1;
    wire data_in_18_7;
    wire data_in_17_7;
    wire \c0.n6_adj_1918 ;
    wire data_in_1_4;
    wire \c0.data_in_field_18 ;
    wire \c0.n5372 ;
    wire \c0.n2043_cascade_ ;
    wire \c0.data_in_field_107 ;
    wire data_in_13_6;
    wire \c0.n5443 ;
    wire \c0.data_in_field_89 ;
    wire \c0.data_in_field_90 ;
    wire data_in_7_7;
    wire \c0.data_in_field_37 ;
    wire \c0.data_in_frame_18_0 ;
    wire \c0.n2077 ;
    wire \c0.n5707 ;
    wire \c0.n5710 ;
    wire \c0.n6198 ;
    wire \c0.delay_counter_9 ;
    wire \c0.delay_counter_2 ;
    wire \c0.delay_counter_0 ;
    wire \c0.delay_counter_7 ;
    wire data_in_5_0;
    wire data_in_4_0;
    wire data_in_8_4;
    wire data_in_7_4;
    wire data_in_6_4;
    wire data_in_5_6;
    wire n5646_cascade_;
    wire n5645;
    wire LED_c;
    wire \c0.data_in_field_110 ;
    wire \c0.n5533 ;
    wire data_out_18_6;
    wire \c0.n17_adj_1913_cascade_ ;
    wire \c0.tx.n5883 ;
    wire \c0.n1253_cascade_ ;
    wire \c0.n5830 ;
    wire \c0.n22_adj_1914_cascade_ ;
    wire tx_data_6_N_keep;
    wire \c0.n5827 ;
    wire \c0.n1253 ;
    wire tx_data_7_N_keep;
    wire data_out_18_0;
    wire data_out_19_0;
    wire \c0.n1198 ;
    wire \c0.n5810_cascade_ ;
    wire \c0.tx_data_0_N ;
    wire \c0.tx.n14_adj_1869_cascade_ ;
    wire \c0.tx.r_SM_Main_2_N_1767_1_cascade_ ;
    wire \c0.tx.n5821 ;
    wire \c0.tx.r_Clock_Count_5 ;
    wire n315;
    wire r_Clock_Count_6;
    wire n317;
    wire r_Clock_Count_4;
    wire \c0.tx.n10_adj_1868 ;
    wire \c0.tx.r_Clock_Count_7 ;
    wire \c0.tx.n5627 ;
    wire n11_adj_1979_cascade_;
    wire \c0.tx.n5629 ;
    wire \c0.tx.n3120 ;
    wire \c0.tx.r_Clock_Count_2 ;
    wire \c0.tx.n3120_cascade_ ;
    wire n313;
    wire n782_cascade_;
    wire r_Clock_Count_8;
    wire data_in_9_2;
    wire \c0.n5384 ;
    wire \c0.n5476 ;
    wire \c0.n5427 ;
    wire \c0.n5521 ;
    wire \c0.n24_adj_1885 ;
    wire \c0.n1866 ;
    wire \c0.data_in_field_113 ;
    wire \c0.data_in_field_57 ;
    wire \c0.n10_cascade_ ;
    wire \c0.n5466 ;
    wire \c0.n5519 ;
    wire data_in_7_6;
    wire data_in_6_6;
    wire data_in_18_0;
    wire \c0.n5548 ;
    wire \c0.n5497 ;
    wire \c0.n5515 ;
    wire \c0.data_in_field_44 ;
    wire \c0.data_in_field_100 ;
    wire \c0.data_in_field_50 ;
    wire \c0.n2053 ;
    wire \c0.n2101 ;
    wire \c0.n2134 ;
    wire \c0.n31_adj_1900_cascade_ ;
    wire \c0.n35 ;
    wire data_in_0_2;
    wire \c0.n14 ;
    wire \c0.n5582 ;
    wire \c0.n13_adj_1899 ;
    wire \c0.n17_adj_1902 ;
    wire \c0.n25_adj_1907 ;
    wire \c0.n4_adj_1920 ;
    wire \c0.data_in_field_122 ;
    wire \c0.n5593 ;
    wire \c0.data_in_field_62 ;
    wire \c0.n5593_cascade_ ;
    wire \c0.n5430 ;
    wire \c0.n33 ;
    wire \c0.n5430_cascade_ ;
    wire \c0.n28_adj_1955 ;
    wire \c0.n37 ;
    wire data_in_1_5;
    wire \c0.data_in_field_13 ;
    wire \c0.n6_adj_1939 ;
    wire data_in_12_4;
    wire data_in_11_4;
    wire \c0.n2089 ;
    wire \c0.n2074 ;
    wire \c0.n5581 ;
    wire \c0.data_in_field_120 ;
    wire \c0.n2107 ;
    wire rx_data_2;
    wire \c0.n6201 ;
    wire \c0.data_in_field_101 ;
    wire \c0.byte_transmit_counter2_3 ;
    wire \c0.byte_transmit_counter2_2 ;
    wire \c0.n5716_cascade_ ;
    wire \c0.n6195 ;
    wire \c0.data_in_field_85 ;
    wire \c0.data_in_field_93 ;
    wire \c0.data_in_field_77 ;
    wire \c0.n6207_cascade_ ;
    wire \c0.data_in_field_69 ;
    wire \c0.n5713 ;
    wire data_in_19_2;
    wire data_in_9_0;
    wire \c0.data_in_field_42 ;
    wire \c0.data_in_field_72 ;
    wire data_in_12_0;
    wire data_in_18_2;
    wire data_in_17_2;
    wire data_in_6_2;
    wire data_in_5_2;
    wire data_in_4_5;
    wire data_in_11_7;
    wire n5448_cascade_;
    wire n4_adj_1975;
    wire data_out_19_4;
    wire data_out_18_4;
    wire \c0.delay_counter_3 ;
    wire \c0.delay_counter_6 ;
    wire \c0.delay_counter_10 ;
    wire \c0.n18_adj_1919 ;
    wire \c0.delay_counter_8 ;
    wire \c0.delay_counter_4 ;
    wire \c0.n20_adj_1922_cascade_ ;
    wire \c0.n16_adj_1921 ;
    wire n4334_cascade_;
    wire n1991;
    wire data_out_19_7;
    wire \c0.n17_adj_1950 ;
    wire n4_adj_1982;
    wire \c0.n17_adj_1908 ;
    wire data_out_18_7;
    wire \c0.n1508 ;
    wire data_out_19_2;
    wire \c0.n1508_cascade_ ;
    wire \c0.n5840 ;
    wire \c0.n6309_cascade_ ;
    wire data_out_18_2;
    wire \c0.n1249 ;
    wire tx_data_4_N_keep;
    wire \c0.tx.n3644 ;
    wire n11_adj_1979;
    wire n5818_cascade_;
    wire n4155;
    wire n318;
    wire r_Clock_Count_3;
    wire n321;
    wire r_Clock_Count_0;
    wire data_out_18_5;
    wire n782;
    wire n320;
    wire r_Clock_Count_1;
    wire rx_data_1;
    wire data_in_14_3;
    wire data_in_13_3;
    wire \c0.data_in_field_55 ;
    wire \c0.data_in_field_63 ;
    wire data_in_14_4;
    wire \c0.data_in_field_48 ;
    wire \c0.data_in_field_32 ;
    wire \c0.data_in_field_40 ;
    wire \c0.n6033_cascade_ ;
    wire \c0.n5791 ;
    wire \c0.n1814 ;
    wire data_in_19_1;
    wire \c0.n2143 ;
    wire \c0.n1814_cascade_ ;
    wire \c0.data_in_field_109 ;
    wire \c0.n32_adj_1901 ;
    wire data_in_8_5;
    wire data_in_17_4;
    wire data_in_5_4;
    wire \c0.n5560 ;
    wire \c0.data_in_field_106 ;
    wire \c0.data_in_field_2 ;
    wire \c0.n5560_cascade_ ;
    wire \c0.n34 ;
    wire data_in_5_7;
    wire \c0.data_in_field_133 ;
    wire \c0.data_in_field_21 ;
    wire \c0.data_in_field_143 ;
    wire \c0.n5378 ;
    wire data_in_11_5;
    wire data_in_2_0;
    wire data_in_13_2;
    wire \c0.data_in_field_88 ;
    wire \c0.data_in_field_98 ;
    wire \c0.data_in_field_28 ;
    wire \c0.data_in_field_121 ;
    wire \c0.n23_adj_1935 ;
    wire \c0.data_in_field_87 ;
    wire \c0.data_in_field_128 ;
    wire \c0.n2068 ;
    wire \c0.data_in_field_46 ;
    wire \c0.n1965_cascade_ ;
    wire \c0.data_in_field_91 ;
    wire \c0.n24_adj_1930 ;
    wire data_in_3_5;
    wire data_in_3_0;
    wire data_in_2_6;
    wire \c0.n28_adj_1925 ;
    wire \c0.byte_transmit_counter2_0 ;
    wire \c0.data_in_field_24 ;
    wire \c0.n6039 ;
    wire n5_cascade_;
    wire \c0.tx_active_prev ;
    wire \c0.tx.r_SM_Main_2_N_1767_1 ;
    wire \c0.tx.n2177 ;
    wire n4333_cascade_;
    wire \c0.n81_adj_1872_cascade_ ;
    wire tx_active;
    wire \c0.tx_transmit ;
    wire n135;
    wire n4_adj_1986_cascade_;
    wire data_out_19_6;
    wire data_out_19_5;
    wire n5440;
    wire \c0.n9 ;
    wire n8_adj_1987;
    wire n5400;
    wire tx_data_2_N_keep;
    wire n5364;
    wire n5482;
    wire n1768;
    wire n5364_cascade_;
    wire n5871;
    wire \c0.n6312 ;
    wire tx_data_3_N_keep;
    wire \c0.n5853 ;
    wire r_Tx_Data_3;
    wire r_Tx_Data_2;
    wire \c0.tx.r_Bit_Index_0 ;
    wire \c0.tx.r_Tx_Data_0 ;
    wire \c0.tx.n6051_cascade_ ;
    wire r_Tx_Data_1;
    wire \c0.tx.r_Bit_Index_2 ;
    wire \c0.tx.n6054 ;
    wire r_SM_Main_0;
    wire \c0.tx.o_Tx_Serial_N_1798_cascade_ ;
    wire r_SM_Main_1;
    wire \c0.tx.n12_cascade_ ;
    wire r_SM_Main_2;
    wire tx_o;
    wire data_in_10_5;
    wire data_in_9_5;
    wire data_in_6_0;
    wire data_in_10_4;
    wire data_in_9_4;
    wire data_in_16_4;
    wire data_in_15_4;
    wire data_in_13_4;
    wire \c0.data_in_field_108 ;
    wire \c0.byte_transmit_counter2_1 ;
    wire \c0.data_in_field_47 ;
    wire \c0.n5997 ;
    wire \c0.n6000 ;
    wire \c0.data_in_field_84 ;
    wire \c0.data_in_field_70 ;
    wire \c0.data_in_field_56 ;
    wire \c0.n5494 ;
    wire \c0.n5554 ;
    wire \c0.n5524 ;
    wire \c0.n5494_cascade_ ;
    wire \c0.n5391 ;
    wire \c0.n26_adj_1927 ;
    wire data_in_8_0;
    wire data_in_7_0;
    wire \c0.data_in_field_74 ;
    wire \c0.data_in_field_1 ;
    wire \c0.data_in_field_16 ;
    wire \c0.n25_adj_1931 ;
    wire \c0.data_in_field_137 ;
    wire \c0.data_in_field_25 ;
    wire \c0.data_in_field_71 ;
    wire \c0.n5542 ;
    wire data_in_17_0;
    wire data_in_10_2;
    wire data_in_4_6;
    wire \c0.data_in_field_38 ;
    wire \c0.data_in_field_136 ;
    wire \c0.data_in_field_31 ;
    wire \c0.n2113 ;
    wire data_in_11_0;
    wire data_in_10_0;
    wire \c0.FRAME_MATCHER_wait_for_transmission ;
    wire \c0.n1729 ;
    wire data_in_4_7;
    wire \c0.data_in_field_39 ;
    wire data_in_10_7;
    wire data_in_9_7;
    wire data_in_14_5;
    wire data_in_12_2;
    wire data_in_11_2;
    wire data_in_4_4;
    wire data_in_9_6;
    wire data_in_8_6;
    wire data_in_3_4;
    wire data_in_2_4;
    wire \c0.n50_adj_1875 ;
    wire bfn_13_23_0_;
    wire \c0.n4703 ;
    wire \c0.n4704 ;
    wire \c0.n4705 ;
    wire \c0.n4706 ;
    wire \c0.byte_transmit_counter_5 ;
    wire \c0.tx_transmit_N_568_5 ;
    wire \c0.n4707 ;
    wire \c0.byte_transmit_counter_6 ;
    wire \c0.tx_transmit_N_568_6 ;
    wire \c0.n4708 ;
    wire \c0.byte_transmit_counter_7 ;
    wire \c0.n4709 ;
    wire \c0.tx_transmit_N_568_7 ;
    wire \c0.tx_transmit_N_568_3 ;
    wire \c0.n95 ;
    wire \c0.n95_cascade_ ;
    wire \c0.n106 ;
    wire n4_adj_1981;
    wire n7_adj_1988;
    wire \c0.n15 ;
    wire \c0.n81_adj_1872 ;
    wire \c0.tx_transmit_N_568_4 ;
    wire \c0.tx_transmit_N_568_2 ;
    wire \c0.n5833 ;
    wire \c0.n31_adj_1912 ;
    wire \c0.n989 ;
    wire \c0.n9_adj_1906_cascade_ ;
    wire \c0.n15_adj_1909 ;
    wire data_out_10_4;
    wire \c0.n2293 ;
    wire n4_adj_1996;
    wire n1519;
    wire tx_data_5_N_keep;
    wire n5421;
    wire data_out_18_1;
    wire data_out_19_3;
    wire \c0.n5837 ;
    wire r_Tx_Data_5;
    wire \c0.tx.r_Bit_Index_1 ;
    wire r_Tx_Data_4;
    wire \c0.tx.n6285 ;
    wire \c0.tx.n6288 ;
    wire n5415;
    wire \c0.n1251 ;
    wire \c0.n5845 ;
    wire \c0.byte_transmit_counter_4 ;
    wire tx_data_1_N_keep;
    wire data_out_11_7;
    wire data_in_13_5;
    wire data_in_12_5;
    wire data_out_10_5;
    wire \c0.n9_adj_1911 ;
    wire data_out_10_0;
    wire \c0.byte_transmit_counter_0 ;
    wire \c0.byte_transmit_counter_3 ;
    wire \c0.byte_transmit_counter_2 ;
    wire \c0.n9_adj_1891_cascade_ ;
    wire \c0.byte_transmit_counter_1 ;
    wire \c0.n15_adj_1893 ;
    wire data_out_11_5;
    wire data_out_10_6;
    wire n4_adj_1976;
    wire n26;
    wire bfn_14_25_0_;
    wire n25;
    wire n4710;
    wire n24;
    wire n4711;
    wire n23;
    wire n4712;
    wire n22;
    wire n4713;
    wire n21;
    wire n4714;
    wire n20;
    wire n4715;
    wire n19;
    wire n4716;
    wire n4717;
    wire n18;
    wire bfn_14_26_0_;
    wire n17;
    wire n4718;
    wire n16;
    wire n4719;
    wire n15;
    wire n4720;
    wire n14;
    wire n4721;
    wire n13;
    wire n4722;
    wire n12;
    wire n4723;
    wire n11;
    wire n4724;
    wire n4725;
    wire n10;
    wire bfn_14_27_0_;
    wire n9;
    wire n4726;
    wire n8;
    wire n4727;
    wire n7;
    wire n4728;
    wire n6;
    wire n4729;
    wire blink_counter_21;
    wire n4730;
    wire blink_counter_22;
    wire n4731;
    wire blink_counter_23;
    wire n4732;
    wire n4733;
    wire blink_counter_24;
    wire bfn_14_28_0_;
    wire n4734;
    wire blink_counter_25;
    wire data_out_10_2;
    wire data_out_11_6;
    wire rx_data_ready;
    wire data_in_16_0;
    wire data_in_15_0;
    wire \c0.n5409 ;
    wire data_out_11_1;
    wire \c0.n5409_cascade_ ;
    wire data_out_11_4;
    wire n4_adj_1978;
    wire n4_adj_1983;
    wire data_out_11_2;
    wire n21_adj_1977;
    wire n4333;
    wire data_out_10_1;
    wire data_out_10_3;
    wire n5424;
    wire data_out_11_0;
    wire data_out_10_7;
    wire n5479;
    wire data_out_11_3;
    wire n8_adj_1984;
    wire n7_adj_1985_cascade_;
    wire data_out_19_1;
    wire data_0;
    wire bfn_15_26_0_;
    wire data_1;
    wire \c0.n4739 ;
    wire data_2;
    wire \c0.n4740 ;
    wire data_3;
    wire \c0.n4741 ;
    wire data_4;
    wire \c0.n4742 ;
    wire data_5;
    wire \c0.n4743 ;
    wire data_6;
    wire \c0.n4744 ;
    wire data_7;
    wire \c0.n4745 ;
    wire \c0.n4746 ;
    wire data_8;
    wire bfn_15_27_0_;
    wire data_9;
    wire \c0.n4747 ;
    wire data_10;
    wire \c0.n4748 ;
    wire data_11;
    wire \c0.n4749 ;
    wire data_12;
    wire \c0.n4750 ;
    wire data_13;
    wire \c0.n4751 ;
    wire data_14;
    wire \c0.n4752 ;
    wire \c0.n4753 ;
    wire data_15;
    wire n1579;
    wire n5433;
    wire n4334;
    wire data_out_18_3;
    wire CLK_c;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__37951),
            .DIN(N__37950),
            .DOUT(N__37949),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__37951),
            .PADOUT(N__37950),
            .PADIN(N__37949),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__23712),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__37942),
            .DIN(N__37941),
            .DOUT(N__37940),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__37942),
            .PADOUT(N__37941),
            .PADIN(N__37940),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__37933),
            .DIN(N__37932),
            .DOUT(N__37931),
            .PACKAGEPIN(PIN_2));
    defparam rx_input_preio.PIN_TYPE=6'b000000;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__37933),
            .PADOUT(N__37932),
            .PADIN(N__37931),
            .CLOCKENABLE(VCCG0),
            .DIN0(\c0.rx.r_Rx_Data_R ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__37589),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx2_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx2_output_iopad.PULLUP=1'b1;
    IO_PAD tx2_output_iopad (
            .OE(N__37924),
            .DIN(N__37923),
            .DOUT(N__37922),
            .PACKAGEPIN(PIN_3));
    defparam tx2_output_preio.PIN_TYPE=6'b101001;
    defparam tx2_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx2_output_preio (
            .PADOEN(N__37924),
            .PADOUT(N__37923),
            .PADIN(N__37922),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12705),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__12675));
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__37915),
            .DIN(N__37914),
            .DOUT(N__37913),
            .PACKAGEPIN(PIN_1));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__37915),
            .PADOUT(N__37914),
            .PADIN(N__37913),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__28890),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15213));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__37906),
            .DIN(N__37905),
            .DOUT(N__37904),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__37906),
            .PADOUT(N__37905),
            .PADIN(N__37904),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__9582 (
            .O(N__37887),
            .I(N__37884));
    InMux I__9581 (
            .O(N__37884),
            .I(N__37881));
    LocalMux I__9580 (
            .O(N__37881),
            .I(N__37877));
    InMux I__9579 (
            .O(N__37880),
            .I(N__37874));
    Odrv12 I__9578 (
            .O(N__37877),
            .I(data_11));
    LocalMux I__9577 (
            .O(N__37874),
            .I(data_11));
    InMux I__9576 (
            .O(N__37869),
            .I(\c0.n4749 ));
    CascadeMux I__9575 (
            .O(N__37866),
            .I(N__37863));
    InMux I__9574 (
            .O(N__37863),
            .I(N__37860));
    LocalMux I__9573 (
            .O(N__37860),
            .I(N__37857));
    Span4Mux_h I__9572 (
            .O(N__37857),
            .I(N__37853));
    InMux I__9571 (
            .O(N__37856),
            .I(N__37850));
    Odrv4 I__9570 (
            .O(N__37853),
            .I(data_12));
    LocalMux I__9569 (
            .O(N__37850),
            .I(data_12));
    InMux I__9568 (
            .O(N__37845),
            .I(\c0.n4750 ));
    CascadeMux I__9567 (
            .O(N__37842),
            .I(N__37839));
    InMux I__9566 (
            .O(N__37839),
            .I(N__37836));
    LocalMux I__9565 (
            .O(N__37836),
            .I(N__37833));
    Span4Mux_h I__9564 (
            .O(N__37833),
            .I(N__37829));
    InMux I__9563 (
            .O(N__37832),
            .I(N__37826));
    Odrv4 I__9562 (
            .O(N__37829),
            .I(data_13));
    LocalMux I__9561 (
            .O(N__37826),
            .I(data_13));
    InMux I__9560 (
            .O(N__37821),
            .I(\c0.n4751 ));
    CascadeMux I__9559 (
            .O(N__37818),
            .I(N__37815));
    InMux I__9558 (
            .O(N__37815),
            .I(N__37812));
    LocalMux I__9557 (
            .O(N__37812),
            .I(N__37809));
    Span4Mux_v I__9556 (
            .O(N__37809),
            .I(N__37805));
    InMux I__9555 (
            .O(N__37808),
            .I(N__37802));
    Odrv4 I__9554 (
            .O(N__37805),
            .I(data_14));
    LocalMux I__9553 (
            .O(N__37802),
            .I(data_14));
    InMux I__9552 (
            .O(N__37797),
            .I(\c0.n4752 ));
    InMux I__9551 (
            .O(N__37794),
            .I(\c0.n4753 ));
    InMux I__9550 (
            .O(N__37791),
            .I(N__37787));
    InMux I__9549 (
            .O(N__37790),
            .I(N__37784));
    LocalMux I__9548 (
            .O(N__37787),
            .I(N__37781));
    LocalMux I__9547 (
            .O(N__37784),
            .I(data_15));
    Odrv12 I__9546 (
            .O(N__37781),
            .I(data_15));
    InMux I__9545 (
            .O(N__37776),
            .I(N__37773));
    LocalMux I__9544 (
            .O(N__37773),
            .I(N__37770));
    Span4Mux_v I__9543 (
            .O(N__37770),
            .I(N__37767));
    Odrv4 I__9542 (
            .O(N__37767),
            .I(n1579));
    CascadeMux I__9541 (
            .O(N__37764),
            .I(N__37761));
    InMux I__9540 (
            .O(N__37761),
            .I(N__37758));
    LocalMux I__9539 (
            .O(N__37758),
            .I(N__37754));
    CascadeMux I__9538 (
            .O(N__37757),
            .I(N__37751));
    Span4Mux_v I__9537 (
            .O(N__37754),
            .I(N__37748));
    InMux I__9536 (
            .O(N__37751),
            .I(N__37745));
    Span4Mux_h I__9535 (
            .O(N__37748),
            .I(N__37740));
    LocalMux I__9534 (
            .O(N__37745),
            .I(N__37740));
    Odrv4 I__9533 (
            .O(N__37740),
            .I(n5433));
    InMux I__9532 (
            .O(N__37737),
            .I(N__37731));
    InMux I__9531 (
            .O(N__37736),
            .I(N__37728));
    InMux I__9530 (
            .O(N__37735),
            .I(N__37721));
    InMux I__9529 (
            .O(N__37734),
            .I(N__37721));
    LocalMux I__9528 (
            .O(N__37731),
            .I(N__37718));
    LocalMux I__9527 (
            .O(N__37728),
            .I(N__37712));
    InMux I__9526 (
            .O(N__37727),
            .I(N__37709));
    InMux I__9525 (
            .O(N__37726),
            .I(N__37699));
    LocalMux I__9524 (
            .O(N__37721),
            .I(N__37696));
    Span4Mux_v I__9523 (
            .O(N__37718),
            .I(N__37693));
    InMux I__9522 (
            .O(N__37717),
            .I(N__37686));
    InMux I__9521 (
            .O(N__37716),
            .I(N__37686));
    InMux I__9520 (
            .O(N__37715),
            .I(N__37686));
    Span4Mux_h I__9519 (
            .O(N__37712),
            .I(N__37681));
    LocalMux I__9518 (
            .O(N__37709),
            .I(N__37681));
    InMux I__9517 (
            .O(N__37708),
            .I(N__37676));
    InMux I__9516 (
            .O(N__37707),
            .I(N__37676));
    InMux I__9515 (
            .O(N__37706),
            .I(N__37673));
    InMux I__9514 (
            .O(N__37705),
            .I(N__37666));
    InMux I__9513 (
            .O(N__37704),
            .I(N__37666));
    InMux I__9512 (
            .O(N__37703),
            .I(N__37666));
    InMux I__9511 (
            .O(N__37702),
            .I(N__37663));
    LocalMux I__9510 (
            .O(N__37699),
            .I(N__37658));
    Span4Mux_h I__9509 (
            .O(N__37696),
            .I(N__37658));
    Odrv4 I__9508 (
            .O(N__37693),
            .I(n4334));
    LocalMux I__9507 (
            .O(N__37686),
            .I(n4334));
    Odrv4 I__9506 (
            .O(N__37681),
            .I(n4334));
    LocalMux I__9505 (
            .O(N__37676),
            .I(n4334));
    LocalMux I__9504 (
            .O(N__37673),
            .I(n4334));
    LocalMux I__9503 (
            .O(N__37666),
            .I(n4334));
    LocalMux I__9502 (
            .O(N__37663),
            .I(n4334));
    Odrv4 I__9501 (
            .O(N__37658),
            .I(n4334));
    InMux I__9500 (
            .O(N__37641),
            .I(N__37638));
    LocalMux I__9499 (
            .O(N__37638),
            .I(N__37634));
    InMux I__9498 (
            .O(N__37637),
            .I(N__37631));
    Span4Mux_h I__9497 (
            .O(N__37634),
            .I(N__37628));
    LocalMux I__9496 (
            .O(N__37631),
            .I(data_out_18_3));
    Odrv4 I__9495 (
            .O(N__37628),
            .I(data_out_18_3));
    ClkMux I__9494 (
            .O(N__37623),
            .I(N__37137));
    ClkMux I__9493 (
            .O(N__37622),
            .I(N__37137));
    ClkMux I__9492 (
            .O(N__37621),
            .I(N__37137));
    ClkMux I__9491 (
            .O(N__37620),
            .I(N__37137));
    ClkMux I__9490 (
            .O(N__37619),
            .I(N__37137));
    ClkMux I__9489 (
            .O(N__37618),
            .I(N__37137));
    ClkMux I__9488 (
            .O(N__37617),
            .I(N__37137));
    ClkMux I__9487 (
            .O(N__37616),
            .I(N__37137));
    ClkMux I__9486 (
            .O(N__37615),
            .I(N__37137));
    ClkMux I__9485 (
            .O(N__37614),
            .I(N__37137));
    ClkMux I__9484 (
            .O(N__37613),
            .I(N__37137));
    ClkMux I__9483 (
            .O(N__37612),
            .I(N__37137));
    ClkMux I__9482 (
            .O(N__37611),
            .I(N__37137));
    ClkMux I__9481 (
            .O(N__37610),
            .I(N__37137));
    ClkMux I__9480 (
            .O(N__37609),
            .I(N__37137));
    ClkMux I__9479 (
            .O(N__37608),
            .I(N__37137));
    ClkMux I__9478 (
            .O(N__37607),
            .I(N__37137));
    ClkMux I__9477 (
            .O(N__37606),
            .I(N__37137));
    ClkMux I__9476 (
            .O(N__37605),
            .I(N__37137));
    ClkMux I__9475 (
            .O(N__37604),
            .I(N__37137));
    ClkMux I__9474 (
            .O(N__37603),
            .I(N__37137));
    ClkMux I__9473 (
            .O(N__37602),
            .I(N__37137));
    ClkMux I__9472 (
            .O(N__37601),
            .I(N__37137));
    ClkMux I__9471 (
            .O(N__37600),
            .I(N__37137));
    ClkMux I__9470 (
            .O(N__37599),
            .I(N__37137));
    ClkMux I__9469 (
            .O(N__37598),
            .I(N__37137));
    ClkMux I__9468 (
            .O(N__37597),
            .I(N__37137));
    ClkMux I__9467 (
            .O(N__37596),
            .I(N__37137));
    ClkMux I__9466 (
            .O(N__37595),
            .I(N__37137));
    ClkMux I__9465 (
            .O(N__37594),
            .I(N__37137));
    ClkMux I__9464 (
            .O(N__37593),
            .I(N__37137));
    ClkMux I__9463 (
            .O(N__37592),
            .I(N__37137));
    ClkMux I__9462 (
            .O(N__37591),
            .I(N__37137));
    ClkMux I__9461 (
            .O(N__37590),
            .I(N__37137));
    ClkMux I__9460 (
            .O(N__37589),
            .I(N__37137));
    ClkMux I__9459 (
            .O(N__37588),
            .I(N__37137));
    ClkMux I__9458 (
            .O(N__37587),
            .I(N__37137));
    ClkMux I__9457 (
            .O(N__37586),
            .I(N__37137));
    ClkMux I__9456 (
            .O(N__37585),
            .I(N__37137));
    ClkMux I__9455 (
            .O(N__37584),
            .I(N__37137));
    ClkMux I__9454 (
            .O(N__37583),
            .I(N__37137));
    ClkMux I__9453 (
            .O(N__37582),
            .I(N__37137));
    ClkMux I__9452 (
            .O(N__37581),
            .I(N__37137));
    ClkMux I__9451 (
            .O(N__37580),
            .I(N__37137));
    ClkMux I__9450 (
            .O(N__37579),
            .I(N__37137));
    ClkMux I__9449 (
            .O(N__37578),
            .I(N__37137));
    ClkMux I__9448 (
            .O(N__37577),
            .I(N__37137));
    ClkMux I__9447 (
            .O(N__37576),
            .I(N__37137));
    ClkMux I__9446 (
            .O(N__37575),
            .I(N__37137));
    ClkMux I__9445 (
            .O(N__37574),
            .I(N__37137));
    ClkMux I__9444 (
            .O(N__37573),
            .I(N__37137));
    ClkMux I__9443 (
            .O(N__37572),
            .I(N__37137));
    ClkMux I__9442 (
            .O(N__37571),
            .I(N__37137));
    ClkMux I__9441 (
            .O(N__37570),
            .I(N__37137));
    ClkMux I__9440 (
            .O(N__37569),
            .I(N__37137));
    ClkMux I__9439 (
            .O(N__37568),
            .I(N__37137));
    ClkMux I__9438 (
            .O(N__37567),
            .I(N__37137));
    ClkMux I__9437 (
            .O(N__37566),
            .I(N__37137));
    ClkMux I__9436 (
            .O(N__37565),
            .I(N__37137));
    ClkMux I__9435 (
            .O(N__37564),
            .I(N__37137));
    ClkMux I__9434 (
            .O(N__37563),
            .I(N__37137));
    ClkMux I__9433 (
            .O(N__37562),
            .I(N__37137));
    ClkMux I__9432 (
            .O(N__37561),
            .I(N__37137));
    ClkMux I__9431 (
            .O(N__37560),
            .I(N__37137));
    ClkMux I__9430 (
            .O(N__37559),
            .I(N__37137));
    ClkMux I__9429 (
            .O(N__37558),
            .I(N__37137));
    ClkMux I__9428 (
            .O(N__37557),
            .I(N__37137));
    ClkMux I__9427 (
            .O(N__37556),
            .I(N__37137));
    ClkMux I__9426 (
            .O(N__37555),
            .I(N__37137));
    ClkMux I__9425 (
            .O(N__37554),
            .I(N__37137));
    ClkMux I__9424 (
            .O(N__37553),
            .I(N__37137));
    ClkMux I__9423 (
            .O(N__37552),
            .I(N__37137));
    ClkMux I__9422 (
            .O(N__37551),
            .I(N__37137));
    ClkMux I__9421 (
            .O(N__37550),
            .I(N__37137));
    ClkMux I__9420 (
            .O(N__37549),
            .I(N__37137));
    ClkMux I__9419 (
            .O(N__37548),
            .I(N__37137));
    ClkMux I__9418 (
            .O(N__37547),
            .I(N__37137));
    ClkMux I__9417 (
            .O(N__37546),
            .I(N__37137));
    ClkMux I__9416 (
            .O(N__37545),
            .I(N__37137));
    ClkMux I__9415 (
            .O(N__37544),
            .I(N__37137));
    ClkMux I__9414 (
            .O(N__37543),
            .I(N__37137));
    ClkMux I__9413 (
            .O(N__37542),
            .I(N__37137));
    ClkMux I__9412 (
            .O(N__37541),
            .I(N__37137));
    ClkMux I__9411 (
            .O(N__37540),
            .I(N__37137));
    ClkMux I__9410 (
            .O(N__37539),
            .I(N__37137));
    ClkMux I__9409 (
            .O(N__37538),
            .I(N__37137));
    ClkMux I__9408 (
            .O(N__37537),
            .I(N__37137));
    ClkMux I__9407 (
            .O(N__37536),
            .I(N__37137));
    ClkMux I__9406 (
            .O(N__37535),
            .I(N__37137));
    ClkMux I__9405 (
            .O(N__37534),
            .I(N__37137));
    ClkMux I__9404 (
            .O(N__37533),
            .I(N__37137));
    ClkMux I__9403 (
            .O(N__37532),
            .I(N__37137));
    ClkMux I__9402 (
            .O(N__37531),
            .I(N__37137));
    ClkMux I__9401 (
            .O(N__37530),
            .I(N__37137));
    ClkMux I__9400 (
            .O(N__37529),
            .I(N__37137));
    ClkMux I__9399 (
            .O(N__37528),
            .I(N__37137));
    ClkMux I__9398 (
            .O(N__37527),
            .I(N__37137));
    ClkMux I__9397 (
            .O(N__37526),
            .I(N__37137));
    ClkMux I__9396 (
            .O(N__37525),
            .I(N__37137));
    ClkMux I__9395 (
            .O(N__37524),
            .I(N__37137));
    ClkMux I__9394 (
            .O(N__37523),
            .I(N__37137));
    ClkMux I__9393 (
            .O(N__37522),
            .I(N__37137));
    ClkMux I__9392 (
            .O(N__37521),
            .I(N__37137));
    ClkMux I__9391 (
            .O(N__37520),
            .I(N__37137));
    ClkMux I__9390 (
            .O(N__37519),
            .I(N__37137));
    ClkMux I__9389 (
            .O(N__37518),
            .I(N__37137));
    ClkMux I__9388 (
            .O(N__37517),
            .I(N__37137));
    ClkMux I__9387 (
            .O(N__37516),
            .I(N__37137));
    ClkMux I__9386 (
            .O(N__37515),
            .I(N__37137));
    ClkMux I__9385 (
            .O(N__37514),
            .I(N__37137));
    ClkMux I__9384 (
            .O(N__37513),
            .I(N__37137));
    ClkMux I__9383 (
            .O(N__37512),
            .I(N__37137));
    ClkMux I__9382 (
            .O(N__37511),
            .I(N__37137));
    ClkMux I__9381 (
            .O(N__37510),
            .I(N__37137));
    ClkMux I__9380 (
            .O(N__37509),
            .I(N__37137));
    ClkMux I__9379 (
            .O(N__37508),
            .I(N__37137));
    ClkMux I__9378 (
            .O(N__37507),
            .I(N__37137));
    ClkMux I__9377 (
            .O(N__37506),
            .I(N__37137));
    ClkMux I__9376 (
            .O(N__37505),
            .I(N__37137));
    ClkMux I__9375 (
            .O(N__37504),
            .I(N__37137));
    ClkMux I__9374 (
            .O(N__37503),
            .I(N__37137));
    ClkMux I__9373 (
            .O(N__37502),
            .I(N__37137));
    ClkMux I__9372 (
            .O(N__37501),
            .I(N__37137));
    ClkMux I__9371 (
            .O(N__37500),
            .I(N__37137));
    ClkMux I__9370 (
            .O(N__37499),
            .I(N__37137));
    ClkMux I__9369 (
            .O(N__37498),
            .I(N__37137));
    ClkMux I__9368 (
            .O(N__37497),
            .I(N__37137));
    ClkMux I__9367 (
            .O(N__37496),
            .I(N__37137));
    ClkMux I__9366 (
            .O(N__37495),
            .I(N__37137));
    ClkMux I__9365 (
            .O(N__37494),
            .I(N__37137));
    ClkMux I__9364 (
            .O(N__37493),
            .I(N__37137));
    ClkMux I__9363 (
            .O(N__37492),
            .I(N__37137));
    ClkMux I__9362 (
            .O(N__37491),
            .I(N__37137));
    ClkMux I__9361 (
            .O(N__37490),
            .I(N__37137));
    ClkMux I__9360 (
            .O(N__37489),
            .I(N__37137));
    ClkMux I__9359 (
            .O(N__37488),
            .I(N__37137));
    ClkMux I__9358 (
            .O(N__37487),
            .I(N__37137));
    ClkMux I__9357 (
            .O(N__37486),
            .I(N__37137));
    ClkMux I__9356 (
            .O(N__37485),
            .I(N__37137));
    ClkMux I__9355 (
            .O(N__37484),
            .I(N__37137));
    ClkMux I__9354 (
            .O(N__37483),
            .I(N__37137));
    ClkMux I__9353 (
            .O(N__37482),
            .I(N__37137));
    ClkMux I__9352 (
            .O(N__37481),
            .I(N__37137));
    ClkMux I__9351 (
            .O(N__37480),
            .I(N__37137));
    ClkMux I__9350 (
            .O(N__37479),
            .I(N__37137));
    ClkMux I__9349 (
            .O(N__37478),
            .I(N__37137));
    ClkMux I__9348 (
            .O(N__37477),
            .I(N__37137));
    ClkMux I__9347 (
            .O(N__37476),
            .I(N__37137));
    ClkMux I__9346 (
            .O(N__37475),
            .I(N__37137));
    ClkMux I__9345 (
            .O(N__37474),
            .I(N__37137));
    ClkMux I__9344 (
            .O(N__37473),
            .I(N__37137));
    ClkMux I__9343 (
            .O(N__37472),
            .I(N__37137));
    ClkMux I__9342 (
            .O(N__37471),
            .I(N__37137));
    ClkMux I__9341 (
            .O(N__37470),
            .I(N__37137));
    ClkMux I__9340 (
            .O(N__37469),
            .I(N__37137));
    ClkMux I__9339 (
            .O(N__37468),
            .I(N__37137));
    ClkMux I__9338 (
            .O(N__37467),
            .I(N__37137));
    ClkMux I__9337 (
            .O(N__37466),
            .I(N__37137));
    ClkMux I__9336 (
            .O(N__37465),
            .I(N__37137));
    ClkMux I__9335 (
            .O(N__37464),
            .I(N__37137));
    ClkMux I__9334 (
            .O(N__37463),
            .I(N__37137));
    ClkMux I__9333 (
            .O(N__37462),
            .I(N__37137));
    GlobalMux I__9332 (
            .O(N__37137),
            .I(N__37134));
    gio2CtrlBuf I__9331 (
            .O(N__37134),
            .I(CLK_c));
    CascadeMux I__9330 (
            .O(N__37131),
            .I(N__37128));
    InMux I__9329 (
            .O(N__37128),
            .I(N__37125));
    LocalMux I__9328 (
            .O(N__37125),
            .I(N__37121));
    InMux I__9327 (
            .O(N__37124),
            .I(N__37118));
    Odrv12 I__9326 (
            .O(N__37121),
            .I(data_3));
    LocalMux I__9325 (
            .O(N__37118),
            .I(data_3));
    InMux I__9324 (
            .O(N__37113),
            .I(\c0.n4741 ));
    CascadeMux I__9323 (
            .O(N__37110),
            .I(N__37107));
    InMux I__9322 (
            .O(N__37107),
            .I(N__37104));
    LocalMux I__9321 (
            .O(N__37104),
            .I(N__37101));
    Span4Mux_h I__9320 (
            .O(N__37101),
            .I(N__37097));
    InMux I__9319 (
            .O(N__37100),
            .I(N__37094));
    Odrv4 I__9318 (
            .O(N__37097),
            .I(data_4));
    LocalMux I__9317 (
            .O(N__37094),
            .I(data_4));
    InMux I__9316 (
            .O(N__37089),
            .I(\c0.n4742 ));
    CascadeMux I__9315 (
            .O(N__37086),
            .I(N__37083));
    InMux I__9314 (
            .O(N__37083),
            .I(N__37080));
    LocalMux I__9313 (
            .O(N__37080),
            .I(N__37076));
    InMux I__9312 (
            .O(N__37079),
            .I(N__37073));
    Odrv4 I__9311 (
            .O(N__37076),
            .I(data_5));
    LocalMux I__9310 (
            .O(N__37073),
            .I(data_5));
    InMux I__9309 (
            .O(N__37068),
            .I(\c0.n4743 ));
    CascadeMux I__9308 (
            .O(N__37065),
            .I(N__37062));
    InMux I__9307 (
            .O(N__37062),
            .I(N__37059));
    LocalMux I__9306 (
            .O(N__37059),
            .I(N__37055));
    InMux I__9305 (
            .O(N__37058),
            .I(N__37052));
    Odrv4 I__9304 (
            .O(N__37055),
            .I(data_6));
    LocalMux I__9303 (
            .O(N__37052),
            .I(data_6));
    InMux I__9302 (
            .O(N__37047),
            .I(\c0.n4744 ));
    CascadeMux I__9301 (
            .O(N__37044),
            .I(N__37041));
    InMux I__9300 (
            .O(N__37041),
            .I(N__37038));
    LocalMux I__9299 (
            .O(N__37038),
            .I(N__37034));
    InMux I__9298 (
            .O(N__37037),
            .I(N__37031));
    Odrv4 I__9297 (
            .O(N__37034),
            .I(data_7));
    LocalMux I__9296 (
            .O(N__37031),
            .I(data_7));
    InMux I__9295 (
            .O(N__37026),
            .I(\c0.n4745 ));
    InMux I__9294 (
            .O(N__37023),
            .I(N__37020));
    LocalMux I__9293 (
            .O(N__37020),
            .I(N__37016));
    InMux I__9292 (
            .O(N__37019),
            .I(N__37013));
    Odrv4 I__9291 (
            .O(N__37016),
            .I(data_8));
    LocalMux I__9290 (
            .O(N__37013),
            .I(data_8));
    InMux I__9289 (
            .O(N__37008),
            .I(bfn_15_27_0_));
    InMux I__9288 (
            .O(N__37005),
            .I(N__37002));
    LocalMux I__9287 (
            .O(N__37002),
            .I(N__36999));
    Span4Mux_h I__9286 (
            .O(N__36999),
            .I(N__36995));
    InMux I__9285 (
            .O(N__36998),
            .I(N__36992));
    Odrv4 I__9284 (
            .O(N__36995),
            .I(data_9));
    LocalMux I__9283 (
            .O(N__36992),
            .I(data_9));
    InMux I__9282 (
            .O(N__36987),
            .I(\c0.n4747 ));
    CascadeMux I__9281 (
            .O(N__36984),
            .I(N__36981));
    InMux I__9280 (
            .O(N__36981),
            .I(N__36977));
    InMux I__9279 (
            .O(N__36980),
            .I(N__36974));
    LocalMux I__9278 (
            .O(N__36977),
            .I(data_10));
    LocalMux I__9277 (
            .O(N__36974),
            .I(data_10));
    InMux I__9276 (
            .O(N__36969),
            .I(\c0.n4748 ));
    CascadeMux I__9275 (
            .O(N__36966),
            .I(N__36961));
    CascadeMux I__9274 (
            .O(N__36965),
            .I(N__36958));
    CascadeMux I__9273 (
            .O(N__36964),
            .I(N__36955));
    InMux I__9272 (
            .O(N__36961),
            .I(N__36949));
    InMux I__9271 (
            .O(N__36958),
            .I(N__36949));
    InMux I__9270 (
            .O(N__36955),
            .I(N__36946));
    InMux I__9269 (
            .O(N__36954),
            .I(N__36942));
    LocalMux I__9268 (
            .O(N__36949),
            .I(N__36939));
    LocalMux I__9267 (
            .O(N__36946),
            .I(N__36936));
    InMux I__9266 (
            .O(N__36945),
            .I(N__36932));
    LocalMux I__9265 (
            .O(N__36942),
            .I(N__36929));
    Span4Mux_h I__9264 (
            .O(N__36939),
            .I(N__36924));
    Span4Mux_h I__9263 (
            .O(N__36936),
            .I(N__36924));
    InMux I__9262 (
            .O(N__36935),
            .I(N__36921));
    LocalMux I__9261 (
            .O(N__36932),
            .I(data_out_11_2));
    Odrv4 I__9260 (
            .O(N__36929),
            .I(data_out_11_2));
    Odrv4 I__9259 (
            .O(N__36924),
            .I(data_out_11_2));
    LocalMux I__9258 (
            .O(N__36921),
            .I(data_out_11_2));
    CascadeMux I__9257 (
            .O(N__36912),
            .I(N__36906));
    CascadeMux I__9256 (
            .O(N__36911),
            .I(N__36903));
    InMux I__9255 (
            .O(N__36910),
            .I(N__36887));
    InMux I__9254 (
            .O(N__36909),
            .I(N__36887));
    InMux I__9253 (
            .O(N__36906),
            .I(N__36884));
    InMux I__9252 (
            .O(N__36903),
            .I(N__36877));
    InMux I__9251 (
            .O(N__36902),
            .I(N__36877));
    InMux I__9250 (
            .O(N__36901),
            .I(N__36877));
    InMux I__9249 (
            .O(N__36900),
            .I(N__36874));
    InMux I__9248 (
            .O(N__36899),
            .I(N__36871));
    InMux I__9247 (
            .O(N__36898),
            .I(N__36868));
    InMux I__9246 (
            .O(N__36897),
            .I(N__36865));
    InMux I__9245 (
            .O(N__36896),
            .I(N__36862));
    InMux I__9244 (
            .O(N__36895),
            .I(N__36855));
    InMux I__9243 (
            .O(N__36894),
            .I(N__36855));
    InMux I__9242 (
            .O(N__36893),
            .I(N__36855));
    InMux I__9241 (
            .O(N__36892),
            .I(N__36852));
    LocalMux I__9240 (
            .O(N__36887),
            .I(N__36849));
    LocalMux I__9239 (
            .O(N__36884),
            .I(N__36842));
    LocalMux I__9238 (
            .O(N__36877),
            .I(N__36842));
    LocalMux I__9237 (
            .O(N__36874),
            .I(N__36842));
    LocalMux I__9236 (
            .O(N__36871),
            .I(N__36837));
    LocalMux I__9235 (
            .O(N__36868),
            .I(N__36837));
    LocalMux I__9234 (
            .O(N__36865),
            .I(N__36832));
    LocalMux I__9233 (
            .O(N__36862),
            .I(N__36832));
    LocalMux I__9232 (
            .O(N__36855),
            .I(N__36829));
    LocalMux I__9231 (
            .O(N__36852),
            .I(N__36814));
    Span4Mux_h I__9230 (
            .O(N__36849),
            .I(N__36814));
    Span4Mux_v I__9229 (
            .O(N__36842),
            .I(N__36814));
    Span4Mux_v I__9228 (
            .O(N__36837),
            .I(N__36814));
    Span4Mux_v I__9227 (
            .O(N__36832),
            .I(N__36814));
    Span4Mux_h I__9226 (
            .O(N__36829),
            .I(N__36811));
    InMux I__9225 (
            .O(N__36828),
            .I(N__36806));
    InMux I__9224 (
            .O(N__36827),
            .I(N__36806));
    InMux I__9223 (
            .O(N__36826),
            .I(N__36801));
    InMux I__9222 (
            .O(N__36825),
            .I(N__36801));
    Odrv4 I__9221 (
            .O(N__36814),
            .I(n21_adj_1977));
    Odrv4 I__9220 (
            .O(N__36811),
            .I(n21_adj_1977));
    LocalMux I__9219 (
            .O(N__36806),
            .I(n21_adj_1977));
    LocalMux I__9218 (
            .O(N__36801),
            .I(n21_adj_1977));
    CascadeMux I__9217 (
            .O(N__36792),
            .I(N__36780));
    InMux I__9216 (
            .O(N__36791),
            .I(N__36777));
    InMux I__9215 (
            .O(N__36790),
            .I(N__36772));
    InMux I__9214 (
            .O(N__36789),
            .I(N__36772));
    InMux I__9213 (
            .O(N__36788),
            .I(N__36763));
    InMux I__9212 (
            .O(N__36787),
            .I(N__36763));
    InMux I__9211 (
            .O(N__36786),
            .I(N__36756));
    InMux I__9210 (
            .O(N__36785),
            .I(N__36756));
    InMux I__9209 (
            .O(N__36784),
            .I(N__36756));
    InMux I__9208 (
            .O(N__36783),
            .I(N__36753));
    InMux I__9207 (
            .O(N__36780),
            .I(N__36749));
    LocalMux I__9206 (
            .O(N__36777),
            .I(N__36745));
    LocalMux I__9205 (
            .O(N__36772),
            .I(N__36742));
    InMux I__9204 (
            .O(N__36771),
            .I(N__36733));
    InMux I__9203 (
            .O(N__36770),
            .I(N__36733));
    InMux I__9202 (
            .O(N__36769),
            .I(N__36733));
    InMux I__9201 (
            .O(N__36768),
            .I(N__36733));
    LocalMux I__9200 (
            .O(N__36763),
            .I(N__36724));
    LocalMux I__9199 (
            .O(N__36756),
            .I(N__36724));
    LocalMux I__9198 (
            .O(N__36753),
            .I(N__36724));
    InMux I__9197 (
            .O(N__36752),
            .I(N__36721));
    LocalMux I__9196 (
            .O(N__36749),
            .I(N__36718));
    InMux I__9195 (
            .O(N__36748),
            .I(N__36715));
    Span4Mux_v I__9194 (
            .O(N__36745),
            .I(N__36708));
    Span4Mux_h I__9193 (
            .O(N__36742),
            .I(N__36708));
    LocalMux I__9192 (
            .O(N__36733),
            .I(N__36708));
    InMux I__9191 (
            .O(N__36732),
            .I(N__36703));
    InMux I__9190 (
            .O(N__36731),
            .I(N__36703));
    Span4Mux_v I__9189 (
            .O(N__36724),
            .I(N__36696));
    LocalMux I__9188 (
            .O(N__36721),
            .I(N__36696));
    Span4Mux_v I__9187 (
            .O(N__36718),
            .I(N__36696));
    LocalMux I__9186 (
            .O(N__36715),
            .I(n4333));
    Odrv4 I__9185 (
            .O(N__36708),
            .I(n4333));
    LocalMux I__9184 (
            .O(N__36703),
            .I(n4333));
    Odrv4 I__9183 (
            .O(N__36696),
            .I(n4333));
    InMux I__9182 (
            .O(N__36687),
            .I(N__36684));
    LocalMux I__9181 (
            .O(N__36684),
            .I(N__36677));
    InMux I__9180 (
            .O(N__36683),
            .I(N__36674));
    InMux I__9179 (
            .O(N__36682),
            .I(N__36671));
    InMux I__9178 (
            .O(N__36681),
            .I(N__36668));
    InMux I__9177 (
            .O(N__36680),
            .I(N__36663));
    Span4Mux_v I__9176 (
            .O(N__36677),
            .I(N__36654));
    LocalMux I__9175 (
            .O(N__36674),
            .I(N__36654));
    LocalMux I__9174 (
            .O(N__36671),
            .I(N__36654));
    LocalMux I__9173 (
            .O(N__36668),
            .I(N__36654));
    InMux I__9172 (
            .O(N__36667),
            .I(N__36649));
    InMux I__9171 (
            .O(N__36666),
            .I(N__36649));
    LocalMux I__9170 (
            .O(N__36663),
            .I(data_out_10_1));
    Odrv4 I__9169 (
            .O(N__36654),
            .I(data_out_10_1));
    LocalMux I__9168 (
            .O(N__36649),
            .I(data_out_10_1));
    InMux I__9167 (
            .O(N__36642),
            .I(N__36636));
    InMux I__9166 (
            .O(N__36641),
            .I(N__36632));
    InMux I__9165 (
            .O(N__36640),
            .I(N__36629));
    InMux I__9164 (
            .O(N__36639),
            .I(N__36626));
    LocalMux I__9163 (
            .O(N__36636),
            .I(N__36623));
    InMux I__9162 (
            .O(N__36635),
            .I(N__36620));
    LocalMux I__9161 (
            .O(N__36632),
            .I(N__36615));
    LocalMux I__9160 (
            .O(N__36629),
            .I(N__36615));
    LocalMux I__9159 (
            .O(N__36626),
            .I(N__36609));
    Span4Mux_v I__9158 (
            .O(N__36623),
            .I(N__36609));
    LocalMux I__9157 (
            .O(N__36620),
            .I(N__36606));
    Span4Mux_h I__9156 (
            .O(N__36615),
            .I(N__36603));
    InMux I__9155 (
            .O(N__36614),
            .I(N__36600));
    Odrv4 I__9154 (
            .O(N__36609),
            .I(data_out_10_3));
    Odrv4 I__9153 (
            .O(N__36606),
            .I(data_out_10_3));
    Odrv4 I__9152 (
            .O(N__36603),
            .I(data_out_10_3));
    LocalMux I__9151 (
            .O(N__36600),
            .I(data_out_10_3));
    CascadeMux I__9150 (
            .O(N__36591),
            .I(N__36588));
    InMux I__9149 (
            .O(N__36588),
            .I(N__36584));
    CascadeMux I__9148 (
            .O(N__36587),
            .I(N__36581));
    LocalMux I__9147 (
            .O(N__36584),
            .I(N__36578));
    InMux I__9146 (
            .O(N__36581),
            .I(N__36575));
    Span4Mux_v I__9145 (
            .O(N__36578),
            .I(N__36570));
    LocalMux I__9144 (
            .O(N__36575),
            .I(N__36570));
    Odrv4 I__9143 (
            .O(N__36570),
            .I(n5424));
    InMux I__9142 (
            .O(N__36567),
            .I(N__36561));
    InMux I__9141 (
            .O(N__36566),
            .I(N__36558));
    InMux I__9140 (
            .O(N__36565),
            .I(N__36555));
    CascadeMux I__9139 (
            .O(N__36564),
            .I(N__36551));
    LocalMux I__9138 (
            .O(N__36561),
            .I(N__36547));
    LocalMux I__9137 (
            .O(N__36558),
            .I(N__36542));
    LocalMux I__9136 (
            .O(N__36555),
            .I(N__36542));
    InMux I__9135 (
            .O(N__36554),
            .I(N__36537));
    InMux I__9134 (
            .O(N__36551),
            .I(N__36537));
    InMux I__9133 (
            .O(N__36550),
            .I(N__36534));
    Span4Mux_h I__9132 (
            .O(N__36547),
            .I(N__36531));
    Span4Mux_h I__9131 (
            .O(N__36542),
            .I(N__36526));
    LocalMux I__9130 (
            .O(N__36537),
            .I(N__36526));
    LocalMux I__9129 (
            .O(N__36534),
            .I(data_out_11_0));
    Odrv4 I__9128 (
            .O(N__36531),
            .I(data_out_11_0));
    Odrv4 I__9127 (
            .O(N__36526),
            .I(data_out_11_0));
    CascadeMux I__9126 (
            .O(N__36519),
            .I(N__36515));
    InMux I__9125 (
            .O(N__36518),
            .I(N__36512));
    InMux I__9124 (
            .O(N__36515),
            .I(N__36509));
    LocalMux I__9123 (
            .O(N__36512),
            .I(N__36501));
    LocalMux I__9122 (
            .O(N__36509),
            .I(N__36501));
    CascadeMux I__9121 (
            .O(N__36508),
            .I(N__36496));
    InMux I__9120 (
            .O(N__36507),
            .I(N__36492));
    InMux I__9119 (
            .O(N__36506),
            .I(N__36489));
    Span4Mux_v I__9118 (
            .O(N__36501),
            .I(N__36486));
    CascadeMux I__9117 (
            .O(N__36500),
            .I(N__36483));
    InMux I__9116 (
            .O(N__36499),
            .I(N__36480));
    InMux I__9115 (
            .O(N__36496),
            .I(N__36475));
    InMux I__9114 (
            .O(N__36495),
            .I(N__36475));
    LocalMux I__9113 (
            .O(N__36492),
            .I(N__36472));
    LocalMux I__9112 (
            .O(N__36489),
            .I(N__36469));
    Span4Mux_h I__9111 (
            .O(N__36486),
            .I(N__36466));
    InMux I__9110 (
            .O(N__36483),
            .I(N__36463));
    LocalMux I__9109 (
            .O(N__36480),
            .I(N__36458));
    LocalMux I__9108 (
            .O(N__36475),
            .I(N__36458));
    Span4Mux_h I__9107 (
            .O(N__36472),
            .I(N__36455));
    Span4Mux_v I__9106 (
            .O(N__36469),
            .I(N__36450));
    Span4Mux_h I__9105 (
            .O(N__36466),
            .I(N__36450));
    LocalMux I__9104 (
            .O(N__36463),
            .I(data_out_10_7));
    Odrv4 I__9103 (
            .O(N__36458),
            .I(data_out_10_7));
    Odrv4 I__9102 (
            .O(N__36455),
            .I(data_out_10_7));
    Odrv4 I__9101 (
            .O(N__36450),
            .I(data_out_10_7));
    InMux I__9100 (
            .O(N__36441),
            .I(N__36437));
    InMux I__9099 (
            .O(N__36440),
            .I(N__36434));
    LocalMux I__9098 (
            .O(N__36437),
            .I(N__36431));
    LocalMux I__9097 (
            .O(N__36434),
            .I(N__36427));
    Span4Mux_h I__9096 (
            .O(N__36431),
            .I(N__36424));
    InMux I__9095 (
            .O(N__36430),
            .I(N__36421));
    Odrv4 I__9094 (
            .O(N__36427),
            .I(n5479));
    Odrv4 I__9093 (
            .O(N__36424),
            .I(n5479));
    LocalMux I__9092 (
            .O(N__36421),
            .I(n5479));
    CascadeMux I__9091 (
            .O(N__36414),
            .I(N__36409));
    InMux I__9090 (
            .O(N__36413),
            .I(N__36403));
    InMux I__9089 (
            .O(N__36412),
            .I(N__36403));
    InMux I__9088 (
            .O(N__36409),
            .I(N__36400));
    InMux I__9087 (
            .O(N__36408),
            .I(N__36396));
    LocalMux I__9086 (
            .O(N__36403),
            .I(N__36393));
    LocalMux I__9085 (
            .O(N__36400),
            .I(N__36387));
    InMux I__9084 (
            .O(N__36399),
            .I(N__36384));
    LocalMux I__9083 (
            .O(N__36396),
            .I(N__36381));
    Span4Mux_h I__9082 (
            .O(N__36393),
            .I(N__36378));
    InMux I__9081 (
            .O(N__36392),
            .I(N__36371));
    InMux I__9080 (
            .O(N__36391),
            .I(N__36371));
    InMux I__9079 (
            .O(N__36390),
            .I(N__36371));
    Span4Mux_h I__9078 (
            .O(N__36387),
            .I(N__36368));
    LocalMux I__9077 (
            .O(N__36384),
            .I(data_out_11_3));
    Odrv4 I__9076 (
            .O(N__36381),
            .I(data_out_11_3));
    Odrv4 I__9075 (
            .O(N__36378),
            .I(data_out_11_3));
    LocalMux I__9074 (
            .O(N__36371),
            .I(data_out_11_3));
    Odrv4 I__9073 (
            .O(N__36368),
            .I(data_out_11_3));
    InMux I__9072 (
            .O(N__36357),
            .I(N__36354));
    LocalMux I__9071 (
            .O(N__36354),
            .I(n8_adj_1984));
    CascadeMux I__9070 (
            .O(N__36351),
            .I(n7_adj_1985_cascade_));
    CascadeMux I__9069 (
            .O(N__36348),
            .I(N__36345));
    InMux I__9068 (
            .O(N__36345),
            .I(N__36342));
    LocalMux I__9067 (
            .O(N__36342),
            .I(N__36338));
    InMux I__9066 (
            .O(N__36341),
            .I(N__36335));
    Span4Mux_h I__9065 (
            .O(N__36338),
            .I(N__36332));
    LocalMux I__9064 (
            .O(N__36335),
            .I(data_out_19_1));
    Odrv4 I__9063 (
            .O(N__36332),
            .I(data_out_19_1));
    CascadeMux I__9062 (
            .O(N__36327),
            .I(N__36324));
    InMux I__9061 (
            .O(N__36324),
            .I(N__36321));
    LocalMux I__9060 (
            .O(N__36321),
            .I(N__36318));
    Span4Mux_h I__9059 (
            .O(N__36318),
            .I(N__36314));
    InMux I__9058 (
            .O(N__36317),
            .I(N__36311));
    Odrv4 I__9057 (
            .O(N__36314),
            .I(data_0));
    LocalMux I__9056 (
            .O(N__36311),
            .I(data_0));
    InMux I__9055 (
            .O(N__36306),
            .I(bfn_15_26_0_));
    InMux I__9054 (
            .O(N__36303),
            .I(N__36300));
    LocalMux I__9053 (
            .O(N__36300),
            .I(N__36297));
    Span4Mux_h I__9052 (
            .O(N__36297),
            .I(N__36293));
    InMux I__9051 (
            .O(N__36296),
            .I(N__36290));
    Odrv4 I__9050 (
            .O(N__36293),
            .I(data_1));
    LocalMux I__9049 (
            .O(N__36290),
            .I(data_1));
    InMux I__9048 (
            .O(N__36285),
            .I(\c0.n4739 ));
    CascadeMux I__9047 (
            .O(N__36282),
            .I(N__36279));
    InMux I__9046 (
            .O(N__36279),
            .I(N__36276));
    LocalMux I__9045 (
            .O(N__36276),
            .I(N__36272));
    InMux I__9044 (
            .O(N__36275),
            .I(N__36269));
    Odrv4 I__9043 (
            .O(N__36272),
            .I(data_2));
    LocalMux I__9042 (
            .O(N__36269),
            .I(data_2));
    InMux I__9041 (
            .O(N__36264),
            .I(\c0.n4740 ));
    CascadeMux I__9040 (
            .O(N__36261),
            .I(N__36257));
    InMux I__9039 (
            .O(N__36260),
            .I(N__36252));
    InMux I__9038 (
            .O(N__36257),
            .I(N__36252));
    LocalMux I__9037 (
            .O(N__36252),
            .I(N__36249));
    Span4Mux_h I__9036 (
            .O(N__36249),
            .I(N__36245));
    InMux I__9035 (
            .O(N__36248),
            .I(N__36242));
    Odrv4 I__9034 (
            .O(N__36245),
            .I(blink_counter_23));
    LocalMux I__9033 (
            .O(N__36242),
            .I(blink_counter_23));
    InMux I__9032 (
            .O(N__36237),
            .I(n4732));
    CascadeMux I__9031 (
            .O(N__36234),
            .I(N__36231));
    InMux I__9030 (
            .O(N__36231),
            .I(N__36225));
    InMux I__9029 (
            .O(N__36230),
            .I(N__36225));
    LocalMux I__9028 (
            .O(N__36225),
            .I(N__36222));
    Span12Mux_h I__9027 (
            .O(N__36222),
            .I(N__36218));
    InMux I__9026 (
            .O(N__36221),
            .I(N__36215));
    Odrv12 I__9025 (
            .O(N__36218),
            .I(blink_counter_24));
    LocalMux I__9024 (
            .O(N__36215),
            .I(blink_counter_24));
    InMux I__9023 (
            .O(N__36210),
            .I(bfn_14_28_0_));
    InMux I__9022 (
            .O(N__36207),
            .I(n4734));
    InMux I__9021 (
            .O(N__36204),
            .I(N__36201));
    LocalMux I__9020 (
            .O(N__36201),
            .I(N__36198));
    Span4Mux_h I__9019 (
            .O(N__36198),
            .I(N__36195));
    Span4Mux_v I__9018 (
            .O(N__36195),
            .I(N__36191));
    InMux I__9017 (
            .O(N__36194),
            .I(N__36188));
    Odrv4 I__9016 (
            .O(N__36191),
            .I(blink_counter_25));
    LocalMux I__9015 (
            .O(N__36188),
            .I(blink_counter_25));
    CascadeMux I__9014 (
            .O(N__36183),
            .I(N__36180));
    InMux I__9013 (
            .O(N__36180),
            .I(N__36177));
    LocalMux I__9012 (
            .O(N__36177),
            .I(N__36170));
    InMux I__9011 (
            .O(N__36176),
            .I(N__36166));
    InMux I__9010 (
            .O(N__36175),
            .I(N__36163));
    InMux I__9009 (
            .O(N__36174),
            .I(N__36160));
    InMux I__9008 (
            .O(N__36173),
            .I(N__36157));
    Span4Mux_v I__9007 (
            .O(N__36170),
            .I(N__36154));
    InMux I__9006 (
            .O(N__36169),
            .I(N__36151));
    LocalMux I__9005 (
            .O(N__36166),
            .I(N__36147));
    LocalMux I__9004 (
            .O(N__36163),
            .I(N__36140));
    LocalMux I__9003 (
            .O(N__36160),
            .I(N__36140));
    LocalMux I__9002 (
            .O(N__36157),
            .I(N__36140));
    Span4Mux_h I__9001 (
            .O(N__36154),
            .I(N__36135));
    LocalMux I__9000 (
            .O(N__36151),
            .I(N__36135));
    InMux I__8999 (
            .O(N__36150),
            .I(N__36132));
    Span4Mux_h I__8998 (
            .O(N__36147),
            .I(N__36125));
    Span4Mux_v I__8997 (
            .O(N__36140),
            .I(N__36125));
    Span4Mux_h I__8996 (
            .O(N__36135),
            .I(N__36125));
    LocalMux I__8995 (
            .O(N__36132),
            .I(data_out_10_2));
    Odrv4 I__8994 (
            .O(N__36125),
            .I(data_out_10_2));
    InMux I__8993 (
            .O(N__36120),
            .I(N__36116));
    InMux I__8992 (
            .O(N__36119),
            .I(N__36113));
    LocalMux I__8991 (
            .O(N__36116),
            .I(N__36105));
    LocalMux I__8990 (
            .O(N__36113),
            .I(N__36102));
    InMux I__8989 (
            .O(N__36112),
            .I(N__36097));
    InMux I__8988 (
            .O(N__36111),
            .I(N__36097));
    InMux I__8987 (
            .O(N__36110),
            .I(N__36094));
    InMux I__8986 (
            .O(N__36109),
            .I(N__36089));
    InMux I__8985 (
            .O(N__36108),
            .I(N__36089));
    Span4Mux_v I__8984 (
            .O(N__36105),
            .I(N__36082));
    Span4Mux_h I__8983 (
            .O(N__36102),
            .I(N__36082));
    LocalMux I__8982 (
            .O(N__36097),
            .I(N__36082));
    LocalMux I__8981 (
            .O(N__36094),
            .I(data_out_11_6));
    LocalMux I__8980 (
            .O(N__36089),
            .I(data_out_11_6));
    Odrv4 I__8979 (
            .O(N__36082),
            .I(data_out_11_6));
    CascadeMux I__8978 (
            .O(N__36075),
            .I(N__36065));
    InMux I__8977 (
            .O(N__36074),
            .I(N__36059));
    CascadeMux I__8976 (
            .O(N__36073),
            .I(N__36049));
    InMux I__8975 (
            .O(N__36072),
            .I(N__36040));
    InMux I__8974 (
            .O(N__36071),
            .I(N__36035));
    InMux I__8973 (
            .O(N__36070),
            .I(N__36035));
    InMux I__8972 (
            .O(N__36069),
            .I(N__36032));
    InMux I__8971 (
            .O(N__36068),
            .I(N__36025));
    InMux I__8970 (
            .O(N__36065),
            .I(N__36025));
    InMux I__8969 (
            .O(N__36064),
            .I(N__36025));
    CascadeMux I__8968 (
            .O(N__36063),
            .I(N__36016));
    InMux I__8967 (
            .O(N__36062),
            .I(N__36011));
    LocalMux I__8966 (
            .O(N__36059),
            .I(N__36008));
    InMux I__8965 (
            .O(N__36058),
            .I(N__36001));
    InMux I__8964 (
            .O(N__36057),
            .I(N__36001));
    InMux I__8963 (
            .O(N__36056),
            .I(N__36001));
    InMux I__8962 (
            .O(N__36055),
            .I(N__35992));
    InMux I__8961 (
            .O(N__36054),
            .I(N__35992));
    InMux I__8960 (
            .O(N__36053),
            .I(N__35992));
    InMux I__8959 (
            .O(N__36052),
            .I(N__35987));
    InMux I__8958 (
            .O(N__36049),
            .I(N__35987));
    InMux I__8957 (
            .O(N__36048),
            .I(N__35984));
    InMux I__8956 (
            .O(N__36047),
            .I(N__35971));
    InMux I__8955 (
            .O(N__36046),
            .I(N__35966));
    InMux I__8954 (
            .O(N__36045),
            .I(N__35966));
    InMux I__8953 (
            .O(N__36044),
            .I(N__35957));
    InMux I__8952 (
            .O(N__36043),
            .I(N__35957));
    LocalMux I__8951 (
            .O(N__36040),
            .I(N__35948));
    LocalMux I__8950 (
            .O(N__36035),
            .I(N__35948));
    LocalMux I__8949 (
            .O(N__36032),
            .I(N__35948));
    LocalMux I__8948 (
            .O(N__36025),
            .I(N__35948));
    InMux I__8947 (
            .O(N__36024),
            .I(N__35945));
    CascadeMux I__8946 (
            .O(N__36023),
            .I(N__35936));
    CascadeMux I__8945 (
            .O(N__36022),
            .I(N__35920));
    InMux I__8944 (
            .O(N__36021),
            .I(N__35911));
    InMux I__8943 (
            .O(N__36020),
            .I(N__35911));
    InMux I__8942 (
            .O(N__36019),
            .I(N__35911));
    InMux I__8941 (
            .O(N__36016),
            .I(N__35908));
    InMux I__8940 (
            .O(N__36015),
            .I(N__35894));
    InMux I__8939 (
            .O(N__36014),
            .I(N__35894));
    LocalMux I__8938 (
            .O(N__36011),
            .I(N__35887));
    Span4Mux_v I__8937 (
            .O(N__36008),
            .I(N__35887));
    LocalMux I__8936 (
            .O(N__36001),
            .I(N__35887));
    InMux I__8935 (
            .O(N__36000),
            .I(N__35884));
    InMux I__8934 (
            .O(N__35999),
            .I(N__35881));
    LocalMux I__8933 (
            .O(N__35992),
            .I(N__35869));
    LocalMux I__8932 (
            .O(N__35987),
            .I(N__35869));
    LocalMux I__8931 (
            .O(N__35984),
            .I(N__35869));
    InMux I__8930 (
            .O(N__35983),
            .I(N__35862));
    InMux I__8929 (
            .O(N__35982),
            .I(N__35862));
    InMux I__8928 (
            .O(N__35981),
            .I(N__35862));
    InMux I__8927 (
            .O(N__35980),
            .I(N__35857));
    InMux I__8926 (
            .O(N__35979),
            .I(N__35857));
    InMux I__8925 (
            .O(N__35978),
            .I(N__35854));
    InMux I__8924 (
            .O(N__35977),
            .I(N__35850));
    InMux I__8923 (
            .O(N__35976),
            .I(N__35847));
    InMux I__8922 (
            .O(N__35975),
            .I(N__35844));
    InMux I__8921 (
            .O(N__35974),
            .I(N__35841));
    LocalMux I__8920 (
            .O(N__35971),
            .I(N__35836));
    LocalMux I__8919 (
            .O(N__35966),
            .I(N__35836));
    InMux I__8918 (
            .O(N__35965),
            .I(N__35831));
    InMux I__8917 (
            .O(N__35964),
            .I(N__35831));
    CascadeMux I__8916 (
            .O(N__35963),
            .I(N__35813));
    InMux I__8915 (
            .O(N__35962),
            .I(N__35809));
    LocalMux I__8914 (
            .O(N__35957),
            .I(N__35802));
    Span4Mux_v I__8913 (
            .O(N__35948),
            .I(N__35802));
    LocalMux I__8912 (
            .O(N__35945),
            .I(N__35802));
    InMux I__8911 (
            .O(N__35944),
            .I(N__35797));
    InMux I__8910 (
            .O(N__35943),
            .I(N__35797));
    InMux I__8909 (
            .O(N__35942),
            .I(N__35792));
    InMux I__8908 (
            .O(N__35941),
            .I(N__35792));
    InMux I__8907 (
            .O(N__35940),
            .I(N__35789));
    InMux I__8906 (
            .O(N__35939),
            .I(N__35782));
    InMux I__8905 (
            .O(N__35936),
            .I(N__35782));
    InMux I__8904 (
            .O(N__35935),
            .I(N__35782));
    InMux I__8903 (
            .O(N__35934),
            .I(N__35775));
    InMux I__8902 (
            .O(N__35933),
            .I(N__35775));
    InMux I__8901 (
            .O(N__35932),
            .I(N__35775));
    InMux I__8900 (
            .O(N__35931),
            .I(N__35766));
    InMux I__8899 (
            .O(N__35930),
            .I(N__35766));
    InMux I__8898 (
            .O(N__35929),
            .I(N__35766));
    InMux I__8897 (
            .O(N__35928),
            .I(N__35766));
    InMux I__8896 (
            .O(N__35927),
            .I(N__35761));
    InMux I__8895 (
            .O(N__35926),
            .I(N__35761));
    InMux I__8894 (
            .O(N__35925),
            .I(N__35757));
    InMux I__8893 (
            .O(N__35924),
            .I(N__35754));
    InMux I__8892 (
            .O(N__35923),
            .I(N__35751));
    InMux I__8891 (
            .O(N__35920),
            .I(N__35744));
    InMux I__8890 (
            .O(N__35919),
            .I(N__35744));
    InMux I__8889 (
            .O(N__35918),
            .I(N__35744));
    LocalMux I__8888 (
            .O(N__35911),
            .I(N__35741));
    LocalMux I__8887 (
            .O(N__35908),
            .I(N__35738));
    InMux I__8886 (
            .O(N__35907),
            .I(N__35731));
    InMux I__8885 (
            .O(N__35906),
            .I(N__35731));
    InMux I__8884 (
            .O(N__35905),
            .I(N__35731));
    InMux I__8883 (
            .O(N__35904),
            .I(N__35728));
    InMux I__8882 (
            .O(N__35903),
            .I(N__35725));
    InMux I__8881 (
            .O(N__35902),
            .I(N__35720));
    InMux I__8880 (
            .O(N__35901),
            .I(N__35720));
    InMux I__8879 (
            .O(N__35900),
            .I(N__35716));
    InMux I__8878 (
            .O(N__35899),
            .I(N__35713));
    LocalMux I__8877 (
            .O(N__35894),
            .I(N__35704));
    Span4Mux_v I__8876 (
            .O(N__35887),
            .I(N__35704));
    LocalMux I__8875 (
            .O(N__35884),
            .I(N__35704));
    LocalMux I__8874 (
            .O(N__35881),
            .I(N__35704));
    InMux I__8873 (
            .O(N__35880),
            .I(N__35699));
    InMux I__8872 (
            .O(N__35879),
            .I(N__35699));
    InMux I__8871 (
            .O(N__35878),
            .I(N__35694));
    InMux I__8870 (
            .O(N__35877),
            .I(N__35694));
    CascadeMux I__8869 (
            .O(N__35876),
            .I(N__35690));
    Span4Mux_v I__8868 (
            .O(N__35869),
            .I(N__35674));
    LocalMux I__8867 (
            .O(N__35862),
            .I(N__35674));
    LocalMux I__8866 (
            .O(N__35857),
            .I(N__35674));
    LocalMux I__8865 (
            .O(N__35854),
            .I(N__35671));
    InMux I__8864 (
            .O(N__35853),
            .I(N__35668));
    LocalMux I__8863 (
            .O(N__35850),
            .I(N__35659));
    LocalMux I__8862 (
            .O(N__35847),
            .I(N__35659));
    LocalMux I__8861 (
            .O(N__35844),
            .I(N__35659));
    LocalMux I__8860 (
            .O(N__35841),
            .I(N__35659));
    Span4Mux_v I__8859 (
            .O(N__35836),
            .I(N__35654));
    LocalMux I__8858 (
            .O(N__35831),
            .I(N__35654));
    InMux I__8857 (
            .O(N__35830),
            .I(N__35651));
    InMux I__8856 (
            .O(N__35829),
            .I(N__35642));
    InMux I__8855 (
            .O(N__35828),
            .I(N__35642));
    InMux I__8854 (
            .O(N__35827),
            .I(N__35642));
    InMux I__8853 (
            .O(N__35826),
            .I(N__35642));
    CascadeMux I__8852 (
            .O(N__35825),
            .I(N__35637));
    InMux I__8851 (
            .O(N__35824),
            .I(N__35623));
    InMux I__8850 (
            .O(N__35823),
            .I(N__35623));
    InMux I__8849 (
            .O(N__35822),
            .I(N__35616));
    InMux I__8848 (
            .O(N__35821),
            .I(N__35616));
    InMux I__8847 (
            .O(N__35820),
            .I(N__35616));
    InMux I__8846 (
            .O(N__35819),
            .I(N__35607));
    InMux I__8845 (
            .O(N__35818),
            .I(N__35607));
    InMux I__8844 (
            .O(N__35817),
            .I(N__35607));
    InMux I__8843 (
            .O(N__35816),
            .I(N__35607));
    InMux I__8842 (
            .O(N__35813),
            .I(N__35604));
    InMux I__8841 (
            .O(N__35812),
            .I(N__35601));
    LocalMux I__8840 (
            .O(N__35809),
            .I(N__35594));
    Span4Mux_v I__8839 (
            .O(N__35802),
            .I(N__35594));
    LocalMux I__8838 (
            .O(N__35797),
            .I(N__35594));
    LocalMux I__8837 (
            .O(N__35792),
            .I(N__35591));
    LocalMux I__8836 (
            .O(N__35789),
            .I(N__35584));
    LocalMux I__8835 (
            .O(N__35782),
            .I(N__35584));
    LocalMux I__8834 (
            .O(N__35775),
            .I(N__35584));
    LocalMux I__8833 (
            .O(N__35766),
            .I(N__35581));
    LocalMux I__8832 (
            .O(N__35761),
            .I(N__35578));
    InMux I__8831 (
            .O(N__35760),
            .I(N__35575));
    LocalMux I__8830 (
            .O(N__35757),
            .I(N__35570));
    LocalMux I__8829 (
            .O(N__35754),
            .I(N__35570));
    LocalMux I__8828 (
            .O(N__35751),
            .I(N__35559));
    LocalMux I__8827 (
            .O(N__35744),
            .I(N__35559));
    Span4Mux_v I__8826 (
            .O(N__35741),
            .I(N__35559));
    Span4Mux_v I__8825 (
            .O(N__35738),
            .I(N__35559));
    LocalMux I__8824 (
            .O(N__35731),
            .I(N__35559));
    LocalMux I__8823 (
            .O(N__35728),
            .I(N__35550));
    LocalMux I__8822 (
            .O(N__35725),
            .I(N__35550));
    LocalMux I__8821 (
            .O(N__35720),
            .I(N__35550));
    InMux I__8820 (
            .O(N__35719),
            .I(N__35547));
    LocalMux I__8819 (
            .O(N__35716),
            .I(N__35536));
    LocalMux I__8818 (
            .O(N__35713),
            .I(N__35536));
    Span4Mux_h I__8817 (
            .O(N__35704),
            .I(N__35536));
    LocalMux I__8816 (
            .O(N__35699),
            .I(N__35536));
    LocalMux I__8815 (
            .O(N__35694),
            .I(N__35536));
    InMux I__8814 (
            .O(N__35693),
            .I(N__35533));
    InMux I__8813 (
            .O(N__35690),
            .I(N__35524));
    InMux I__8812 (
            .O(N__35689),
            .I(N__35524));
    InMux I__8811 (
            .O(N__35688),
            .I(N__35524));
    InMux I__8810 (
            .O(N__35687),
            .I(N__35524));
    InMux I__8809 (
            .O(N__35686),
            .I(N__35519));
    InMux I__8808 (
            .O(N__35685),
            .I(N__35519));
    CascadeMux I__8807 (
            .O(N__35684),
            .I(N__35512));
    InMux I__8806 (
            .O(N__35683),
            .I(N__35506));
    InMux I__8805 (
            .O(N__35682),
            .I(N__35503));
    InMux I__8804 (
            .O(N__35681),
            .I(N__35496));
    Span4Mux_h I__8803 (
            .O(N__35674),
            .I(N__35489));
    Span4Mux_v I__8802 (
            .O(N__35671),
            .I(N__35489));
    LocalMux I__8801 (
            .O(N__35668),
            .I(N__35489));
    Span4Mux_v I__8800 (
            .O(N__35659),
            .I(N__35486));
    Span4Mux_v I__8799 (
            .O(N__35654),
            .I(N__35479));
    LocalMux I__8798 (
            .O(N__35651),
            .I(N__35479));
    LocalMux I__8797 (
            .O(N__35642),
            .I(N__35479));
    InMux I__8796 (
            .O(N__35641),
            .I(N__35474));
    InMux I__8795 (
            .O(N__35640),
            .I(N__35471));
    InMux I__8794 (
            .O(N__35637),
            .I(N__35466));
    InMux I__8793 (
            .O(N__35636),
            .I(N__35466));
    InMux I__8792 (
            .O(N__35635),
            .I(N__35457));
    InMux I__8791 (
            .O(N__35634),
            .I(N__35457));
    InMux I__8790 (
            .O(N__35633),
            .I(N__35457));
    InMux I__8789 (
            .O(N__35632),
            .I(N__35457));
    InMux I__8788 (
            .O(N__35631),
            .I(N__35454));
    InMux I__8787 (
            .O(N__35630),
            .I(N__35451));
    InMux I__8786 (
            .O(N__35629),
            .I(N__35443));
    InMux I__8785 (
            .O(N__35628),
            .I(N__35443));
    LocalMux I__8784 (
            .O(N__35623),
            .I(N__35436));
    LocalMux I__8783 (
            .O(N__35616),
            .I(N__35436));
    LocalMux I__8782 (
            .O(N__35607),
            .I(N__35436));
    LocalMux I__8781 (
            .O(N__35604),
            .I(N__35433));
    LocalMux I__8780 (
            .O(N__35601),
            .I(N__35430));
    Span4Mux_v I__8779 (
            .O(N__35594),
            .I(N__35427));
    Span4Mux_s3_h I__8778 (
            .O(N__35591),
            .I(N__35422));
    Span4Mux_v I__8777 (
            .O(N__35584),
            .I(N__35422));
    Span4Mux_v I__8776 (
            .O(N__35581),
            .I(N__35419));
    Span4Mux_v I__8775 (
            .O(N__35578),
            .I(N__35416));
    LocalMux I__8774 (
            .O(N__35575),
            .I(N__35413));
    Span4Mux_v I__8773 (
            .O(N__35570),
            .I(N__35408));
    Span4Mux_v I__8772 (
            .O(N__35559),
            .I(N__35408));
    CascadeMux I__8771 (
            .O(N__35558),
            .I(N__35402));
    InMux I__8770 (
            .O(N__35557),
            .I(N__35398));
    Span4Mux_v I__8769 (
            .O(N__35550),
            .I(N__35385));
    LocalMux I__8768 (
            .O(N__35547),
            .I(N__35385));
    Span4Mux_v I__8767 (
            .O(N__35536),
            .I(N__35385));
    LocalMux I__8766 (
            .O(N__35533),
            .I(N__35385));
    LocalMux I__8765 (
            .O(N__35524),
            .I(N__35385));
    LocalMux I__8764 (
            .O(N__35519),
            .I(N__35385));
    InMux I__8763 (
            .O(N__35518),
            .I(N__35381));
    InMux I__8762 (
            .O(N__35517),
            .I(N__35378));
    InMux I__8761 (
            .O(N__35516),
            .I(N__35373));
    InMux I__8760 (
            .O(N__35515),
            .I(N__35373));
    InMux I__8759 (
            .O(N__35512),
            .I(N__35368));
    InMux I__8758 (
            .O(N__35511),
            .I(N__35368));
    InMux I__8757 (
            .O(N__35510),
            .I(N__35363));
    InMux I__8756 (
            .O(N__35509),
            .I(N__35363));
    LocalMux I__8755 (
            .O(N__35506),
            .I(N__35358));
    LocalMux I__8754 (
            .O(N__35503),
            .I(N__35358));
    InMux I__8753 (
            .O(N__35502),
            .I(N__35353));
    InMux I__8752 (
            .O(N__35501),
            .I(N__35353));
    InMux I__8751 (
            .O(N__35500),
            .I(N__35350));
    InMux I__8750 (
            .O(N__35499),
            .I(N__35339));
    LocalMux I__8749 (
            .O(N__35496),
            .I(N__35330));
    Span4Mux_h I__8748 (
            .O(N__35489),
            .I(N__35330));
    Span4Mux_s1_h I__8747 (
            .O(N__35486),
            .I(N__35330));
    Span4Mux_v I__8746 (
            .O(N__35479),
            .I(N__35330));
    InMux I__8745 (
            .O(N__35478),
            .I(N__35325));
    InMux I__8744 (
            .O(N__35477),
            .I(N__35325));
    LocalMux I__8743 (
            .O(N__35474),
            .I(N__35322));
    LocalMux I__8742 (
            .O(N__35471),
            .I(N__35311));
    LocalMux I__8741 (
            .O(N__35466),
            .I(N__35311));
    LocalMux I__8740 (
            .O(N__35457),
            .I(N__35311));
    LocalMux I__8739 (
            .O(N__35454),
            .I(N__35311));
    LocalMux I__8738 (
            .O(N__35451),
            .I(N__35311));
    InMux I__8737 (
            .O(N__35450),
            .I(N__35306));
    InMux I__8736 (
            .O(N__35449),
            .I(N__35306));
    InMux I__8735 (
            .O(N__35448),
            .I(N__35303));
    LocalMux I__8734 (
            .O(N__35443),
            .I(N__35296));
    Span4Mux_h I__8733 (
            .O(N__35436),
            .I(N__35296));
    Span4Mux_v I__8732 (
            .O(N__35433),
            .I(N__35296));
    Span4Mux_h I__8731 (
            .O(N__35430),
            .I(N__35289));
    Span4Mux_v I__8730 (
            .O(N__35427),
            .I(N__35289));
    Span4Mux_v I__8729 (
            .O(N__35422),
            .I(N__35289));
    Span4Mux_v I__8728 (
            .O(N__35419),
            .I(N__35284));
    Span4Mux_v I__8727 (
            .O(N__35416),
            .I(N__35284));
    Span4Mux_v I__8726 (
            .O(N__35413),
            .I(N__35279));
    Span4Mux_v I__8725 (
            .O(N__35408),
            .I(N__35279));
    InMux I__8724 (
            .O(N__35407),
            .I(N__35270));
    InMux I__8723 (
            .O(N__35406),
            .I(N__35270));
    InMux I__8722 (
            .O(N__35405),
            .I(N__35270));
    InMux I__8721 (
            .O(N__35402),
            .I(N__35270));
    InMux I__8720 (
            .O(N__35401),
            .I(N__35267));
    LocalMux I__8719 (
            .O(N__35398),
            .I(N__35262));
    Span4Mux_h I__8718 (
            .O(N__35385),
            .I(N__35262));
    InMux I__8717 (
            .O(N__35384),
            .I(N__35252));
    LocalMux I__8716 (
            .O(N__35381),
            .I(N__35245));
    LocalMux I__8715 (
            .O(N__35378),
            .I(N__35245));
    LocalMux I__8714 (
            .O(N__35373),
            .I(N__35245));
    LocalMux I__8713 (
            .O(N__35368),
            .I(N__35242));
    LocalMux I__8712 (
            .O(N__35363),
            .I(N__35237));
    Span4Mux_v I__8711 (
            .O(N__35358),
            .I(N__35237));
    LocalMux I__8710 (
            .O(N__35353),
            .I(N__35234));
    LocalMux I__8709 (
            .O(N__35350),
            .I(N__35231));
    InMux I__8708 (
            .O(N__35349),
            .I(N__35228));
    InMux I__8707 (
            .O(N__35348),
            .I(N__35225));
    InMux I__8706 (
            .O(N__35347),
            .I(N__35220));
    InMux I__8705 (
            .O(N__35346),
            .I(N__35220));
    InMux I__8704 (
            .O(N__35345),
            .I(N__35211));
    InMux I__8703 (
            .O(N__35344),
            .I(N__35211));
    InMux I__8702 (
            .O(N__35343),
            .I(N__35211));
    InMux I__8701 (
            .O(N__35342),
            .I(N__35211));
    LocalMux I__8700 (
            .O(N__35339),
            .I(N__35208));
    Sp12to4 I__8699 (
            .O(N__35330),
            .I(N__35205));
    LocalMux I__8698 (
            .O(N__35325),
            .I(N__35196));
    Sp12to4 I__8697 (
            .O(N__35322),
            .I(N__35196));
    Span12Mux_h I__8696 (
            .O(N__35311),
            .I(N__35196));
    LocalMux I__8695 (
            .O(N__35306),
            .I(N__35196));
    LocalMux I__8694 (
            .O(N__35303),
            .I(N__35185));
    Span4Mux_v I__8693 (
            .O(N__35296),
            .I(N__35185));
    Span4Mux_v I__8692 (
            .O(N__35289),
            .I(N__35185));
    Span4Mux_v I__8691 (
            .O(N__35284),
            .I(N__35185));
    Span4Mux_h I__8690 (
            .O(N__35279),
            .I(N__35185));
    LocalMux I__8689 (
            .O(N__35270),
            .I(N__35178));
    LocalMux I__8688 (
            .O(N__35267),
            .I(N__35178));
    Sp12to4 I__8687 (
            .O(N__35262),
            .I(N__35178));
    InMux I__8686 (
            .O(N__35261),
            .I(N__35175));
    InMux I__8685 (
            .O(N__35260),
            .I(N__35170));
    InMux I__8684 (
            .O(N__35259),
            .I(N__35170));
    InMux I__8683 (
            .O(N__35258),
            .I(N__35163));
    InMux I__8682 (
            .O(N__35257),
            .I(N__35163));
    InMux I__8681 (
            .O(N__35256),
            .I(N__35163));
    InMux I__8680 (
            .O(N__35255),
            .I(N__35160));
    LocalMux I__8679 (
            .O(N__35252),
            .I(N__35157));
    Span4Mux_v I__8678 (
            .O(N__35245),
            .I(N__35154));
    Span4Mux_v I__8677 (
            .O(N__35242),
            .I(N__35145));
    Span4Mux_s1_h I__8676 (
            .O(N__35237),
            .I(N__35145));
    Span4Mux_v I__8675 (
            .O(N__35234),
            .I(N__35145));
    Span4Mux_v I__8674 (
            .O(N__35231),
            .I(N__35145));
    LocalMux I__8673 (
            .O(N__35228),
            .I(N__35132));
    LocalMux I__8672 (
            .O(N__35225),
            .I(N__35132));
    LocalMux I__8671 (
            .O(N__35220),
            .I(N__35132));
    LocalMux I__8670 (
            .O(N__35211),
            .I(N__35132));
    Span12Mux_h I__8669 (
            .O(N__35208),
            .I(N__35132));
    Span12Mux_s4_h I__8668 (
            .O(N__35205),
            .I(N__35132));
    Span12Mux_v I__8667 (
            .O(N__35196),
            .I(N__35129));
    Sp12to4 I__8666 (
            .O(N__35185),
            .I(N__35124));
    Span12Mux_v I__8665 (
            .O(N__35178),
            .I(N__35124));
    LocalMux I__8664 (
            .O(N__35175),
            .I(rx_data_ready));
    LocalMux I__8663 (
            .O(N__35170),
            .I(rx_data_ready));
    LocalMux I__8662 (
            .O(N__35163),
            .I(rx_data_ready));
    LocalMux I__8661 (
            .O(N__35160),
            .I(rx_data_ready));
    Odrv4 I__8660 (
            .O(N__35157),
            .I(rx_data_ready));
    Odrv4 I__8659 (
            .O(N__35154),
            .I(rx_data_ready));
    Odrv4 I__8658 (
            .O(N__35145),
            .I(rx_data_ready));
    Odrv12 I__8657 (
            .O(N__35132),
            .I(rx_data_ready));
    Odrv12 I__8656 (
            .O(N__35129),
            .I(rx_data_ready));
    Odrv12 I__8655 (
            .O(N__35124),
            .I(rx_data_ready));
    CascadeMux I__8654 (
            .O(N__35103),
            .I(N__35100));
    InMux I__8653 (
            .O(N__35100),
            .I(N__35096));
    InMux I__8652 (
            .O(N__35099),
            .I(N__35093));
    LocalMux I__8651 (
            .O(N__35096),
            .I(N__35090));
    LocalMux I__8650 (
            .O(N__35093),
            .I(N__35087));
    Span4Mux_v I__8649 (
            .O(N__35090),
            .I(N__35081));
    Span4Mux_v I__8648 (
            .O(N__35087),
            .I(N__35081));
    InMux I__8647 (
            .O(N__35086),
            .I(N__35078));
    Odrv4 I__8646 (
            .O(N__35081),
            .I(data_in_16_0));
    LocalMux I__8645 (
            .O(N__35078),
            .I(data_in_16_0));
    CascadeMux I__8644 (
            .O(N__35073),
            .I(N__35070));
    InMux I__8643 (
            .O(N__35070),
            .I(N__35066));
    InMux I__8642 (
            .O(N__35069),
            .I(N__35063));
    LocalMux I__8641 (
            .O(N__35066),
            .I(N__35060));
    LocalMux I__8640 (
            .O(N__35063),
            .I(N__35057));
    Span4Mux_v I__8639 (
            .O(N__35060),
            .I(N__35052));
    Span4Mux_h I__8638 (
            .O(N__35057),
            .I(N__35052));
    Span4Mux_h I__8637 (
            .O(N__35052),
            .I(N__35048));
    InMux I__8636 (
            .O(N__35051),
            .I(N__35045));
    Odrv4 I__8635 (
            .O(N__35048),
            .I(data_in_15_0));
    LocalMux I__8634 (
            .O(N__35045),
            .I(data_in_15_0));
    InMux I__8633 (
            .O(N__35040),
            .I(N__35031));
    InMux I__8632 (
            .O(N__35039),
            .I(N__35031));
    InMux I__8631 (
            .O(N__35038),
            .I(N__35031));
    LocalMux I__8630 (
            .O(N__35031),
            .I(N__35028));
    Span4Mux_h I__8629 (
            .O(N__35028),
            .I(N__35025));
    Span4Mux_h I__8628 (
            .O(N__35025),
            .I(N__35022));
    Odrv4 I__8627 (
            .O(N__35022),
            .I(\c0.n5409 ));
    InMux I__8626 (
            .O(N__35019),
            .I(N__35015));
    CascadeMux I__8625 (
            .O(N__35018),
            .I(N__35009));
    LocalMux I__8624 (
            .O(N__35015),
            .I(N__35004));
    InMux I__8623 (
            .O(N__35014),
            .I(N__35001));
    InMux I__8622 (
            .O(N__35013),
            .I(N__34998));
    InMux I__8621 (
            .O(N__35012),
            .I(N__34993));
    InMux I__8620 (
            .O(N__35009),
            .I(N__34993));
    InMux I__8619 (
            .O(N__35008),
            .I(N__34988));
    InMux I__8618 (
            .O(N__35007),
            .I(N__34988));
    Span4Mux_h I__8617 (
            .O(N__35004),
            .I(N__34983));
    LocalMux I__8616 (
            .O(N__35001),
            .I(N__34983));
    LocalMux I__8615 (
            .O(N__34998),
            .I(data_out_11_1));
    LocalMux I__8614 (
            .O(N__34993),
            .I(data_out_11_1));
    LocalMux I__8613 (
            .O(N__34988),
            .I(data_out_11_1));
    Odrv4 I__8612 (
            .O(N__34983),
            .I(data_out_11_1));
    CascadeMux I__8611 (
            .O(N__34974),
            .I(\c0.n5409_cascade_ ));
    InMux I__8610 (
            .O(N__34971),
            .I(N__34963));
    InMux I__8609 (
            .O(N__34970),
            .I(N__34963));
    CascadeMux I__8608 (
            .O(N__34969),
            .I(N__34958));
    CascadeMux I__8607 (
            .O(N__34968),
            .I(N__34955));
    LocalMux I__8606 (
            .O(N__34963),
            .I(N__34952));
    InMux I__8605 (
            .O(N__34962),
            .I(N__34949));
    InMux I__8604 (
            .O(N__34961),
            .I(N__34946));
    InMux I__8603 (
            .O(N__34958),
            .I(N__34940));
    InMux I__8602 (
            .O(N__34955),
            .I(N__34940));
    Span4Mux_h I__8601 (
            .O(N__34952),
            .I(N__34937));
    LocalMux I__8600 (
            .O(N__34949),
            .I(N__34932));
    LocalMux I__8599 (
            .O(N__34946),
            .I(N__34932));
    InMux I__8598 (
            .O(N__34945),
            .I(N__34929));
    LocalMux I__8597 (
            .O(N__34940),
            .I(N__34926));
    Odrv4 I__8596 (
            .O(N__34937),
            .I(data_out_11_4));
    Odrv4 I__8595 (
            .O(N__34932),
            .I(data_out_11_4));
    LocalMux I__8594 (
            .O(N__34929),
            .I(data_out_11_4));
    Odrv4 I__8593 (
            .O(N__34926),
            .I(data_out_11_4));
    InMux I__8592 (
            .O(N__34917),
            .I(N__34914));
    LocalMux I__8591 (
            .O(N__34914),
            .I(N__34911));
    Span4Mux_h I__8590 (
            .O(N__34911),
            .I(N__34908));
    Odrv4 I__8589 (
            .O(N__34908),
            .I(n4_adj_1978));
    CascadeMux I__8588 (
            .O(N__34905),
            .I(N__34902));
    InMux I__8587 (
            .O(N__34902),
            .I(N__34899));
    LocalMux I__8586 (
            .O(N__34899),
            .I(N__34896));
    Span4Mux_v I__8585 (
            .O(N__34896),
            .I(N__34893));
    Odrv4 I__8584 (
            .O(N__34893),
            .I(n4_adj_1983));
    InMux I__8583 (
            .O(N__34890),
            .I(N__34887));
    LocalMux I__8582 (
            .O(N__34887),
            .I(n11));
    InMux I__8581 (
            .O(N__34884),
            .I(n4724));
    InMux I__8580 (
            .O(N__34881),
            .I(N__34878));
    LocalMux I__8579 (
            .O(N__34878),
            .I(n10));
    InMux I__8578 (
            .O(N__34875),
            .I(bfn_14_27_0_));
    InMux I__8577 (
            .O(N__34872),
            .I(N__34869));
    LocalMux I__8576 (
            .O(N__34869),
            .I(n9));
    InMux I__8575 (
            .O(N__34866),
            .I(n4726));
    InMux I__8574 (
            .O(N__34863),
            .I(N__34860));
    LocalMux I__8573 (
            .O(N__34860),
            .I(n8));
    InMux I__8572 (
            .O(N__34857),
            .I(n4727));
    InMux I__8571 (
            .O(N__34854),
            .I(N__34851));
    LocalMux I__8570 (
            .O(N__34851),
            .I(n7));
    InMux I__8569 (
            .O(N__34848),
            .I(n4728));
    InMux I__8568 (
            .O(N__34845),
            .I(N__34842));
    LocalMux I__8567 (
            .O(N__34842),
            .I(n6));
    InMux I__8566 (
            .O(N__34839),
            .I(n4729));
    InMux I__8565 (
            .O(N__34836),
            .I(N__34830));
    InMux I__8564 (
            .O(N__34835),
            .I(N__34830));
    LocalMux I__8563 (
            .O(N__34830),
            .I(N__34827));
    Span4Mux_v I__8562 (
            .O(N__34827),
            .I(N__34824));
    Span4Mux_h I__8561 (
            .O(N__34824),
            .I(N__34820));
    InMux I__8560 (
            .O(N__34823),
            .I(N__34817));
    Odrv4 I__8559 (
            .O(N__34820),
            .I(blink_counter_21));
    LocalMux I__8558 (
            .O(N__34817),
            .I(blink_counter_21));
    InMux I__8557 (
            .O(N__34812),
            .I(n4730));
    InMux I__8556 (
            .O(N__34809),
            .I(N__34803));
    InMux I__8555 (
            .O(N__34808),
            .I(N__34803));
    LocalMux I__8554 (
            .O(N__34803),
            .I(N__34800));
    Span4Mux_v I__8553 (
            .O(N__34800),
            .I(N__34797));
    Sp12to4 I__8552 (
            .O(N__34797),
            .I(N__34793));
    InMux I__8551 (
            .O(N__34796),
            .I(N__34790));
    Odrv12 I__8550 (
            .O(N__34793),
            .I(blink_counter_22));
    LocalMux I__8549 (
            .O(N__34790),
            .I(blink_counter_22));
    InMux I__8548 (
            .O(N__34785),
            .I(n4731));
    InMux I__8547 (
            .O(N__34782),
            .I(n4715));
    InMux I__8546 (
            .O(N__34779),
            .I(N__34776));
    LocalMux I__8545 (
            .O(N__34776),
            .I(n19));
    InMux I__8544 (
            .O(N__34773),
            .I(n4716));
    InMux I__8543 (
            .O(N__34770),
            .I(N__34767));
    LocalMux I__8542 (
            .O(N__34767),
            .I(n18));
    InMux I__8541 (
            .O(N__34764),
            .I(bfn_14_26_0_));
    InMux I__8540 (
            .O(N__34761),
            .I(N__34758));
    LocalMux I__8539 (
            .O(N__34758),
            .I(n17));
    InMux I__8538 (
            .O(N__34755),
            .I(n4718));
    InMux I__8537 (
            .O(N__34752),
            .I(N__34749));
    LocalMux I__8536 (
            .O(N__34749),
            .I(n16));
    InMux I__8535 (
            .O(N__34746),
            .I(n4719));
    InMux I__8534 (
            .O(N__34743),
            .I(N__34740));
    LocalMux I__8533 (
            .O(N__34740),
            .I(n15));
    InMux I__8532 (
            .O(N__34737),
            .I(n4720));
    InMux I__8531 (
            .O(N__34734),
            .I(N__34731));
    LocalMux I__8530 (
            .O(N__34731),
            .I(n14));
    InMux I__8529 (
            .O(N__34728),
            .I(n4721));
    InMux I__8528 (
            .O(N__34725),
            .I(N__34722));
    LocalMux I__8527 (
            .O(N__34722),
            .I(n13));
    InMux I__8526 (
            .O(N__34719),
            .I(n4722));
    InMux I__8525 (
            .O(N__34716),
            .I(N__34713));
    LocalMux I__8524 (
            .O(N__34713),
            .I(n12));
    InMux I__8523 (
            .O(N__34710),
            .I(n4723));
    InMux I__8522 (
            .O(N__34707),
            .I(N__34702));
    InMux I__8521 (
            .O(N__34706),
            .I(N__34697));
    InMux I__8520 (
            .O(N__34705),
            .I(N__34697));
    LocalMux I__8519 (
            .O(N__34702),
            .I(N__34691));
    LocalMux I__8518 (
            .O(N__34697),
            .I(N__34688));
    InMux I__8517 (
            .O(N__34696),
            .I(N__34683));
    InMux I__8516 (
            .O(N__34695),
            .I(N__34683));
    InMux I__8515 (
            .O(N__34694),
            .I(N__34679));
    Span4Mux_v I__8514 (
            .O(N__34691),
            .I(N__34676));
    Span4Mux_v I__8513 (
            .O(N__34688),
            .I(N__34671));
    LocalMux I__8512 (
            .O(N__34683),
            .I(N__34671));
    InMux I__8511 (
            .O(N__34682),
            .I(N__34668));
    LocalMux I__8510 (
            .O(N__34679),
            .I(data_out_11_5));
    Odrv4 I__8509 (
            .O(N__34676),
            .I(data_out_11_5));
    Odrv4 I__8508 (
            .O(N__34671),
            .I(data_out_11_5));
    LocalMux I__8507 (
            .O(N__34668),
            .I(data_out_11_5));
    InMux I__8506 (
            .O(N__34659),
            .I(N__34654));
    InMux I__8505 (
            .O(N__34658),
            .I(N__34651));
    InMux I__8504 (
            .O(N__34657),
            .I(N__34646));
    LocalMux I__8503 (
            .O(N__34654),
            .I(N__34643));
    LocalMux I__8502 (
            .O(N__34651),
            .I(N__34638));
    InMux I__8501 (
            .O(N__34650),
            .I(N__34635));
    InMux I__8500 (
            .O(N__34649),
            .I(N__34632));
    LocalMux I__8499 (
            .O(N__34646),
            .I(N__34629));
    Span4Mux_v I__8498 (
            .O(N__34643),
            .I(N__34626));
    InMux I__8497 (
            .O(N__34642),
            .I(N__34621));
    InMux I__8496 (
            .O(N__34641),
            .I(N__34621));
    Span4Mux_h I__8495 (
            .O(N__34638),
            .I(N__34618));
    LocalMux I__8494 (
            .O(N__34635),
            .I(N__34613));
    LocalMux I__8493 (
            .O(N__34632),
            .I(N__34613));
    Odrv12 I__8492 (
            .O(N__34629),
            .I(data_out_10_6));
    Odrv4 I__8491 (
            .O(N__34626),
            .I(data_out_10_6));
    LocalMux I__8490 (
            .O(N__34621),
            .I(data_out_10_6));
    Odrv4 I__8489 (
            .O(N__34618),
            .I(data_out_10_6));
    Odrv4 I__8488 (
            .O(N__34613),
            .I(data_out_10_6));
    InMux I__8487 (
            .O(N__34602),
            .I(N__34599));
    LocalMux I__8486 (
            .O(N__34599),
            .I(N__34596));
    Odrv12 I__8485 (
            .O(N__34596),
            .I(n4_adj_1976));
    InMux I__8484 (
            .O(N__34593),
            .I(N__34590));
    LocalMux I__8483 (
            .O(N__34590),
            .I(n26));
    InMux I__8482 (
            .O(N__34587),
            .I(bfn_14_25_0_));
    InMux I__8481 (
            .O(N__34584),
            .I(N__34581));
    LocalMux I__8480 (
            .O(N__34581),
            .I(n25));
    InMux I__8479 (
            .O(N__34578),
            .I(n4710));
    InMux I__8478 (
            .O(N__34575),
            .I(N__34572));
    LocalMux I__8477 (
            .O(N__34572),
            .I(n24));
    InMux I__8476 (
            .O(N__34569),
            .I(n4711));
    InMux I__8475 (
            .O(N__34566),
            .I(N__34563));
    LocalMux I__8474 (
            .O(N__34563),
            .I(n23));
    InMux I__8473 (
            .O(N__34560),
            .I(n4712));
    InMux I__8472 (
            .O(N__34557),
            .I(N__34554));
    LocalMux I__8471 (
            .O(N__34554),
            .I(n22));
    InMux I__8470 (
            .O(N__34551),
            .I(n4713));
    InMux I__8469 (
            .O(N__34548),
            .I(N__34545));
    LocalMux I__8468 (
            .O(N__34545),
            .I(n21));
    InMux I__8467 (
            .O(N__34542),
            .I(n4714));
    InMux I__8466 (
            .O(N__34539),
            .I(N__34536));
    LocalMux I__8465 (
            .O(N__34536),
            .I(n20));
    InMux I__8464 (
            .O(N__34533),
            .I(N__34528));
    InMux I__8463 (
            .O(N__34532),
            .I(N__34525));
    InMux I__8462 (
            .O(N__34531),
            .I(N__34522));
    LocalMux I__8461 (
            .O(N__34528),
            .I(N__34515));
    LocalMux I__8460 (
            .O(N__34525),
            .I(N__34512));
    LocalMux I__8459 (
            .O(N__34522),
            .I(N__34509));
    InMux I__8458 (
            .O(N__34521),
            .I(N__34500));
    InMux I__8457 (
            .O(N__34520),
            .I(N__34500));
    InMux I__8456 (
            .O(N__34519),
            .I(N__34500));
    InMux I__8455 (
            .O(N__34518),
            .I(N__34500));
    Odrv4 I__8454 (
            .O(N__34515),
            .I(data_out_11_7));
    Odrv4 I__8453 (
            .O(N__34512),
            .I(data_out_11_7));
    Odrv4 I__8452 (
            .O(N__34509),
            .I(data_out_11_7));
    LocalMux I__8451 (
            .O(N__34500),
            .I(data_out_11_7));
    CascadeMux I__8450 (
            .O(N__34491),
            .I(N__34488));
    InMux I__8449 (
            .O(N__34488),
            .I(N__34485));
    LocalMux I__8448 (
            .O(N__34485),
            .I(N__34482));
    Span4Mux_h I__8447 (
            .O(N__34482),
            .I(N__34479));
    Span4Mux_h I__8446 (
            .O(N__34479),
            .I(N__34474));
    InMux I__8445 (
            .O(N__34478),
            .I(N__34471));
    InMux I__8444 (
            .O(N__34477),
            .I(N__34468));
    Odrv4 I__8443 (
            .O(N__34474),
            .I(data_in_13_5));
    LocalMux I__8442 (
            .O(N__34471),
            .I(data_in_13_5));
    LocalMux I__8441 (
            .O(N__34468),
            .I(data_in_13_5));
    CascadeMux I__8440 (
            .O(N__34461),
            .I(N__34458));
    InMux I__8439 (
            .O(N__34458),
            .I(N__34454));
    InMux I__8438 (
            .O(N__34457),
            .I(N__34451));
    LocalMux I__8437 (
            .O(N__34454),
            .I(N__34448));
    LocalMux I__8436 (
            .O(N__34451),
            .I(N__34445));
    Span4Mux_h I__8435 (
            .O(N__34448),
            .I(N__34439));
    Span4Mux_h I__8434 (
            .O(N__34445),
            .I(N__34439));
    InMux I__8433 (
            .O(N__34444),
            .I(N__34436));
    Odrv4 I__8432 (
            .O(N__34439),
            .I(data_in_12_5));
    LocalMux I__8431 (
            .O(N__34436),
            .I(data_in_12_5));
    InMux I__8430 (
            .O(N__34431),
            .I(N__34426));
    InMux I__8429 (
            .O(N__34430),
            .I(N__34423));
    InMux I__8428 (
            .O(N__34429),
            .I(N__34420));
    LocalMux I__8427 (
            .O(N__34426),
            .I(N__34412));
    LocalMux I__8426 (
            .O(N__34423),
            .I(N__34412));
    LocalMux I__8425 (
            .O(N__34420),
            .I(N__34412));
    InMux I__8424 (
            .O(N__34419),
            .I(N__34408));
    Span4Mux_v I__8423 (
            .O(N__34412),
            .I(N__34405));
    InMux I__8422 (
            .O(N__34411),
            .I(N__34402));
    LocalMux I__8421 (
            .O(N__34408),
            .I(data_out_10_5));
    Odrv4 I__8420 (
            .O(N__34405),
            .I(data_out_10_5));
    LocalMux I__8419 (
            .O(N__34402),
            .I(data_out_10_5));
    CascadeMux I__8418 (
            .O(N__34395),
            .I(N__34392));
    InMux I__8417 (
            .O(N__34392),
            .I(N__34389));
    LocalMux I__8416 (
            .O(N__34389),
            .I(N__34386));
    Odrv4 I__8415 (
            .O(N__34386),
            .I(\c0.n9_adj_1911 ));
    CascadeMux I__8414 (
            .O(N__34383),
            .I(N__34376));
    InMux I__8413 (
            .O(N__34382),
            .I(N__34370));
    InMux I__8412 (
            .O(N__34381),
            .I(N__34370));
    InMux I__8411 (
            .O(N__34380),
            .I(N__34367));
    InMux I__8410 (
            .O(N__34379),
            .I(N__34364));
    InMux I__8409 (
            .O(N__34376),
            .I(N__34361));
    InMux I__8408 (
            .O(N__34375),
            .I(N__34358));
    LocalMux I__8407 (
            .O(N__34370),
            .I(N__34355));
    LocalMux I__8406 (
            .O(N__34367),
            .I(N__34352));
    LocalMux I__8405 (
            .O(N__34364),
            .I(N__34349));
    LocalMux I__8404 (
            .O(N__34361),
            .I(N__34342));
    LocalMux I__8403 (
            .O(N__34358),
            .I(N__34342));
    Span4Mux_h I__8402 (
            .O(N__34355),
            .I(N__34342));
    Span4Mux_h I__8401 (
            .O(N__34352),
            .I(N__34339));
    Odrv4 I__8400 (
            .O(N__34349),
            .I(data_out_10_0));
    Odrv4 I__8399 (
            .O(N__34342),
            .I(data_out_10_0));
    Odrv4 I__8398 (
            .O(N__34339),
            .I(data_out_10_0));
    InMux I__8397 (
            .O(N__34332),
            .I(N__34316));
    InMux I__8396 (
            .O(N__34331),
            .I(N__34309));
    InMux I__8395 (
            .O(N__34330),
            .I(N__34309));
    InMux I__8394 (
            .O(N__34329),
            .I(N__34309));
    InMux I__8393 (
            .O(N__34328),
            .I(N__34304));
    InMux I__8392 (
            .O(N__34327),
            .I(N__34304));
    InMux I__8391 (
            .O(N__34326),
            .I(N__34296));
    InMux I__8390 (
            .O(N__34325),
            .I(N__34296));
    InMux I__8389 (
            .O(N__34324),
            .I(N__34291));
    InMux I__8388 (
            .O(N__34323),
            .I(N__34291));
    InMux I__8387 (
            .O(N__34322),
            .I(N__34286));
    InMux I__8386 (
            .O(N__34321),
            .I(N__34286));
    InMux I__8385 (
            .O(N__34320),
            .I(N__34283));
    InMux I__8384 (
            .O(N__34319),
            .I(N__34280));
    LocalMux I__8383 (
            .O(N__34316),
            .I(N__34271));
    LocalMux I__8382 (
            .O(N__34309),
            .I(N__34271));
    LocalMux I__8381 (
            .O(N__34304),
            .I(N__34271));
    InMux I__8380 (
            .O(N__34303),
            .I(N__34262));
    InMux I__8379 (
            .O(N__34302),
            .I(N__34262));
    InMux I__8378 (
            .O(N__34301),
            .I(N__34262));
    LocalMux I__8377 (
            .O(N__34296),
            .I(N__34257));
    LocalMux I__8376 (
            .O(N__34291),
            .I(N__34257));
    LocalMux I__8375 (
            .O(N__34286),
            .I(N__34250));
    LocalMux I__8374 (
            .O(N__34283),
            .I(N__34250));
    LocalMux I__8373 (
            .O(N__34280),
            .I(N__34250));
    InMux I__8372 (
            .O(N__34279),
            .I(N__34247));
    CascadeMux I__8371 (
            .O(N__34278),
            .I(N__34244));
    Span4Mux_v I__8370 (
            .O(N__34271),
            .I(N__34241));
    InMux I__8369 (
            .O(N__34270),
            .I(N__34238));
    InMux I__8368 (
            .O(N__34269),
            .I(N__34235));
    LocalMux I__8367 (
            .O(N__34262),
            .I(N__34226));
    Span4Mux_h I__8366 (
            .O(N__34257),
            .I(N__34226));
    Span4Mux_v I__8365 (
            .O(N__34250),
            .I(N__34226));
    LocalMux I__8364 (
            .O(N__34247),
            .I(N__34226));
    InMux I__8363 (
            .O(N__34244),
            .I(N__34223));
    Odrv4 I__8362 (
            .O(N__34241),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__8361 (
            .O(N__34238),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__8360 (
            .O(N__34235),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__8359 (
            .O(N__34226),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__8358 (
            .O(N__34223),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__8357 (
            .O(N__34212),
            .I(N__34208));
    InMux I__8356 (
            .O(N__34211),
            .I(N__34201));
    LocalMux I__8355 (
            .O(N__34208),
            .I(N__34198));
    InMux I__8354 (
            .O(N__34207),
            .I(N__34188));
    InMux I__8353 (
            .O(N__34206),
            .I(N__34188));
    InMux I__8352 (
            .O(N__34205),
            .I(N__34188));
    InMux I__8351 (
            .O(N__34204),
            .I(N__34188));
    LocalMux I__8350 (
            .O(N__34201),
            .I(N__34183));
    Span4Mux_h I__8349 (
            .O(N__34198),
            .I(N__34180));
    InMux I__8348 (
            .O(N__34197),
            .I(N__34177));
    LocalMux I__8347 (
            .O(N__34188),
            .I(N__34174));
    CascadeMux I__8346 (
            .O(N__34187),
            .I(N__34168));
    InMux I__8345 (
            .O(N__34186),
            .I(N__34165));
    Span4Mux_h I__8344 (
            .O(N__34183),
            .I(N__34162));
    Span4Mux_h I__8343 (
            .O(N__34180),
            .I(N__34155));
    LocalMux I__8342 (
            .O(N__34177),
            .I(N__34155));
    Span4Mux_h I__8341 (
            .O(N__34174),
            .I(N__34155));
    InMux I__8340 (
            .O(N__34173),
            .I(N__34148));
    InMux I__8339 (
            .O(N__34172),
            .I(N__34148));
    InMux I__8338 (
            .O(N__34171),
            .I(N__34148));
    InMux I__8337 (
            .O(N__34168),
            .I(N__34145));
    LocalMux I__8336 (
            .O(N__34165),
            .I(\c0.byte_transmit_counter_3 ));
    Odrv4 I__8335 (
            .O(N__34162),
            .I(\c0.byte_transmit_counter_3 ));
    Odrv4 I__8334 (
            .O(N__34155),
            .I(\c0.byte_transmit_counter_3 ));
    LocalMux I__8333 (
            .O(N__34148),
            .I(\c0.byte_transmit_counter_3 ));
    LocalMux I__8332 (
            .O(N__34145),
            .I(\c0.byte_transmit_counter_3 ));
    InMux I__8331 (
            .O(N__34134),
            .I(N__34123));
    InMux I__8330 (
            .O(N__34133),
            .I(N__34123));
    InMux I__8329 (
            .O(N__34132),
            .I(N__34123));
    InMux I__8328 (
            .O(N__34131),
            .I(N__34118));
    InMux I__8327 (
            .O(N__34130),
            .I(N__34118));
    LocalMux I__8326 (
            .O(N__34123),
            .I(N__34109));
    LocalMux I__8325 (
            .O(N__34118),
            .I(N__34109));
    InMux I__8324 (
            .O(N__34117),
            .I(N__34105));
    InMux I__8323 (
            .O(N__34116),
            .I(N__34098));
    InMux I__8322 (
            .O(N__34115),
            .I(N__34098));
    InMux I__8321 (
            .O(N__34114),
            .I(N__34098));
    Span4Mux_h I__8320 (
            .O(N__34109),
            .I(N__34095));
    InMux I__8319 (
            .O(N__34108),
            .I(N__34092));
    LocalMux I__8318 (
            .O(N__34105),
            .I(\c0.byte_transmit_counter_2 ));
    LocalMux I__8317 (
            .O(N__34098),
            .I(\c0.byte_transmit_counter_2 ));
    Odrv4 I__8316 (
            .O(N__34095),
            .I(\c0.byte_transmit_counter_2 ));
    LocalMux I__8315 (
            .O(N__34092),
            .I(\c0.byte_transmit_counter_2 ));
    CascadeMux I__8314 (
            .O(N__34083),
            .I(\c0.n9_adj_1891_cascade_ ));
    InMux I__8313 (
            .O(N__34080),
            .I(N__34076));
    InMux I__8312 (
            .O(N__34079),
            .I(N__34073));
    LocalMux I__8311 (
            .O(N__34076),
            .I(N__34061));
    LocalMux I__8310 (
            .O(N__34073),
            .I(N__34061));
    InMux I__8309 (
            .O(N__34072),
            .I(N__34050));
    InMux I__8308 (
            .O(N__34071),
            .I(N__34050));
    InMux I__8307 (
            .O(N__34070),
            .I(N__34050));
    InMux I__8306 (
            .O(N__34069),
            .I(N__34043));
    InMux I__8305 (
            .O(N__34068),
            .I(N__34043));
    InMux I__8304 (
            .O(N__34067),
            .I(N__34043));
    InMux I__8303 (
            .O(N__34066),
            .I(N__34040));
    Span4Mux_v I__8302 (
            .O(N__34061),
            .I(N__34037));
    InMux I__8301 (
            .O(N__34060),
            .I(N__34031));
    InMux I__8300 (
            .O(N__34059),
            .I(N__34031));
    InMux I__8299 (
            .O(N__34058),
            .I(N__34026));
    InMux I__8298 (
            .O(N__34057),
            .I(N__34026));
    LocalMux I__8297 (
            .O(N__34050),
            .I(N__34023));
    LocalMux I__8296 (
            .O(N__34043),
            .I(N__34018));
    LocalMux I__8295 (
            .O(N__34040),
            .I(N__34018));
    Span4Mux_h I__8294 (
            .O(N__34037),
            .I(N__34014));
    InMux I__8293 (
            .O(N__34036),
            .I(N__34011));
    LocalMux I__8292 (
            .O(N__34031),
            .I(N__34008));
    LocalMux I__8291 (
            .O(N__34026),
            .I(N__34003));
    Span4Mux_h I__8290 (
            .O(N__34023),
            .I(N__34003));
    Span4Mux_v I__8289 (
            .O(N__34018),
            .I(N__34000));
    InMux I__8288 (
            .O(N__34017),
            .I(N__33997));
    Odrv4 I__8287 (
            .O(N__34014),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__8286 (
            .O(N__34011),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv12 I__8285 (
            .O(N__34008),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__8284 (
            .O(N__34003),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__8283 (
            .O(N__34000),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__8282 (
            .O(N__33997),
            .I(\c0.byte_transmit_counter_1 ));
    InMux I__8281 (
            .O(N__33984),
            .I(N__33981));
    LocalMux I__8280 (
            .O(N__33981),
            .I(N__33978));
    Span4Mux_v I__8279 (
            .O(N__33978),
            .I(N__33975));
    Odrv4 I__8278 (
            .O(N__33975),
            .I(\c0.n15_adj_1893 ));
    InMux I__8277 (
            .O(N__33972),
            .I(N__33968));
    InMux I__8276 (
            .O(N__33971),
            .I(N__33964));
    LocalMux I__8275 (
            .O(N__33968),
            .I(N__33961));
    InMux I__8274 (
            .O(N__33967),
            .I(N__33958));
    LocalMux I__8273 (
            .O(N__33964),
            .I(n5421));
    Odrv4 I__8272 (
            .O(N__33961),
            .I(n5421));
    LocalMux I__8271 (
            .O(N__33958),
            .I(n5421));
    InMux I__8270 (
            .O(N__33951),
            .I(N__33947));
    InMux I__8269 (
            .O(N__33950),
            .I(N__33944));
    LocalMux I__8268 (
            .O(N__33947),
            .I(N__33941));
    LocalMux I__8267 (
            .O(N__33944),
            .I(data_out_18_1));
    Odrv4 I__8266 (
            .O(N__33941),
            .I(data_out_18_1));
    CascadeMux I__8265 (
            .O(N__33936),
            .I(N__33933));
    InMux I__8264 (
            .O(N__33933),
            .I(N__33930));
    LocalMux I__8263 (
            .O(N__33930),
            .I(N__33927));
    Span4Mux_h I__8262 (
            .O(N__33927),
            .I(N__33923));
    InMux I__8261 (
            .O(N__33926),
            .I(N__33920));
    Sp12to4 I__8260 (
            .O(N__33923),
            .I(N__33917));
    LocalMux I__8259 (
            .O(N__33920),
            .I(data_out_19_3));
    Odrv12 I__8258 (
            .O(N__33917),
            .I(data_out_19_3));
    InMux I__8257 (
            .O(N__33912),
            .I(N__33909));
    LocalMux I__8256 (
            .O(N__33909),
            .I(\c0.n5837 ));
    InMux I__8255 (
            .O(N__33906),
            .I(N__33902));
    InMux I__8254 (
            .O(N__33905),
            .I(N__33899));
    LocalMux I__8253 (
            .O(N__33902),
            .I(r_Tx_Data_5));
    LocalMux I__8252 (
            .O(N__33899),
            .I(r_Tx_Data_5));
    CascadeMux I__8251 (
            .O(N__33894),
            .I(N__33889));
    CascadeMux I__8250 (
            .O(N__33893),
            .I(N__33885));
    InMux I__8249 (
            .O(N__33892),
            .I(N__33878));
    InMux I__8248 (
            .O(N__33889),
            .I(N__33878));
    InMux I__8247 (
            .O(N__33888),
            .I(N__33873));
    InMux I__8246 (
            .O(N__33885),
            .I(N__33873));
    CascadeMux I__8245 (
            .O(N__33884),
            .I(N__33870));
    InMux I__8244 (
            .O(N__33883),
            .I(N__33865));
    LocalMux I__8243 (
            .O(N__33878),
            .I(N__33862));
    LocalMux I__8242 (
            .O(N__33873),
            .I(N__33859));
    InMux I__8241 (
            .O(N__33870),
            .I(N__33854));
    InMux I__8240 (
            .O(N__33869),
            .I(N__33854));
    InMux I__8239 (
            .O(N__33868),
            .I(N__33851));
    LocalMux I__8238 (
            .O(N__33865),
            .I(N__33848));
    Span4Mux_h I__8237 (
            .O(N__33862),
            .I(N__33843));
    Span4Mux_v I__8236 (
            .O(N__33859),
            .I(N__33843));
    LocalMux I__8235 (
            .O(N__33854),
            .I(\c0.tx.r_Bit_Index_1 ));
    LocalMux I__8234 (
            .O(N__33851),
            .I(\c0.tx.r_Bit_Index_1 ));
    Odrv12 I__8233 (
            .O(N__33848),
            .I(\c0.tx.r_Bit_Index_1 ));
    Odrv4 I__8232 (
            .O(N__33843),
            .I(\c0.tx.r_Bit_Index_1 ));
    CascadeMux I__8231 (
            .O(N__33834),
            .I(N__33830));
    InMux I__8230 (
            .O(N__33833),
            .I(N__33827));
    InMux I__8229 (
            .O(N__33830),
            .I(N__33824));
    LocalMux I__8228 (
            .O(N__33827),
            .I(N__33819));
    LocalMux I__8227 (
            .O(N__33824),
            .I(N__33819));
    Odrv4 I__8226 (
            .O(N__33819),
            .I(r_Tx_Data_4));
    InMux I__8225 (
            .O(N__33816),
            .I(N__33813));
    LocalMux I__8224 (
            .O(N__33813),
            .I(N__33810));
    Span4Mux_h I__8223 (
            .O(N__33810),
            .I(N__33807));
    Odrv4 I__8222 (
            .O(N__33807),
            .I(\c0.tx.n6285 ));
    InMux I__8221 (
            .O(N__33804),
            .I(N__33801));
    LocalMux I__8220 (
            .O(N__33801),
            .I(\c0.tx.n6288 ));
    CascadeMux I__8219 (
            .O(N__33798),
            .I(N__33795));
    InMux I__8218 (
            .O(N__33795),
            .I(N__33792));
    LocalMux I__8217 (
            .O(N__33792),
            .I(N__33789));
    Span4Mux_h I__8216 (
            .O(N__33789),
            .I(N__33786));
    Odrv4 I__8215 (
            .O(N__33786),
            .I(n5415));
    InMux I__8214 (
            .O(N__33783),
            .I(N__33777));
    CascadeMux I__8213 (
            .O(N__33782),
            .I(N__33774));
    InMux I__8212 (
            .O(N__33781),
            .I(N__33769));
    InMux I__8211 (
            .O(N__33780),
            .I(N__33769));
    LocalMux I__8210 (
            .O(N__33777),
            .I(N__33766));
    InMux I__8209 (
            .O(N__33774),
            .I(N__33763));
    LocalMux I__8208 (
            .O(N__33769),
            .I(N__33760));
    Odrv12 I__8207 (
            .O(N__33766),
            .I(\c0.n1251 ));
    LocalMux I__8206 (
            .O(N__33763),
            .I(\c0.n1251 ));
    Odrv4 I__8205 (
            .O(N__33760),
            .I(\c0.n1251 ));
    CascadeMux I__8204 (
            .O(N__33753),
            .I(N__33750));
    InMux I__8203 (
            .O(N__33750),
            .I(N__33747));
    LocalMux I__8202 (
            .O(N__33747),
            .I(\c0.n5845 ));
    InMux I__8201 (
            .O(N__33744),
            .I(N__33741));
    LocalMux I__8200 (
            .O(N__33741),
            .I(N__33733));
    InMux I__8199 (
            .O(N__33740),
            .I(N__33724));
    InMux I__8198 (
            .O(N__33739),
            .I(N__33724));
    InMux I__8197 (
            .O(N__33738),
            .I(N__33724));
    InMux I__8196 (
            .O(N__33737),
            .I(N__33724));
    InMux I__8195 (
            .O(N__33736),
            .I(N__33719));
    Span4Mux_h I__8194 (
            .O(N__33733),
            .I(N__33714));
    LocalMux I__8193 (
            .O(N__33724),
            .I(N__33714));
    InMux I__8192 (
            .O(N__33723),
            .I(N__33710));
    InMux I__8191 (
            .O(N__33722),
            .I(N__33707));
    LocalMux I__8190 (
            .O(N__33719),
            .I(N__33704));
    Span4Mux_v I__8189 (
            .O(N__33714),
            .I(N__33701));
    InMux I__8188 (
            .O(N__33713),
            .I(N__33698));
    LocalMux I__8187 (
            .O(N__33710),
            .I(\c0.byte_transmit_counter_4 ));
    LocalMux I__8186 (
            .O(N__33707),
            .I(\c0.byte_transmit_counter_4 ));
    Odrv4 I__8185 (
            .O(N__33704),
            .I(\c0.byte_transmit_counter_4 ));
    Odrv4 I__8184 (
            .O(N__33701),
            .I(\c0.byte_transmit_counter_4 ));
    LocalMux I__8183 (
            .O(N__33698),
            .I(\c0.byte_transmit_counter_4 ));
    InMux I__8182 (
            .O(N__33687),
            .I(N__33684));
    LocalMux I__8181 (
            .O(N__33684),
            .I(tx_data_1_N_keep));
    CascadeMux I__8180 (
            .O(N__33681),
            .I(\c0.n9_adj_1906_cascade_ ));
    InMux I__8179 (
            .O(N__33678),
            .I(N__33675));
    LocalMux I__8178 (
            .O(N__33675),
            .I(N__33672));
    Odrv4 I__8177 (
            .O(N__33672),
            .I(\c0.n15_adj_1909 ));
    InMux I__8176 (
            .O(N__33669),
            .I(N__33666));
    LocalMux I__8175 (
            .O(N__33666),
            .I(N__33661));
    InMux I__8174 (
            .O(N__33665),
            .I(N__33658));
    InMux I__8173 (
            .O(N__33664),
            .I(N__33652));
    Span12Mux_v I__8172 (
            .O(N__33661),
            .I(N__33647));
    LocalMux I__8171 (
            .O(N__33658),
            .I(N__33647));
    InMux I__8170 (
            .O(N__33657),
            .I(N__33640));
    InMux I__8169 (
            .O(N__33656),
            .I(N__33640));
    InMux I__8168 (
            .O(N__33655),
            .I(N__33640));
    LocalMux I__8167 (
            .O(N__33652),
            .I(data_out_10_4));
    Odrv12 I__8166 (
            .O(N__33647),
            .I(data_out_10_4));
    LocalMux I__8165 (
            .O(N__33640),
            .I(data_out_10_4));
    InMux I__8164 (
            .O(N__33633),
            .I(N__33630));
    LocalMux I__8163 (
            .O(N__33630),
            .I(N__33627));
    Odrv12 I__8162 (
            .O(N__33627),
            .I(\c0.n2293 ));
    InMux I__8161 (
            .O(N__33624),
            .I(N__33621));
    LocalMux I__8160 (
            .O(N__33621),
            .I(N__33618));
    Span4Mux_v I__8159 (
            .O(N__33618),
            .I(N__33615));
    Odrv4 I__8158 (
            .O(N__33615),
            .I(n4_adj_1996));
    CascadeMux I__8157 (
            .O(N__33612),
            .I(N__33606));
    InMux I__8156 (
            .O(N__33611),
            .I(N__33602));
    InMux I__8155 (
            .O(N__33610),
            .I(N__33599));
    InMux I__8154 (
            .O(N__33609),
            .I(N__33595));
    InMux I__8153 (
            .O(N__33606),
            .I(N__33592));
    InMux I__8152 (
            .O(N__33605),
            .I(N__33589));
    LocalMux I__8151 (
            .O(N__33602),
            .I(N__33586));
    LocalMux I__8150 (
            .O(N__33599),
            .I(N__33583));
    InMux I__8149 (
            .O(N__33598),
            .I(N__33580));
    LocalMux I__8148 (
            .O(N__33595),
            .I(N__33577));
    LocalMux I__8147 (
            .O(N__33592),
            .I(N__33572));
    LocalMux I__8146 (
            .O(N__33589),
            .I(N__33572));
    Span4Mux_v I__8145 (
            .O(N__33586),
            .I(N__33563));
    Span4Mux_v I__8144 (
            .O(N__33583),
            .I(N__33563));
    LocalMux I__8143 (
            .O(N__33580),
            .I(N__33563));
    Span4Mux_v I__8142 (
            .O(N__33577),
            .I(N__33558));
    Span4Mux_v I__8141 (
            .O(N__33572),
            .I(N__33558));
    InMux I__8140 (
            .O(N__33571),
            .I(N__33555));
    InMux I__8139 (
            .O(N__33570),
            .I(N__33552));
    Span4Mux_h I__8138 (
            .O(N__33563),
            .I(N__33549));
    Sp12to4 I__8137 (
            .O(N__33558),
            .I(N__33544));
    LocalMux I__8136 (
            .O(N__33555),
            .I(N__33544));
    LocalMux I__8135 (
            .O(N__33552),
            .I(N__33541));
    Odrv4 I__8134 (
            .O(N__33549),
            .I(n1519));
    Odrv12 I__8133 (
            .O(N__33544),
            .I(n1519));
    Odrv4 I__8132 (
            .O(N__33541),
            .I(n1519));
    InMux I__8131 (
            .O(N__33534),
            .I(N__33531));
    LocalMux I__8130 (
            .O(N__33531),
            .I(tx_data_5_N_keep));
    CascadeMux I__8129 (
            .O(N__33528),
            .I(\c0.n95_cascade_ ));
    InMux I__8128 (
            .O(N__33525),
            .I(N__33519));
    InMux I__8127 (
            .O(N__33524),
            .I(N__33519));
    LocalMux I__8126 (
            .O(N__33519),
            .I(\c0.n106 ));
    CascadeMux I__8125 (
            .O(N__33516),
            .I(N__33513));
    InMux I__8124 (
            .O(N__33513),
            .I(N__33510));
    LocalMux I__8123 (
            .O(N__33510),
            .I(N__33507));
    Odrv12 I__8122 (
            .O(N__33507),
            .I(n4_adj_1981));
    CascadeMux I__8121 (
            .O(N__33504),
            .I(N__33501));
    InMux I__8120 (
            .O(N__33501),
            .I(N__33498));
    LocalMux I__8119 (
            .O(N__33498),
            .I(N__33495));
    Odrv4 I__8118 (
            .O(N__33495),
            .I(n7_adj_1988));
    InMux I__8117 (
            .O(N__33492),
            .I(N__33483));
    InMux I__8116 (
            .O(N__33491),
            .I(N__33483));
    InMux I__8115 (
            .O(N__33490),
            .I(N__33476));
    InMux I__8114 (
            .O(N__33489),
            .I(N__33476));
    InMux I__8113 (
            .O(N__33488),
            .I(N__33476));
    LocalMux I__8112 (
            .O(N__33483),
            .I(\c0.n15 ));
    LocalMux I__8111 (
            .O(N__33476),
            .I(\c0.n15 ));
    CascadeMux I__8110 (
            .O(N__33471),
            .I(N__33468));
    InMux I__8109 (
            .O(N__33468),
            .I(N__33461));
    InMux I__8108 (
            .O(N__33467),
            .I(N__33461));
    InMux I__8107 (
            .O(N__33466),
            .I(N__33458));
    LocalMux I__8106 (
            .O(N__33461),
            .I(N__33451));
    LocalMux I__8105 (
            .O(N__33458),
            .I(N__33451));
    InMux I__8104 (
            .O(N__33457),
            .I(N__33448));
    InMux I__8103 (
            .O(N__33456),
            .I(N__33445));
    Odrv4 I__8102 (
            .O(N__33451),
            .I(\c0.n81_adj_1872 ));
    LocalMux I__8101 (
            .O(N__33448),
            .I(\c0.n81_adj_1872 ));
    LocalMux I__8100 (
            .O(N__33445),
            .I(\c0.n81_adj_1872 ));
    CascadeMux I__8099 (
            .O(N__33438),
            .I(N__33433));
    InMux I__8098 (
            .O(N__33437),
            .I(N__33429));
    InMux I__8097 (
            .O(N__33436),
            .I(N__33422));
    InMux I__8096 (
            .O(N__33433),
            .I(N__33422));
    InMux I__8095 (
            .O(N__33432),
            .I(N__33422));
    LocalMux I__8094 (
            .O(N__33429),
            .I(\c0.tx_transmit_N_568_4 ));
    LocalMux I__8093 (
            .O(N__33422),
            .I(\c0.tx_transmit_N_568_4 ));
    InMux I__8092 (
            .O(N__33417),
            .I(N__33411));
    InMux I__8091 (
            .O(N__33416),
            .I(N__33411));
    LocalMux I__8090 (
            .O(N__33411),
            .I(\c0.tx_transmit_N_568_2 ));
    CascadeMux I__8089 (
            .O(N__33408),
            .I(N__33405));
    InMux I__8088 (
            .O(N__33405),
            .I(N__33402));
    LocalMux I__8087 (
            .O(N__33402),
            .I(N__33399));
    Odrv12 I__8086 (
            .O(N__33399),
            .I(\c0.n5833 ));
    CascadeMux I__8085 (
            .O(N__33396),
            .I(N__33393));
    InMux I__8084 (
            .O(N__33393),
            .I(N__33390));
    LocalMux I__8083 (
            .O(N__33390),
            .I(N__33387));
    Span4Mux_h I__8082 (
            .O(N__33387),
            .I(N__33384));
    Odrv4 I__8081 (
            .O(N__33384),
            .I(\c0.n31_adj_1912 ));
    InMux I__8080 (
            .O(N__33381),
            .I(N__33378));
    LocalMux I__8079 (
            .O(N__33378),
            .I(\c0.n989 ));
    InMux I__8078 (
            .O(N__33375),
            .I(\c0.n4703 ));
    InMux I__8077 (
            .O(N__33372),
            .I(\c0.n4704 ));
    InMux I__8076 (
            .O(N__33369),
            .I(\c0.n4705 ));
    InMux I__8075 (
            .O(N__33366),
            .I(\c0.n4706 ));
    InMux I__8074 (
            .O(N__33363),
            .I(N__33360));
    LocalMux I__8073 (
            .O(N__33360),
            .I(\c0.byte_transmit_counter_5 ));
    InMux I__8072 (
            .O(N__33357),
            .I(N__33351));
    InMux I__8071 (
            .O(N__33356),
            .I(N__33351));
    LocalMux I__8070 (
            .O(N__33351),
            .I(\c0.tx_transmit_N_568_5 ));
    InMux I__8069 (
            .O(N__33348),
            .I(\c0.n4707 ));
    InMux I__8068 (
            .O(N__33345),
            .I(N__33342));
    LocalMux I__8067 (
            .O(N__33342),
            .I(N__33339));
    Odrv4 I__8066 (
            .O(N__33339),
            .I(\c0.byte_transmit_counter_6 ));
    InMux I__8065 (
            .O(N__33336),
            .I(N__33333));
    LocalMux I__8064 (
            .O(N__33333),
            .I(N__33329));
    InMux I__8063 (
            .O(N__33332),
            .I(N__33326));
    Odrv4 I__8062 (
            .O(N__33329),
            .I(\c0.tx_transmit_N_568_6 ));
    LocalMux I__8061 (
            .O(N__33326),
            .I(\c0.tx_transmit_N_568_6 ));
    InMux I__8060 (
            .O(N__33321),
            .I(\c0.n4708 ));
    InMux I__8059 (
            .O(N__33318),
            .I(N__33315));
    LocalMux I__8058 (
            .O(N__33315),
            .I(N__33312));
    Odrv4 I__8057 (
            .O(N__33312),
            .I(\c0.byte_transmit_counter_7 ));
    InMux I__8056 (
            .O(N__33309),
            .I(\c0.n4709 ));
    InMux I__8055 (
            .O(N__33306),
            .I(N__33303));
    LocalMux I__8054 (
            .O(N__33303),
            .I(N__33299));
    InMux I__8053 (
            .O(N__33302),
            .I(N__33296));
    Odrv4 I__8052 (
            .O(N__33299),
            .I(\c0.tx_transmit_N_568_7 ));
    LocalMux I__8051 (
            .O(N__33296),
            .I(\c0.tx_transmit_N_568_7 ));
    InMux I__8050 (
            .O(N__33291),
            .I(N__33285));
    InMux I__8049 (
            .O(N__33290),
            .I(N__33285));
    LocalMux I__8048 (
            .O(N__33285),
            .I(\c0.tx_transmit_N_568_3 ));
    InMux I__8047 (
            .O(N__33282),
            .I(N__33279));
    LocalMux I__8046 (
            .O(N__33279),
            .I(\c0.n95 ));
    CascadeMux I__8045 (
            .O(N__33276),
            .I(N__33264));
    CascadeMux I__8044 (
            .O(N__33275),
            .I(N__33258));
    CascadeMux I__8043 (
            .O(N__33274),
            .I(N__33255));
    CascadeMux I__8042 (
            .O(N__33273),
            .I(N__33247));
    CascadeMux I__8041 (
            .O(N__33272),
            .I(N__33235));
    InMux I__8040 (
            .O(N__33271),
            .I(N__33220));
    InMux I__8039 (
            .O(N__33270),
            .I(N__33220));
    InMux I__8038 (
            .O(N__33269),
            .I(N__33220));
    InMux I__8037 (
            .O(N__33268),
            .I(N__33212));
    InMux I__8036 (
            .O(N__33267),
            .I(N__33212));
    InMux I__8035 (
            .O(N__33264),
            .I(N__33203));
    InMux I__8034 (
            .O(N__33263),
            .I(N__33203));
    InMux I__8033 (
            .O(N__33262),
            .I(N__33203));
    InMux I__8032 (
            .O(N__33261),
            .I(N__33203));
    InMux I__8031 (
            .O(N__33258),
            .I(N__33198));
    InMux I__8030 (
            .O(N__33255),
            .I(N__33198));
    InMux I__8029 (
            .O(N__33254),
            .I(N__33191));
    InMux I__8028 (
            .O(N__33253),
            .I(N__33191));
    InMux I__8027 (
            .O(N__33252),
            .I(N__33191));
    InMux I__8026 (
            .O(N__33251),
            .I(N__33186));
    InMux I__8025 (
            .O(N__33250),
            .I(N__33186));
    InMux I__8024 (
            .O(N__33247),
            .I(N__33183));
    InMux I__8023 (
            .O(N__33246),
            .I(N__33180));
    CascadeMux I__8022 (
            .O(N__33245),
            .I(N__33177));
    CascadeMux I__8021 (
            .O(N__33244),
            .I(N__33170));
    CascadeMux I__8020 (
            .O(N__33243),
            .I(N__33167));
    CascadeMux I__8019 (
            .O(N__33242),
            .I(N__33160));
    InMux I__8018 (
            .O(N__33241),
            .I(N__33144));
    InMux I__8017 (
            .O(N__33240),
            .I(N__33144));
    InMux I__8016 (
            .O(N__33239),
            .I(N__33144));
    InMux I__8015 (
            .O(N__33238),
            .I(N__33144));
    InMux I__8014 (
            .O(N__33235),
            .I(N__33139));
    InMux I__8013 (
            .O(N__33234),
            .I(N__33139));
    CascadeMux I__8012 (
            .O(N__33233),
            .I(N__33132));
    CascadeMux I__8011 (
            .O(N__33232),
            .I(N__33126));
    InMux I__8010 (
            .O(N__33231),
            .I(N__33112));
    InMux I__8009 (
            .O(N__33230),
            .I(N__33112));
    CascadeMux I__8008 (
            .O(N__33229),
            .I(N__33109));
    CascadeMux I__8007 (
            .O(N__33228),
            .I(N__33099));
    InMux I__8006 (
            .O(N__33227),
            .I(N__33091));
    LocalMux I__8005 (
            .O(N__33220),
            .I(N__33088));
    CascadeMux I__8004 (
            .O(N__33219),
            .I(N__33078));
    CascadeMux I__8003 (
            .O(N__33218),
            .I(N__33071));
    CascadeMux I__8002 (
            .O(N__33217),
            .I(N__33065));
    LocalMux I__8001 (
            .O(N__33212),
            .I(N__33062));
    LocalMux I__8000 (
            .O(N__33203),
            .I(N__33055));
    LocalMux I__7999 (
            .O(N__33198),
            .I(N__33055));
    LocalMux I__7998 (
            .O(N__33191),
            .I(N__33055));
    LocalMux I__7997 (
            .O(N__33186),
            .I(N__33050));
    LocalMux I__7996 (
            .O(N__33183),
            .I(N__33050));
    LocalMux I__7995 (
            .O(N__33180),
            .I(N__33047));
    InMux I__7994 (
            .O(N__33177),
            .I(N__33038));
    InMux I__7993 (
            .O(N__33176),
            .I(N__33038));
    InMux I__7992 (
            .O(N__33175),
            .I(N__33038));
    InMux I__7991 (
            .O(N__33174),
            .I(N__33038));
    InMux I__7990 (
            .O(N__33173),
            .I(N__33027));
    InMux I__7989 (
            .O(N__33170),
            .I(N__33027));
    InMux I__7988 (
            .O(N__33167),
            .I(N__33027));
    InMux I__7987 (
            .O(N__33166),
            .I(N__33027));
    InMux I__7986 (
            .O(N__33165),
            .I(N__33027));
    InMux I__7985 (
            .O(N__33164),
            .I(N__33015));
    InMux I__7984 (
            .O(N__33163),
            .I(N__33015));
    InMux I__7983 (
            .O(N__33160),
            .I(N__33015));
    InMux I__7982 (
            .O(N__33159),
            .I(N__33015));
    InMux I__7981 (
            .O(N__33158),
            .I(N__33015));
    InMux I__7980 (
            .O(N__33157),
            .I(N__33010));
    InMux I__7979 (
            .O(N__33156),
            .I(N__33010));
    CascadeMux I__7978 (
            .O(N__33155),
            .I(N__33007));
    InMux I__7977 (
            .O(N__33154),
            .I(N__33000));
    InMux I__7976 (
            .O(N__33153),
            .I(N__33000));
    LocalMux I__7975 (
            .O(N__33144),
            .I(N__32995));
    LocalMux I__7974 (
            .O(N__33139),
            .I(N__32995));
    InMux I__7973 (
            .O(N__33138),
            .I(N__32979));
    CascadeMux I__7972 (
            .O(N__33137),
            .I(N__32974));
    CascadeMux I__7971 (
            .O(N__33136),
            .I(N__32971));
    InMux I__7970 (
            .O(N__33135),
            .I(N__32958));
    InMux I__7969 (
            .O(N__33132),
            .I(N__32958));
    InMux I__7968 (
            .O(N__33131),
            .I(N__32958));
    InMux I__7967 (
            .O(N__33130),
            .I(N__32958));
    InMux I__7966 (
            .O(N__33129),
            .I(N__32958));
    InMux I__7965 (
            .O(N__33126),
            .I(N__32953));
    InMux I__7964 (
            .O(N__33125),
            .I(N__32953));
    InMux I__7963 (
            .O(N__33124),
            .I(N__32944));
    InMux I__7962 (
            .O(N__33123),
            .I(N__32944));
    InMux I__7961 (
            .O(N__33122),
            .I(N__32944));
    InMux I__7960 (
            .O(N__33121),
            .I(N__32944));
    InMux I__7959 (
            .O(N__33120),
            .I(N__32935));
    InMux I__7958 (
            .O(N__33119),
            .I(N__32935));
    InMux I__7957 (
            .O(N__33118),
            .I(N__32935));
    InMux I__7956 (
            .O(N__33117),
            .I(N__32935));
    LocalMux I__7955 (
            .O(N__33112),
            .I(N__32932));
    InMux I__7954 (
            .O(N__33109),
            .I(N__32925));
    InMux I__7953 (
            .O(N__33108),
            .I(N__32925));
    InMux I__7952 (
            .O(N__33107),
            .I(N__32925));
    InMux I__7951 (
            .O(N__33106),
            .I(N__32920));
    InMux I__7950 (
            .O(N__33105),
            .I(N__32920));
    InMux I__7949 (
            .O(N__33104),
            .I(N__32917));
    InMux I__7948 (
            .O(N__33103),
            .I(N__32913));
    InMux I__7947 (
            .O(N__33102),
            .I(N__32910));
    InMux I__7946 (
            .O(N__33099),
            .I(N__32905));
    InMux I__7945 (
            .O(N__33098),
            .I(N__32905));
    InMux I__7944 (
            .O(N__33097),
            .I(N__32896));
    InMux I__7943 (
            .O(N__33096),
            .I(N__32896));
    InMux I__7942 (
            .O(N__33095),
            .I(N__32896));
    InMux I__7941 (
            .O(N__33094),
            .I(N__32896));
    LocalMux I__7940 (
            .O(N__33091),
            .I(N__32891));
    Span4Mux_v I__7939 (
            .O(N__33088),
            .I(N__32888));
    InMux I__7938 (
            .O(N__33087),
            .I(N__32881));
    InMux I__7937 (
            .O(N__33086),
            .I(N__32881));
    InMux I__7936 (
            .O(N__33085),
            .I(N__32881));
    InMux I__7935 (
            .O(N__33084),
            .I(N__32878));
    InMux I__7934 (
            .O(N__33083),
            .I(N__32875));
    InMux I__7933 (
            .O(N__33082),
            .I(N__32870));
    InMux I__7932 (
            .O(N__33081),
            .I(N__32870));
    InMux I__7931 (
            .O(N__33078),
            .I(N__32865));
    InMux I__7930 (
            .O(N__33077),
            .I(N__32862));
    InMux I__7929 (
            .O(N__33076),
            .I(N__32853));
    InMux I__7928 (
            .O(N__33075),
            .I(N__32853));
    InMux I__7927 (
            .O(N__33074),
            .I(N__32853));
    InMux I__7926 (
            .O(N__33071),
            .I(N__32848));
    InMux I__7925 (
            .O(N__33070),
            .I(N__32848));
    CascadeMux I__7924 (
            .O(N__33069),
            .I(N__32843));
    CascadeMux I__7923 (
            .O(N__33068),
            .I(N__32840));
    InMux I__7922 (
            .O(N__33065),
            .I(N__32835));
    Span4Mux_v I__7921 (
            .O(N__33062),
            .I(N__32824));
    Span4Mux_v I__7920 (
            .O(N__33055),
            .I(N__32824));
    Span4Mux_v I__7919 (
            .O(N__33050),
            .I(N__32824));
    Span4Mux_v I__7918 (
            .O(N__33047),
            .I(N__32824));
    LocalMux I__7917 (
            .O(N__33038),
            .I(N__32824));
    LocalMux I__7916 (
            .O(N__33027),
            .I(N__32821));
    InMux I__7915 (
            .O(N__33026),
            .I(N__32818));
    LocalMux I__7914 (
            .O(N__33015),
            .I(N__32813));
    LocalMux I__7913 (
            .O(N__33010),
            .I(N__32813));
    InMux I__7912 (
            .O(N__33007),
            .I(N__32808));
    InMux I__7911 (
            .O(N__33006),
            .I(N__32808));
    InMux I__7910 (
            .O(N__33005),
            .I(N__32801));
    LocalMux I__7909 (
            .O(N__33000),
            .I(N__32798));
    Span4Mux_h I__7908 (
            .O(N__32995),
            .I(N__32795));
    InMux I__7907 (
            .O(N__32994),
            .I(N__32784));
    InMux I__7906 (
            .O(N__32993),
            .I(N__32784));
    InMux I__7905 (
            .O(N__32992),
            .I(N__32784));
    InMux I__7904 (
            .O(N__32991),
            .I(N__32784));
    InMux I__7903 (
            .O(N__32990),
            .I(N__32784));
    InMux I__7902 (
            .O(N__32989),
            .I(N__32781));
    CascadeMux I__7901 (
            .O(N__32988),
            .I(N__32774));
    CascadeMux I__7900 (
            .O(N__32987),
            .I(N__32770));
    CascadeMux I__7899 (
            .O(N__32986),
            .I(N__32764));
    InMux I__7898 (
            .O(N__32985),
            .I(N__32747));
    InMux I__7897 (
            .O(N__32984),
            .I(N__32747));
    InMux I__7896 (
            .O(N__32983),
            .I(N__32747));
    InMux I__7895 (
            .O(N__32982),
            .I(N__32747));
    LocalMux I__7894 (
            .O(N__32979),
            .I(N__32744));
    InMux I__7893 (
            .O(N__32978),
            .I(N__32739));
    InMux I__7892 (
            .O(N__32977),
            .I(N__32739));
    InMux I__7891 (
            .O(N__32974),
            .I(N__32734));
    InMux I__7890 (
            .O(N__32971),
            .I(N__32734));
    InMux I__7889 (
            .O(N__32970),
            .I(N__32729));
    InMux I__7888 (
            .O(N__32969),
            .I(N__32729));
    LocalMux I__7887 (
            .O(N__32958),
            .I(N__32726));
    LocalMux I__7886 (
            .O(N__32953),
            .I(N__32723));
    LocalMux I__7885 (
            .O(N__32944),
            .I(N__32718));
    LocalMux I__7884 (
            .O(N__32935),
            .I(N__32718));
    Span4Mux_v I__7883 (
            .O(N__32932),
            .I(N__32709));
    LocalMux I__7882 (
            .O(N__32925),
            .I(N__32709));
    LocalMux I__7881 (
            .O(N__32920),
            .I(N__32709));
    LocalMux I__7880 (
            .O(N__32917),
            .I(N__32709));
    CascadeMux I__7879 (
            .O(N__32916),
            .I(N__32706));
    LocalMux I__7878 (
            .O(N__32913),
            .I(N__32695));
    LocalMux I__7877 (
            .O(N__32910),
            .I(N__32695));
    LocalMux I__7876 (
            .O(N__32905),
            .I(N__32695));
    LocalMux I__7875 (
            .O(N__32896),
            .I(N__32695));
    InMux I__7874 (
            .O(N__32895),
            .I(N__32690));
    InMux I__7873 (
            .O(N__32894),
            .I(N__32690));
    Span4Mux_v I__7872 (
            .O(N__32891),
            .I(N__32681));
    Span4Mux_v I__7871 (
            .O(N__32888),
            .I(N__32681));
    LocalMux I__7870 (
            .O(N__32881),
            .I(N__32681));
    LocalMux I__7869 (
            .O(N__32878),
            .I(N__32681));
    LocalMux I__7868 (
            .O(N__32875),
            .I(N__32676));
    LocalMux I__7867 (
            .O(N__32870),
            .I(N__32676));
    InMux I__7866 (
            .O(N__32869),
            .I(N__32671));
    InMux I__7865 (
            .O(N__32868),
            .I(N__32671));
    LocalMux I__7864 (
            .O(N__32865),
            .I(N__32666));
    LocalMux I__7863 (
            .O(N__32862),
            .I(N__32666));
    InMux I__7862 (
            .O(N__32861),
            .I(N__32661));
    InMux I__7861 (
            .O(N__32860),
            .I(N__32661));
    LocalMux I__7860 (
            .O(N__32853),
            .I(N__32656));
    LocalMux I__7859 (
            .O(N__32848),
            .I(N__32656));
    InMux I__7858 (
            .O(N__32847),
            .I(N__32649));
    InMux I__7857 (
            .O(N__32846),
            .I(N__32649));
    InMux I__7856 (
            .O(N__32843),
            .I(N__32649));
    InMux I__7855 (
            .O(N__32840),
            .I(N__32644));
    InMux I__7854 (
            .O(N__32839),
            .I(N__32644));
    CascadeMux I__7853 (
            .O(N__32838),
            .I(N__32640));
    LocalMux I__7852 (
            .O(N__32835),
            .I(N__32632));
    Span4Mux_h I__7851 (
            .O(N__32824),
            .I(N__32632));
    Span4Mux_h I__7850 (
            .O(N__32821),
            .I(N__32623));
    LocalMux I__7849 (
            .O(N__32818),
            .I(N__32623));
    Span4Mux_h I__7848 (
            .O(N__32813),
            .I(N__32623));
    LocalMux I__7847 (
            .O(N__32808),
            .I(N__32623));
    InMux I__7846 (
            .O(N__32807),
            .I(N__32614));
    InMux I__7845 (
            .O(N__32806),
            .I(N__32614));
    InMux I__7844 (
            .O(N__32805),
            .I(N__32614));
    InMux I__7843 (
            .O(N__32804),
            .I(N__32614));
    LocalMux I__7842 (
            .O(N__32801),
            .I(N__32603));
    Span4Mux_v I__7841 (
            .O(N__32798),
            .I(N__32603));
    Span4Mux_h I__7840 (
            .O(N__32795),
            .I(N__32603));
    LocalMux I__7839 (
            .O(N__32784),
            .I(N__32603));
    LocalMux I__7838 (
            .O(N__32781),
            .I(N__32603));
    CascadeMux I__7837 (
            .O(N__32780),
            .I(N__32599));
    CascadeMux I__7836 (
            .O(N__32779),
            .I(N__32595));
    CascadeMux I__7835 (
            .O(N__32778),
            .I(N__32592));
    InMux I__7834 (
            .O(N__32777),
            .I(N__32582));
    InMux I__7833 (
            .O(N__32774),
            .I(N__32582));
    InMux I__7832 (
            .O(N__32773),
            .I(N__32575));
    InMux I__7831 (
            .O(N__32770),
            .I(N__32575));
    InMux I__7830 (
            .O(N__32769),
            .I(N__32575));
    InMux I__7829 (
            .O(N__32768),
            .I(N__32572));
    InMux I__7828 (
            .O(N__32767),
            .I(N__32563));
    InMux I__7827 (
            .O(N__32764),
            .I(N__32563));
    InMux I__7826 (
            .O(N__32763),
            .I(N__32563));
    InMux I__7825 (
            .O(N__32762),
            .I(N__32563));
    InMux I__7824 (
            .O(N__32761),
            .I(N__32554));
    InMux I__7823 (
            .O(N__32760),
            .I(N__32554));
    InMux I__7822 (
            .O(N__32759),
            .I(N__32554));
    InMux I__7821 (
            .O(N__32758),
            .I(N__32554));
    InMux I__7820 (
            .O(N__32757),
            .I(N__32549));
    InMux I__7819 (
            .O(N__32756),
            .I(N__32549));
    LocalMux I__7818 (
            .O(N__32747),
            .I(N__32542));
    Span4Mux_v I__7817 (
            .O(N__32744),
            .I(N__32542));
    LocalMux I__7816 (
            .O(N__32739),
            .I(N__32542));
    LocalMux I__7815 (
            .O(N__32734),
            .I(N__32531));
    LocalMux I__7814 (
            .O(N__32729),
            .I(N__32531));
    Span4Mux_v I__7813 (
            .O(N__32726),
            .I(N__32531));
    Span4Mux_h I__7812 (
            .O(N__32723),
            .I(N__32531));
    Span4Mux_v I__7811 (
            .O(N__32718),
            .I(N__32531));
    Span4Mux_v I__7810 (
            .O(N__32709),
            .I(N__32528));
    InMux I__7809 (
            .O(N__32706),
            .I(N__32521));
    InMux I__7808 (
            .O(N__32705),
            .I(N__32521));
    InMux I__7807 (
            .O(N__32704),
            .I(N__32521));
    Span4Mux_h I__7806 (
            .O(N__32695),
            .I(N__32516));
    LocalMux I__7805 (
            .O(N__32690),
            .I(N__32516));
    Span4Mux_h I__7804 (
            .O(N__32681),
            .I(N__32505));
    Span4Mux_h I__7803 (
            .O(N__32676),
            .I(N__32505));
    LocalMux I__7802 (
            .O(N__32671),
            .I(N__32505));
    Span4Mux_v I__7801 (
            .O(N__32666),
            .I(N__32505));
    LocalMux I__7800 (
            .O(N__32661),
            .I(N__32505));
    Span4Mux_v I__7799 (
            .O(N__32656),
            .I(N__32502));
    LocalMux I__7798 (
            .O(N__32649),
            .I(N__32497));
    LocalMux I__7797 (
            .O(N__32644),
            .I(N__32497));
    InMux I__7796 (
            .O(N__32643),
            .I(N__32494));
    InMux I__7795 (
            .O(N__32640),
            .I(N__32485));
    InMux I__7794 (
            .O(N__32639),
            .I(N__32485));
    InMux I__7793 (
            .O(N__32638),
            .I(N__32485));
    InMux I__7792 (
            .O(N__32637),
            .I(N__32485));
    Span4Mux_s1_h I__7791 (
            .O(N__32632),
            .I(N__32480));
    Span4Mux_h I__7790 (
            .O(N__32623),
            .I(N__32480));
    LocalMux I__7789 (
            .O(N__32614),
            .I(N__32475));
    Span4Mux_h I__7788 (
            .O(N__32603),
            .I(N__32475));
    InMux I__7787 (
            .O(N__32602),
            .I(N__32469));
    InMux I__7786 (
            .O(N__32599),
            .I(N__32469));
    InMux I__7785 (
            .O(N__32598),
            .I(N__32462));
    InMux I__7784 (
            .O(N__32595),
            .I(N__32462));
    InMux I__7783 (
            .O(N__32592),
            .I(N__32462));
    InMux I__7782 (
            .O(N__32591),
            .I(N__32459));
    InMux I__7781 (
            .O(N__32590),
            .I(N__32454));
    InMux I__7780 (
            .O(N__32589),
            .I(N__32454));
    InMux I__7779 (
            .O(N__32588),
            .I(N__32449));
    InMux I__7778 (
            .O(N__32587),
            .I(N__32449));
    LocalMux I__7777 (
            .O(N__32582),
            .I(N__32444));
    LocalMux I__7776 (
            .O(N__32575),
            .I(N__32444));
    LocalMux I__7775 (
            .O(N__32572),
            .I(N__32439));
    LocalMux I__7774 (
            .O(N__32563),
            .I(N__32439));
    LocalMux I__7773 (
            .O(N__32554),
            .I(N__32434));
    LocalMux I__7772 (
            .O(N__32549),
            .I(N__32429));
    Span4Mux_v I__7771 (
            .O(N__32542),
            .I(N__32429));
    Span4Mux_v I__7770 (
            .O(N__32531),
            .I(N__32426));
    Span4Mux_v I__7769 (
            .O(N__32528),
            .I(N__32423));
    LocalMux I__7768 (
            .O(N__32521),
            .I(N__32420));
    Span4Mux_v I__7767 (
            .O(N__32516),
            .I(N__32417));
    Span4Mux_v I__7766 (
            .O(N__32505),
            .I(N__32414));
    Span4Mux_v I__7765 (
            .O(N__32502),
            .I(N__32411));
    Span4Mux_v I__7764 (
            .O(N__32497),
            .I(N__32400));
    LocalMux I__7763 (
            .O(N__32494),
            .I(N__32400));
    LocalMux I__7762 (
            .O(N__32485),
            .I(N__32400));
    Span4Mux_v I__7761 (
            .O(N__32480),
            .I(N__32400));
    Span4Mux_h I__7760 (
            .O(N__32475),
            .I(N__32400));
    InMux I__7759 (
            .O(N__32474),
            .I(N__32397));
    LocalMux I__7758 (
            .O(N__32469),
            .I(N__32394));
    LocalMux I__7757 (
            .O(N__32462),
            .I(N__32391));
    LocalMux I__7756 (
            .O(N__32459),
            .I(N__32380));
    LocalMux I__7755 (
            .O(N__32454),
            .I(N__32380));
    LocalMux I__7754 (
            .O(N__32449),
            .I(N__32380));
    Span4Mux_h I__7753 (
            .O(N__32444),
            .I(N__32380));
    Span4Mux_v I__7752 (
            .O(N__32439),
            .I(N__32380));
    CascadeMux I__7751 (
            .O(N__32438),
            .I(N__32376));
    CascadeMux I__7750 (
            .O(N__32437),
            .I(N__32373));
    Span4Mux_v I__7749 (
            .O(N__32434),
            .I(N__32363));
    Span4Mux_v I__7748 (
            .O(N__32429),
            .I(N__32363));
    Span4Mux_h I__7747 (
            .O(N__32426),
            .I(N__32363));
    Span4Mux_h I__7746 (
            .O(N__32423),
            .I(N__32363));
    Span4Mux_v I__7745 (
            .O(N__32420),
            .I(N__32354));
    Span4Mux_v I__7744 (
            .O(N__32417),
            .I(N__32354));
    Span4Mux_v I__7743 (
            .O(N__32414),
            .I(N__32354));
    Span4Mux_h I__7742 (
            .O(N__32411),
            .I(N__32354));
    Span4Mux_h I__7741 (
            .O(N__32400),
            .I(N__32351));
    LocalMux I__7740 (
            .O(N__32397),
            .I(N__32348));
    Span4Mux_h I__7739 (
            .O(N__32394),
            .I(N__32343));
    Span4Mux_v I__7738 (
            .O(N__32391),
            .I(N__32343));
    Span4Mux_v I__7737 (
            .O(N__32380),
            .I(N__32340));
    InMux I__7736 (
            .O(N__32379),
            .I(N__32333));
    InMux I__7735 (
            .O(N__32376),
            .I(N__32333));
    InMux I__7734 (
            .O(N__32373),
            .I(N__32333));
    InMux I__7733 (
            .O(N__32372),
            .I(N__32330));
    Span4Mux_h I__7732 (
            .O(N__32363),
            .I(N__32327));
    Span4Mux_h I__7731 (
            .O(N__32354),
            .I(N__32324));
    Span4Mux_v I__7730 (
            .O(N__32351),
            .I(N__32321));
    Odrv4 I__7729 (
            .O(N__32348),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__7728 (
            .O(N__32343),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__7727 (
            .O(N__32340),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    LocalMux I__7726 (
            .O(N__32333),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    LocalMux I__7725 (
            .O(N__32330),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__7724 (
            .O(N__32327),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__7723 (
            .O(N__32324),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    Odrv4 I__7722 (
            .O(N__32321),
            .I(\c0.FRAME_MATCHER_wait_for_transmission ));
    InMux I__7721 (
            .O(N__32304),
            .I(N__32300));
    CascadeMux I__7720 (
            .O(N__32303),
            .I(N__32297));
    LocalMux I__7719 (
            .O(N__32300),
            .I(N__32279));
    InMux I__7718 (
            .O(N__32297),
            .I(N__32276));
    InMux I__7717 (
            .O(N__32296),
            .I(N__32273));
    InMux I__7716 (
            .O(N__32295),
            .I(N__32268));
    InMux I__7715 (
            .O(N__32294),
            .I(N__32268));
    InMux I__7714 (
            .O(N__32293),
            .I(N__32265));
    InMux I__7713 (
            .O(N__32292),
            .I(N__32258));
    InMux I__7712 (
            .O(N__32291),
            .I(N__32258));
    InMux I__7711 (
            .O(N__32290),
            .I(N__32258));
    InMux I__7710 (
            .O(N__32289),
            .I(N__32251));
    InMux I__7709 (
            .O(N__32288),
            .I(N__32251));
    InMux I__7708 (
            .O(N__32287),
            .I(N__32251));
    InMux I__7707 (
            .O(N__32286),
            .I(N__32246));
    InMux I__7706 (
            .O(N__32285),
            .I(N__32246));
    CascadeMux I__7705 (
            .O(N__32284),
            .I(N__32223));
    CascadeMux I__7704 (
            .O(N__32283),
            .I(N__32213));
    CascadeMux I__7703 (
            .O(N__32282),
            .I(N__32208));
    Span4Mux_h I__7702 (
            .O(N__32279),
            .I(N__32184));
    LocalMux I__7701 (
            .O(N__32276),
            .I(N__32184));
    LocalMux I__7700 (
            .O(N__32273),
            .I(N__32184));
    LocalMux I__7699 (
            .O(N__32268),
            .I(N__32184));
    LocalMux I__7698 (
            .O(N__32265),
            .I(N__32184));
    LocalMux I__7697 (
            .O(N__32258),
            .I(N__32184));
    LocalMux I__7696 (
            .O(N__32251),
            .I(N__32184));
    LocalMux I__7695 (
            .O(N__32246),
            .I(N__32184));
    InMux I__7694 (
            .O(N__32245),
            .I(N__32179));
    InMux I__7693 (
            .O(N__32244),
            .I(N__32179));
    InMux I__7692 (
            .O(N__32243),
            .I(N__32174));
    InMux I__7691 (
            .O(N__32242),
            .I(N__32174));
    CascadeMux I__7690 (
            .O(N__32241),
            .I(N__32166));
    InMux I__7689 (
            .O(N__32240),
            .I(N__32157));
    InMux I__7688 (
            .O(N__32239),
            .I(N__32148));
    InMux I__7687 (
            .O(N__32238),
            .I(N__32148));
    InMux I__7686 (
            .O(N__32237),
            .I(N__32148));
    InMux I__7685 (
            .O(N__32236),
            .I(N__32148));
    CascadeMux I__7684 (
            .O(N__32235),
            .I(N__32145));
    InMux I__7683 (
            .O(N__32234),
            .I(N__32139));
    InMux I__7682 (
            .O(N__32233),
            .I(N__32136));
    InMux I__7681 (
            .O(N__32232),
            .I(N__32117));
    InMux I__7680 (
            .O(N__32231),
            .I(N__32117));
    InMux I__7679 (
            .O(N__32230),
            .I(N__32112));
    InMux I__7678 (
            .O(N__32229),
            .I(N__32112));
    InMux I__7677 (
            .O(N__32228),
            .I(N__32106));
    InMux I__7676 (
            .O(N__32227),
            .I(N__32106));
    InMux I__7675 (
            .O(N__32226),
            .I(N__32101));
    InMux I__7674 (
            .O(N__32223),
            .I(N__32101));
    CascadeMux I__7673 (
            .O(N__32222),
            .I(N__32096));
    CascadeMux I__7672 (
            .O(N__32221),
            .I(N__32093));
    InMux I__7671 (
            .O(N__32220),
            .I(N__32077));
    InMux I__7670 (
            .O(N__32219),
            .I(N__32077));
    InMux I__7669 (
            .O(N__32218),
            .I(N__32077));
    CascadeMux I__7668 (
            .O(N__32217),
            .I(N__32073));
    CascadeMux I__7667 (
            .O(N__32216),
            .I(N__32060));
    InMux I__7666 (
            .O(N__32213),
            .I(N__32049));
    InMux I__7665 (
            .O(N__32212),
            .I(N__32044));
    InMux I__7664 (
            .O(N__32211),
            .I(N__32044));
    InMux I__7663 (
            .O(N__32208),
            .I(N__32039));
    InMux I__7662 (
            .O(N__32207),
            .I(N__32039));
    InMux I__7661 (
            .O(N__32206),
            .I(N__32030));
    InMux I__7660 (
            .O(N__32205),
            .I(N__32030));
    InMux I__7659 (
            .O(N__32204),
            .I(N__32030));
    InMux I__7658 (
            .O(N__32203),
            .I(N__32030));
    InMux I__7657 (
            .O(N__32202),
            .I(N__32025));
    InMux I__7656 (
            .O(N__32201),
            .I(N__32025));
    Span4Mux_v I__7655 (
            .O(N__32184),
            .I(N__32021));
    LocalMux I__7654 (
            .O(N__32179),
            .I(N__32016));
    LocalMux I__7653 (
            .O(N__32174),
            .I(N__32016));
    InMux I__7652 (
            .O(N__32173),
            .I(N__32011));
    InMux I__7651 (
            .O(N__32172),
            .I(N__32011));
    CascadeMux I__7650 (
            .O(N__32171),
            .I(N__32008));
    CascadeMux I__7649 (
            .O(N__32170),
            .I(N__32001));
    InMux I__7648 (
            .O(N__32169),
            .I(N__31991));
    InMux I__7647 (
            .O(N__32166),
            .I(N__31986));
    InMux I__7646 (
            .O(N__32165),
            .I(N__31986));
    InMux I__7645 (
            .O(N__32164),
            .I(N__31975));
    InMux I__7644 (
            .O(N__32163),
            .I(N__31975));
    InMux I__7643 (
            .O(N__32162),
            .I(N__31975));
    InMux I__7642 (
            .O(N__32161),
            .I(N__31975));
    InMux I__7641 (
            .O(N__32160),
            .I(N__31975));
    LocalMux I__7640 (
            .O(N__32157),
            .I(N__31970));
    LocalMux I__7639 (
            .O(N__32148),
            .I(N__31970));
    InMux I__7638 (
            .O(N__32145),
            .I(N__31967));
    InMux I__7637 (
            .O(N__32144),
            .I(N__31964));
    InMux I__7636 (
            .O(N__32143),
            .I(N__31961));
    InMux I__7635 (
            .O(N__32142),
            .I(N__31958));
    LocalMux I__7634 (
            .O(N__32139),
            .I(N__31953));
    LocalMux I__7633 (
            .O(N__32136),
            .I(N__31953));
    InMux I__7632 (
            .O(N__32135),
            .I(N__31948));
    InMux I__7631 (
            .O(N__32134),
            .I(N__31948));
    InMux I__7630 (
            .O(N__32133),
            .I(N__31945));
    CascadeMux I__7629 (
            .O(N__32132),
            .I(N__31933));
    InMux I__7628 (
            .O(N__32131),
            .I(N__31927));
    InMux I__7627 (
            .O(N__32130),
            .I(N__31924));
    InMux I__7626 (
            .O(N__32129),
            .I(N__31919));
    InMux I__7625 (
            .O(N__32128),
            .I(N__31919));
    InMux I__7624 (
            .O(N__32127),
            .I(N__31916));
    InMux I__7623 (
            .O(N__32126),
            .I(N__31912));
    InMux I__7622 (
            .O(N__32125),
            .I(N__31909));
    InMux I__7621 (
            .O(N__32124),
            .I(N__31906));
    InMux I__7620 (
            .O(N__32123),
            .I(N__31901));
    InMux I__7619 (
            .O(N__32122),
            .I(N__31901));
    LocalMux I__7618 (
            .O(N__32117),
            .I(N__31896));
    LocalMux I__7617 (
            .O(N__32112),
            .I(N__31896));
    InMux I__7616 (
            .O(N__32111),
            .I(N__31893));
    LocalMux I__7615 (
            .O(N__32106),
            .I(N__31888));
    LocalMux I__7614 (
            .O(N__32101),
            .I(N__31888));
    CascadeMux I__7613 (
            .O(N__32100),
            .I(N__31884));
    InMux I__7612 (
            .O(N__32099),
            .I(N__31877));
    InMux I__7611 (
            .O(N__32096),
            .I(N__31877));
    InMux I__7610 (
            .O(N__32093),
            .I(N__31868));
    InMux I__7609 (
            .O(N__32092),
            .I(N__31868));
    InMux I__7608 (
            .O(N__32091),
            .I(N__31868));
    InMux I__7607 (
            .O(N__32090),
            .I(N__31868));
    InMux I__7606 (
            .O(N__32089),
            .I(N__31863));
    InMux I__7605 (
            .O(N__32088),
            .I(N__31863));
    InMux I__7604 (
            .O(N__32087),
            .I(N__31854));
    InMux I__7603 (
            .O(N__32086),
            .I(N__31854));
    InMux I__7602 (
            .O(N__32085),
            .I(N__31854));
    InMux I__7601 (
            .O(N__32084),
            .I(N__31854));
    LocalMux I__7600 (
            .O(N__32077),
            .I(N__31851));
    InMux I__7599 (
            .O(N__32076),
            .I(N__31840));
    InMux I__7598 (
            .O(N__32073),
            .I(N__31840));
    InMux I__7597 (
            .O(N__32072),
            .I(N__31835));
    InMux I__7596 (
            .O(N__32071),
            .I(N__31835));
    InMux I__7595 (
            .O(N__32070),
            .I(N__31830));
    InMux I__7594 (
            .O(N__32069),
            .I(N__31830));
    InMux I__7593 (
            .O(N__32068),
            .I(N__31821));
    InMux I__7592 (
            .O(N__32067),
            .I(N__31821));
    InMux I__7591 (
            .O(N__32066),
            .I(N__31821));
    InMux I__7590 (
            .O(N__32065),
            .I(N__31821));
    InMux I__7589 (
            .O(N__32064),
            .I(N__31818));
    InMux I__7588 (
            .O(N__32063),
            .I(N__31815));
    InMux I__7587 (
            .O(N__32060),
            .I(N__31804));
    InMux I__7586 (
            .O(N__32059),
            .I(N__31804));
    InMux I__7585 (
            .O(N__32058),
            .I(N__31804));
    InMux I__7584 (
            .O(N__32057),
            .I(N__31804));
    InMux I__7583 (
            .O(N__32056),
            .I(N__31804));
    InMux I__7582 (
            .O(N__32055),
            .I(N__31795));
    InMux I__7581 (
            .O(N__32054),
            .I(N__31795));
    InMux I__7580 (
            .O(N__32053),
            .I(N__31795));
    InMux I__7579 (
            .O(N__32052),
            .I(N__31795));
    LocalMux I__7578 (
            .O(N__32049),
            .I(N__31788));
    LocalMux I__7577 (
            .O(N__32044),
            .I(N__31788));
    LocalMux I__7576 (
            .O(N__32039),
            .I(N__31788));
    LocalMux I__7575 (
            .O(N__32030),
            .I(N__31785));
    LocalMux I__7574 (
            .O(N__32025),
            .I(N__31782));
    InMux I__7573 (
            .O(N__32024),
            .I(N__31779));
    Span4Mux_h I__7572 (
            .O(N__32021),
            .I(N__31772));
    Span4Mux_v I__7571 (
            .O(N__32016),
            .I(N__31772));
    LocalMux I__7570 (
            .O(N__32011),
            .I(N__31772));
    InMux I__7569 (
            .O(N__32008),
            .I(N__31769));
    InMux I__7568 (
            .O(N__32007),
            .I(N__31762));
    InMux I__7567 (
            .O(N__32006),
            .I(N__31762));
    InMux I__7566 (
            .O(N__32005),
            .I(N__31762));
    InMux I__7565 (
            .O(N__32004),
            .I(N__31751));
    InMux I__7564 (
            .O(N__32001),
            .I(N__31751));
    InMux I__7563 (
            .O(N__32000),
            .I(N__31751));
    InMux I__7562 (
            .O(N__31999),
            .I(N__31751));
    InMux I__7561 (
            .O(N__31998),
            .I(N__31751));
    InMux I__7560 (
            .O(N__31997),
            .I(N__31746));
    InMux I__7559 (
            .O(N__31996),
            .I(N__31746));
    InMux I__7558 (
            .O(N__31995),
            .I(N__31741));
    InMux I__7557 (
            .O(N__31994),
            .I(N__31741));
    LocalMux I__7556 (
            .O(N__31991),
            .I(N__31734));
    LocalMux I__7555 (
            .O(N__31986),
            .I(N__31734));
    LocalMux I__7554 (
            .O(N__31975),
            .I(N__31734));
    Span4Mux_h I__7553 (
            .O(N__31970),
            .I(N__31721));
    LocalMux I__7552 (
            .O(N__31967),
            .I(N__31721));
    LocalMux I__7551 (
            .O(N__31964),
            .I(N__31721));
    LocalMux I__7550 (
            .O(N__31961),
            .I(N__31721));
    LocalMux I__7549 (
            .O(N__31958),
            .I(N__31721));
    Span4Mux_v I__7548 (
            .O(N__31953),
            .I(N__31721));
    LocalMux I__7547 (
            .O(N__31948),
            .I(N__31716));
    LocalMux I__7546 (
            .O(N__31945),
            .I(N__31716));
    CascadeMux I__7545 (
            .O(N__31944),
            .I(N__31701));
    InMux I__7544 (
            .O(N__31943),
            .I(N__31694));
    InMux I__7543 (
            .O(N__31942),
            .I(N__31694));
    InMux I__7542 (
            .O(N__31941),
            .I(N__31689));
    InMux I__7541 (
            .O(N__31940),
            .I(N__31689));
    InMux I__7540 (
            .O(N__31939),
            .I(N__31680));
    InMux I__7539 (
            .O(N__31938),
            .I(N__31680));
    InMux I__7538 (
            .O(N__31937),
            .I(N__31680));
    InMux I__7537 (
            .O(N__31936),
            .I(N__31680));
    InMux I__7536 (
            .O(N__31933),
            .I(N__31671));
    InMux I__7535 (
            .O(N__31932),
            .I(N__31671));
    InMux I__7534 (
            .O(N__31931),
            .I(N__31671));
    InMux I__7533 (
            .O(N__31930),
            .I(N__31671));
    LocalMux I__7532 (
            .O(N__31927),
            .I(N__31662));
    LocalMux I__7531 (
            .O(N__31924),
            .I(N__31662));
    LocalMux I__7530 (
            .O(N__31919),
            .I(N__31662));
    LocalMux I__7529 (
            .O(N__31916),
            .I(N__31662));
    InMux I__7528 (
            .O(N__31915),
            .I(N__31659));
    LocalMux I__7527 (
            .O(N__31912),
            .I(N__31656));
    LocalMux I__7526 (
            .O(N__31909),
            .I(N__31651));
    LocalMux I__7525 (
            .O(N__31906),
            .I(N__31651));
    LocalMux I__7524 (
            .O(N__31901),
            .I(N__31646));
    Span4Mux_v I__7523 (
            .O(N__31896),
            .I(N__31646));
    LocalMux I__7522 (
            .O(N__31893),
            .I(N__31641));
    Span4Mux_v I__7521 (
            .O(N__31888),
            .I(N__31641));
    InMux I__7520 (
            .O(N__31887),
            .I(N__31632));
    InMux I__7519 (
            .O(N__31884),
            .I(N__31632));
    InMux I__7518 (
            .O(N__31883),
            .I(N__31632));
    InMux I__7517 (
            .O(N__31882),
            .I(N__31632));
    LocalMux I__7516 (
            .O(N__31877),
            .I(N__31621));
    LocalMux I__7515 (
            .O(N__31868),
            .I(N__31621));
    LocalMux I__7514 (
            .O(N__31863),
            .I(N__31621));
    LocalMux I__7513 (
            .O(N__31854),
            .I(N__31621));
    Span4Mux_h I__7512 (
            .O(N__31851),
            .I(N__31621));
    InMux I__7511 (
            .O(N__31850),
            .I(N__31618));
    InMux I__7510 (
            .O(N__31849),
            .I(N__31615));
    InMux I__7509 (
            .O(N__31848),
            .I(N__31606));
    InMux I__7508 (
            .O(N__31847),
            .I(N__31606));
    InMux I__7507 (
            .O(N__31846),
            .I(N__31606));
    InMux I__7506 (
            .O(N__31845),
            .I(N__31606));
    LocalMux I__7505 (
            .O(N__31840),
            .I(N__31595));
    LocalMux I__7504 (
            .O(N__31835),
            .I(N__31595));
    LocalMux I__7503 (
            .O(N__31830),
            .I(N__31595));
    LocalMux I__7502 (
            .O(N__31821),
            .I(N__31595));
    LocalMux I__7501 (
            .O(N__31818),
            .I(N__31595));
    LocalMux I__7500 (
            .O(N__31815),
            .I(N__31592));
    LocalMux I__7499 (
            .O(N__31804),
            .I(N__31581));
    LocalMux I__7498 (
            .O(N__31795),
            .I(N__31581));
    Span4Mux_h I__7497 (
            .O(N__31788),
            .I(N__31581));
    Span4Mux_h I__7496 (
            .O(N__31785),
            .I(N__31581));
    Span4Mux_h I__7495 (
            .O(N__31782),
            .I(N__31581));
    LocalMux I__7494 (
            .O(N__31779),
            .I(N__31578));
    Span4Mux_v I__7493 (
            .O(N__31772),
            .I(N__31575));
    LocalMux I__7492 (
            .O(N__31769),
            .I(N__31562));
    LocalMux I__7491 (
            .O(N__31762),
            .I(N__31562));
    LocalMux I__7490 (
            .O(N__31751),
            .I(N__31562));
    LocalMux I__7489 (
            .O(N__31746),
            .I(N__31562));
    LocalMux I__7488 (
            .O(N__31741),
            .I(N__31562));
    Span4Mux_h I__7487 (
            .O(N__31734),
            .I(N__31562));
    Span4Mux_v I__7486 (
            .O(N__31721),
            .I(N__31559));
    Span4Mux_v I__7485 (
            .O(N__31716),
            .I(N__31556));
    InMux I__7484 (
            .O(N__31715),
            .I(N__31551));
    InMux I__7483 (
            .O(N__31714),
            .I(N__31551));
    InMux I__7482 (
            .O(N__31713),
            .I(N__31548));
    InMux I__7481 (
            .O(N__31712),
            .I(N__31541));
    InMux I__7480 (
            .O(N__31711),
            .I(N__31541));
    InMux I__7479 (
            .O(N__31710),
            .I(N__31541));
    InMux I__7478 (
            .O(N__31709),
            .I(N__31530));
    InMux I__7477 (
            .O(N__31708),
            .I(N__31530));
    InMux I__7476 (
            .O(N__31707),
            .I(N__31530));
    InMux I__7475 (
            .O(N__31706),
            .I(N__31530));
    InMux I__7474 (
            .O(N__31705),
            .I(N__31530));
    InMux I__7473 (
            .O(N__31704),
            .I(N__31521));
    InMux I__7472 (
            .O(N__31701),
            .I(N__31521));
    InMux I__7471 (
            .O(N__31700),
            .I(N__31521));
    InMux I__7470 (
            .O(N__31699),
            .I(N__31521));
    LocalMux I__7469 (
            .O(N__31694),
            .I(N__31512));
    LocalMux I__7468 (
            .O(N__31689),
            .I(N__31512));
    LocalMux I__7467 (
            .O(N__31680),
            .I(N__31512));
    LocalMux I__7466 (
            .O(N__31671),
            .I(N__31512));
    Span4Mux_v I__7465 (
            .O(N__31662),
            .I(N__31509));
    LocalMux I__7464 (
            .O(N__31659),
            .I(N__31498));
    Span4Mux_v I__7463 (
            .O(N__31656),
            .I(N__31498));
    Span4Mux_v I__7462 (
            .O(N__31651),
            .I(N__31498));
    Span4Mux_h I__7461 (
            .O(N__31646),
            .I(N__31498));
    Span4Mux_h I__7460 (
            .O(N__31641),
            .I(N__31498));
    LocalMux I__7459 (
            .O(N__31632),
            .I(N__31493));
    Span4Mux_v I__7458 (
            .O(N__31621),
            .I(N__31493));
    LocalMux I__7457 (
            .O(N__31618),
            .I(N__31482));
    LocalMux I__7456 (
            .O(N__31615),
            .I(N__31482));
    LocalMux I__7455 (
            .O(N__31606),
            .I(N__31482));
    Span12Mux_v I__7454 (
            .O(N__31595),
            .I(N__31482));
    Span12Mux_v I__7453 (
            .O(N__31592),
            .I(N__31482));
    Span4Mux_v I__7452 (
            .O(N__31581),
            .I(N__31479));
    Span4Mux_v I__7451 (
            .O(N__31578),
            .I(N__31468));
    Span4Mux_h I__7450 (
            .O(N__31575),
            .I(N__31468));
    Span4Mux_v I__7449 (
            .O(N__31562),
            .I(N__31468));
    Span4Mux_h I__7448 (
            .O(N__31559),
            .I(N__31468));
    Span4Mux_h I__7447 (
            .O(N__31556),
            .I(N__31468));
    LocalMux I__7446 (
            .O(N__31551),
            .I(\c0.n1729 ));
    LocalMux I__7445 (
            .O(N__31548),
            .I(\c0.n1729 ));
    LocalMux I__7444 (
            .O(N__31541),
            .I(\c0.n1729 ));
    LocalMux I__7443 (
            .O(N__31530),
            .I(\c0.n1729 ));
    LocalMux I__7442 (
            .O(N__31521),
            .I(\c0.n1729 ));
    Odrv12 I__7441 (
            .O(N__31512),
            .I(\c0.n1729 ));
    Odrv4 I__7440 (
            .O(N__31509),
            .I(\c0.n1729 ));
    Odrv4 I__7439 (
            .O(N__31498),
            .I(\c0.n1729 ));
    Odrv4 I__7438 (
            .O(N__31493),
            .I(\c0.n1729 ));
    Odrv12 I__7437 (
            .O(N__31482),
            .I(\c0.n1729 ));
    Odrv4 I__7436 (
            .O(N__31479),
            .I(\c0.n1729 ));
    Odrv4 I__7435 (
            .O(N__31468),
            .I(\c0.n1729 ));
    InMux I__7434 (
            .O(N__31443),
            .I(N__31440));
    LocalMux I__7433 (
            .O(N__31440),
            .I(N__31437));
    Span4Mux_h I__7432 (
            .O(N__31437),
            .I(N__31433));
    InMux I__7431 (
            .O(N__31436),
            .I(N__31429));
    Span4Mux_h I__7430 (
            .O(N__31433),
            .I(N__31426));
    InMux I__7429 (
            .O(N__31432),
            .I(N__31423));
    LocalMux I__7428 (
            .O(N__31429),
            .I(data_in_4_7));
    Odrv4 I__7427 (
            .O(N__31426),
            .I(data_in_4_7));
    LocalMux I__7426 (
            .O(N__31423),
            .I(data_in_4_7));
    InMux I__7425 (
            .O(N__31416),
            .I(N__31413));
    LocalMux I__7424 (
            .O(N__31413),
            .I(N__31408));
    CascadeMux I__7423 (
            .O(N__31412),
            .I(N__31404));
    InMux I__7422 (
            .O(N__31411),
            .I(N__31401));
    Span4Mux_v I__7421 (
            .O(N__31408),
            .I(N__31397));
    CascadeMux I__7420 (
            .O(N__31407),
            .I(N__31394));
    InMux I__7419 (
            .O(N__31404),
            .I(N__31391));
    LocalMux I__7418 (
            .O(N__31401),
            .I(N__31388));
    InMux I__7417 (
            .O(N__31400),
            .I(N__31385));
    Span4Mux_h I__7416 (
            .O(N__31397),
            .I(N__31382));
    InMux I__7415 (
            .O(N__31394),
            .I(N__31379));
    LocalMux I__7414 (
            .O(N__31391),
            .I(\c0.data_in_field_39 ));
    Odrv4 I__7413 (
            .O(N__31388),
            .I(\c0.data_in_field_39 ));
    LocalMux I__7412 (
            .O(N__31385),
            .I(\c0.data_in_field_39 ));
    Odrv4 I__7411 (
            .O(N__31382),
            .I(\c0.data_in_field_39 ));
    LocalMux I__7410 (
            .O(N__31379),
            .I(\c0.data_in_field_39 ));
    InMux I__7409 (
            .O(N__31368),
            .I(N__31364));
    InMux I__7408 (
            .O(N__31367),
            .I(N__31361));
    LocalMux I__7407 (
            .O(N__31364),
            .I(N__31358));
    LocalMux I__7406 (
            .O(N__31361),
            .I(N__31354));
    Span4Mux_h I__7405 (
            .O(N__31358),
            .I(N__31351));
    InMux I__7404 (
            .O(N__31357),
            .I(N__31348));
    Odrv12 I__7403 (
            .O(N__31354),
            .I(data_in_10_7));
    Odrv4 I__7402 (
            .O(N__31351),
            .I(data_in_10_7));
    LocalMux I__7401 (
            .O(N__31348),
            .I(data_in_10_7));
    InMux I__7400 (
            .O(N__31341),
            .I(N__31338));
    LocalMux I__7399 (
            .O(N__31338),
            .I(N__31334));
    InMux I__7398 (
            .O(N__31337),
            .I(N__31331));
    Span4Mux_v I__7397 (
            .O(N__31334),
            .I(N__31326));
    LocalMux I__7396 (
            .O(N__31331),
            .I(N__31326));
    Sp12to4 I__7395 (
            .O(N__31326),
            .I(N__31323));
    Span12Mux_s11_v I__7394 (
            .O(N__31323),
            .I(N__31319));
    InMux I__7393 (
            .O(N__31322),
            .I(N__31316));
    Odrv12 I__7392 (
            .O(N__31319),
            .I(data_in_9_7));
    LocalMux I__7391 (
            .O(N__31316),
            .I(data_in_9_7));
    CascadeMux I__7390 (
            .O(N__31311),
            .I(N__31307));
    InMux I__7389 (
            .O(N__31310),
            .I(N__31304));
    InMux I__7388 (
            .O(N__31307),
            .I(N__31301));
    LocalMux I__7387 (
            .O(N__31304),
            .I(N__31298));
    LocalMux I__7386 (
            .O(N__31301),
            .I(N__31294));
    Span4Mux_h I__7385 (
            .O(N__31298),
            .I(N__31291));
    InMux I__7384 (
            .O(N__31297),
            .I(N__31288));
    Odrv12 I__7383 (
            .O(N__31294),
            .I(data_in_14_5));
    Odrv4 I__7382 (
            .O(N__31291),
            .I(data_in_14_5));
    LocalMux I__7381 (
            .O(N__31288),
            .I(data_in_14_5));
    CascadeMux I__7380 (
            .O(N__31281),
            .I(N__31278));
    InMux I__7379 (
            .O(N__31278),
            .I(N__31271));
    InMux I__7378 (
            .O(N__31277),
            .I(N__31271));
    InMux I__7377 (
            .O(N__31276),
            .I(N__31268));
    LocalMux I__7376 (
            .O(N__31271),
            .I(N__31265));
    LocalMux I__7375 (
            .O(N__31268),
            .I(data_in_12_2));
    Odrv4 I__7374 (
            .O(N__31265),
            .I(data_in_12_2));
    CascadeMux I__7373 (
            .O(N__31260),
            .I(N__31257));
    InMux I__7372 (
            .O(N__31257),
            .I(N__31254));
    LocalMux I__7371 (
            .O(N__31254),
            .I(N__31250));
    InMux I__7370 (
            .O(N__31253),
            .I(N__31247));
    Span4Mux_v I__7369 (
            .O(N__31250),
            .I(N__31243));
    LocalMux I__7368 (
            .O(N__31247),
            .I(N__31240));
    InMux I__7367 (
            .O(N__31246),
            .I(N__31237));
    Odrv4 I__7366 (
            .O(N__31243),
            .I(data_in_11_2));
    Odrv4 I__7365 (
            .O(N__31240),
            .I(data_in_11_2));
    LocalMux I__7364 (
            .O(N__31237),
            .I(data_in_11_2));
    CascadeMux I__7363 (
            .O(N__31230),
            .I(N__31227));
    InMux I__7362 (
            .O(N__31227),
            .I(N__31224));
    LocalMux I__7361 (
            .O(N__31224),
            .I(N__31220));
    InMux I__7360 (
            .O(N__31223),
            .I(N__31217));
    Span4Mux_h I__7359 (
            .O(N__31220),
            .I(N__31214));
    LocalMux I__7358 (
            .O(N__31217),
            .I(N__31211));
    Span4Mux_h I__7357 (
            .O(N__31214),
            .I(N__31205));
    Span4Mux_h I__7356 (
            .O(N__31211),
            .I(N__31205));
    InMux I__7355 (
            .O(N__31210),
            .I(N__31202));
    Odrv4 I__7354 (
            .O(N__31205),
            .I(data_in_4_4));
    LocalMux I__7353 (
            .O(N__31202),
            .I(data_in_4_4));
    InMux I__7352 (
            .O(N__31197),
            .I(N__31194));
    LocalMux I__7351 (
            .O(N__31194),
            .I(N__31190));
    InMux I__7350 (
            .O(N__31193),
            .I(N__31187));
    Span4Mux_v I__7349 (
            .O(N__31190),
            .I(N__31184));
    LocalMux I__7348 (
            .O(N__31187),
            .I(N__31178));
    Sp12to4 I__7347 (
            .O(N__31184),
            .I(N__31178));
    InMux I__7346 (
            .O(N__31183),
            .I(N__31175));
    Odrv12 I__7345 (
            .O(N__31178),
            .I(data_in_9_6));
    LocalMux I__7344 (
            .O(N__31175),
            .I(data_in_9_6));
    InMux I__7343 (
            .O(N__31170),
            .I(N__31166));
    CascadeMux I__7342 (
            .O(N__31169),
            .I(N__31163));
    LocalMux I__7341 (
            .O(N__31166),
            .I(N__31160));
    InMux I__7340 (
            .O(N__31163),
            .I(N__31157));
    Span4Mux_v I__7339 (
            .O(N__31160),
            .I(N__31154));
    LocalMux I__7338 (
            .O(N__31157),
            .I(N__31150));
    Span4Mux_h I__7337 (
            .O(N__31154),
            .I(N__31147));
    InMux I__7336 (
            .O(N__31153),
            .I(N__31144));
    Odrv12 I__7335 (
            .O(N__31150),
            .I(data_in_8_6));
    Odrv4 I__7334 (
            .O(N__31147),
            .I(data_in_8_6));
    LocalMux I__7333 (
            .O(N__31144),
            .I(data_in_8_6));
    CascadeMux I__7332 (
            .O(N__31137),
            .I(N__31134));
    InMux I__7331 (
            .O(N__31134),
            .I(N__31131));
    LocalMux I__7330 (
            .O(N__31131),
            .I(N__31127));
    CascadeMux I__7329 (
            .O(N__31130),
            .I(N__31122));
    Span4Mux_h I__7328 (
            .O(N__31127),
            .I(N__31119));
    InMux I__7327 (
            .O(N__31126),
            .I(N__31114));
    InMux I__7326 (
            .O(N__31125),
            .I(N__31114));
    InMux I__7325 (
            .O(N__31122),
            .I(N__31111));
    Odrv4 I__7324 (
            .O(N__31119),
            .I(data_in_3_4));
    LocalMux I__7323 (
            .O(N__31114),
            .I(data_in_3_4));
    LocalMux I__7322 (
            .O(N__31111),
            .I(data_in_3_4));
    InMux I__7321 (
            .O(N__31104),
            .I(N__31099));
    InMux I__7320 (
            .O(N__31103),
            .I(N__31096));
    InMux I__7319 (
            .O(N__31102),
            .I(N__31093));
    LocalMux I__7318 (
            .O(N__31099),
            .I(N__31090));
    LocalMux I__7317 (
            .O(N__31096),
            .I(N__31084));
    LocalMux I__7316 (
            .O(N__31093),
            .I(N__31084));
    Span4Mux_v I__7315 (
            .O(N__31090),
            .I(N__31081));
    InMux I__7314 (
            .O(N__31089),
            .I(N__31078));
    Span4Mux_h I__7313 (
            .O(N__31084),
            .I(N__31075));
    Odrv4 I__7312 (
            .O(N__31081),
            .I(data_in_2_4));
    LocalMux I__7311 (
            .O(N__31078),
            .I(data_in_2_4));
    Odrv4 I__7310 (
            .O(N__31075),
            .I(data_in_2_4));
    InMux I__7309 (
            .O(N__31068),
            .I(N__31065));
    LocalMux I__7308 (
            .O(N__31065),
            .I(\c0.n50_adj_1875 ));
    InMux I__7307 (
            .O(N__31062),
            .I(N__31059));
    LocalMux I__7306 (
            .O(N__31059),
            .I(N__31055));
    InMux I__7305 (
            .O(N__31058),
            .I(N__31052));
    Span4Mux_h I__7304 (
            .O(N__31055),
            .I(N__31049));
    LocalMux I__7303 (
            .O(N__31052),
            .I(N__31046));
    Span4Mux_h I__7302 (
            .O(N__31049),
            .I(N__31040));
    Span4Mux_h I__7301 (
            .O(N__31046),
            .I(N__31040));
    InMux I__7300 (
            .O(N__31045),
            .I(N__31037));
    Odrv4 I__7299 (
            .O(N__31040),
            .I(data_in_8_0));
    LocalMux I__7298 (
            .O(N__31037),
            .I(data_in_8_0));
    CascadeMux I__7297 (
            .O(N__31032),
            .I(N__31028));
    InMux I__7296 (
            .O(N__31031),
            .I(N__31024));
    InMux I__7295 (
            .O(N__31028),
            .I(N__31019));
    InMux I__7294 (
            .O(N__31027),
            .I(N__31019));
    LocalMux I__7293 (
            .O(N__31024),
            .I(data_in_7_0));
    LocalMux I__7292 (
            .O(N__31019),
            .I(data_in_7_0));
    InMux I__7291 (
            .O(N__31014),
            .I(N__31010));
    InMux I__7290 (
            .O(N__31013),
            .I(N__31007));
    LocalMux I__7289 (
            .O(N__31010),
            .I(N__31004));
    LocalMux I__7288 (
            .O(N__31007),
            .I(N__31001));
    Span4Mux_v I__7287 (
            .O(N__31004),
            .I(N__30997));
    Span4Mux_v I__7286 (
            .O(N__31001),
            .I(N__30994));
    InMux I__7285 (
            .O(N__31000),
            .I(N__30990));
    Span4Mux_h I__7284 (
            .O(N__30997),
            .I(N__30985));
    Span4Mux_h I__7283 (
            .O(N__30994),
            .I(N__30985));
    InMux I__7282 (
            .O(N__30993),
            .I(N__30982));
    LocalMux I__7281 (
            .O(N__30990),
            .I(\c0.data_in_field_74 ));
    Odrv4 I__7280 (
            .O(N__30985),
            .I(\c0.data_in_field_74 ));
    LocalMux I__7279 (
            .O(N__30982),
            .I(\c0.data_in_field_74 ));
    InMux I__7278 (
            .O(N__30975),
            .I(N__30971));
    InMux I__7277 (
            .O(N__30974),
            .I(N__30968));
    LocalMux I__7276 (
            .O(N__30971),
            .I(N__30963));
    LocalMux I__7275 (
            .O(N__30968),
            .I(N__30960));
    CascadeMux I__7274 (
            .O(N__30967),
            .I(N__30957));
    InMux I__7273 (
            .O(N__30966),
            .I(N__30954));
    Span4Mux_v I__7272 (
            .O(N__30963),
            .I(N__30951));
    Span12Mux_h I__7271 (
            .O(N__30960),
            .I(N__30948));
    InMux I__7270 (
            .O(N__30957),
            .I(N__30945));
    LocalMux I__7269 (
            .O(N__30954),
            .I(\c0.data_in_field_1 ));
    Odrv4 I__7268 (
            .O(N__30951),
            .I(\c0.data_in_field_1 ));
    Odrv12 I__7267 (
            .O(N__30948),
            .I(\c0.data_in_field_1 ));
    LocalMux I__7266 (
            .O(N__30945),
            .I(\c0.data_in_field_1 ));
    CascadeMux I__7265 (
            .O(N__30936),
            .I(N__30930));
    CascadeMux I__7264 (
            .O(N__30935),
            .I(N__30927));
    InMux I__7263 (
            .O(N__30934),
            .I(N__30923));
    InMux I__7262 (
            .O(N__30933),
            .I(N__30920));
    InMux I__7261 (
            .O(N__30930),
            .I(N__30917));
    InMux I__7260 (
            .O(N__30927),
            .I(N__30912));
    InMux I__7259 (
            .O(N__30926),
            .I(N__30912));
    LocalMux I__7258 (
            .O(N__30923),
            .I(\c0.data_in_field_16 ));
    LocalMux I__7257 (
            .O(N__30920),
            .I(\c0.data_in_field_16 ));
    LocalMux I__7256 (
            .O(N__30917),
            .I(\c0.data_in_field_16 ));
    LocalMux I__7255 (
            .O(N__30912),
            .I(\c0.data_in_field_16 ));
    InMux I__7254 (
            .O(N__30903),
            .I(N__30900));
    LocalMux I__7253 (
            .O(N__30900),
            .I(\c0.n25_adj_1931 ));
    InMux I__7252 (
            .O(N__30897),
            .I(N__30893));
    InMux I__7251 (
            .O(N__30896),
            .I(N__30889));
    LocalMux I__7250 (
            .O(N__30893),
            .I(N__30886));
    InMux I__7249 (
            .O(N__30892),
            .I(N__30883));
    LocalMux I__7248 (
            .O(N__30889),
            .I(N__30878));
    Span4Mux_v I__7247 (
            .O(N__30886),
            .I(N__30875));
    LocalMux I__7246 (
            .O(N__30883),
            .I(N__30872));
    CascadeMux I__7245 (
            .O(N__30882),
            .I(N__30869));
    InMux I__7244 (
            .O(N__30881),
            .I(N__30866));
    Span4Mux_v I__7243 (
            .O(N__30878),
            .I(N__30863));
    Span4Mux_h I__7242 (
            .O(N__30875),
            .I(N__30858));
    Span4Mux_v I__7241 (
            .O(N__30872),
            .I(N__30858));
    InMux I__7240 (
            .O(N__30869),
            .I(N__30855));
    LocalMux I__7239 (
            .O(N__30866),
            .I(\c0.data_in_field_137 ));
    Odrv4 I__7238 (
            .O(N__30863),
            .I(\c0.data_in_field_137 ));
    Odrv4 I__7237 (
            .O(N__30858),
            .I(\c0.data_in_field_137 ));
    LocalMux I__7236 (
            .O(N__30855),
            .I(\c0.data_in_field_137 ));
    CascadeMux I__7235 (
            .O(N__30846),
            .I(N__30842));
    CascadeMux I__7234 (
            .O(N__30845),
            .I(N__30839));
    InMux I__7233 (
            .O(N__30842),
            .I(N__30836));
    InMux I__7232 (
            .O(N__30839),
            .I(N__30833));
    LocalMux I__7231 (
            .O(N__30836),
            .I(N__30830));
    LocalMux I__7230 (
            .O(N__30833),
            .I(N__30825));
    Span4Mux_v I__7229 (
            .O(N__30830),
            .I(N__30822));
    InMux I__7228 (
            .O(N__30829),
            .I(N__30818));
    CascadeMux I__7227 (
            .O(N__30828),
            .I(N__30815));
    Span4Mux_v I__7226 (
            .O(N__30825),
            .I(N__30812));
    Span4Mux_h I__7225 (
            .O(N__30822),
            .I(N__30809));
    CascadeMux I__7224 (
            .O(N__30821),
            .I(N__30806));
    LocalMux I__7223 (
            .O(N__30818),
            .I(N__30803));
    InMux I__7222 (
            .O(N__30815),
            .I(N__30800));
    Span4Mux_v I__7221 (
            .O(N__30812),
            .I(N__30795));
    Span4Mux_h I__7220 (
            .O(N__30809),
            .I(N__30795));
    InMux I__7219 (
            .O(N__30806),
            .I(N__30792));
    Span4Mux_h I__7218 (
            .O(N__30803),
            .I(N__30789));
    LocalMux I__7217 (
            .O(N__30800),
            .I(\c0.data_in_field_25 ));
    Odrv4 I__7216 (
            .O(N__30795),
            .I(\c0.data_in_field_25 ));
    LocalMux I__7215 (
            .O(N__30792),
            .I(\c0.data_in_field_25 ));
    Odrv4 I__7214 (
            .O(N__30789),
            .I(\c0.data_in_field_25 ));
    InMux I__7213 (
            .O(N__30780),
            .I(N__30776));
    InMux I__7212 (
            .O(N__30779),
            .I(N__30772));
    LocalMux I__7211 (
            .O(N__30776),
            .I(N__30769));
    CascadeMux I__7210 (
            .O(N__30775),
            .I(N__30765));
    LocalMux I__7209 (
            .O(N__30772),
            .I(N__30762));
    Span4Mux_v I__7208 (
            .O(N__30769),
            .I(N__30759));
    CascadeMux I__7207 (
            .O(N__30768),
            .I(N__30756));
    InMux I__7206 (
            .O(N__30765),
            .I(N__30753));
    Span4Mux_h I__7205 (
            .O(N__30762),
            .I(N__30750));
    Span4Mux_h I__7204 (
            .O(N__30759),
            .I(N__30747));
    InMux I__7203 (
            .O(N__30756),
            .I(N__30744));
    LocalMux I__7202 (
            .O(N__30753),
            .I(\c0.data_in_field_71 ));
    Odrv4 I__7201 (
            .O(N__30750),
            .I(\c0.data_in_field_71 ));
    Odrv4 I__7200 (
            .O(N__30747),
            .I(\c0.data_in_field_71 ));
    LocalMux I__7199 (
            .O(N__30744),
            .I(\c0.data_in_field_71 ));
    InMux I__7198 (
            .O(N__30735),
            .I(N__30731));
    CascadeMux I__7197 (
            .O(N__30734),
            .I(N__30728));
    LocalMux I__7196 (
            .O(N__30731),
            .I(N__30725));
    InMux I__7195 (
            .O(N__30728),
            .I(N__30722));
    Span4Mux_h I__7194 (
            .O(N__30725),
            .I(N__30719));
    LocalMux I__7193 (
            .O(N__30722),
            .I(N__30716));
    Span4Mux_h I__7192 (
            .O(N__30719),
            .I(N__30713));
    Span4Mux_h I__7191 (
            .O(N__30716),
            .I(N__30710));
    Odrv4 I__7190 (
            .O(N__30713),
            .I(\c0.n5542 ));
    Odrv4 I__7189 (
            .O(N__30710),
            .I(\c0.n5542 ));
    CascadeMux I__7188 (
            .O(N__30705),
            .I(N__30702));
    InMux I__7187 (
            .O(N__30702),
            .I(N__30699));
    LocalMux I__7186 (
            .O(N__30699),
            .I(N__30696));
    Span4Mux_v I__7185 (
            .O(N__30696),
            .I(N__30691));
    InMux I__7184 (
            .O(N__30695),
            .I(N__30688));
    InMux I__7183 (
            .O(N__30694),
            .I(N__30685));
    Odrv4 I__7182 (
            .O(N__30691),
            .I(data_in_17_0));
    LocalMux I__7181 (
            .O(N__30688),
            .I(data_in_17_0));
    LocalMux I__7180 (
            .O(N__30685),
            .I(data_in_17_0));
    CascadeMux I__7179 (
            .O(N__30678),
            .I(N__30675));
    InMux I__7178 (
            .O(N__30675),
            .I(N__30672));
    LocalMux I__7177 (
            .O(N__30672),
            .I(N__30668));
    InMux I__7176 (
            .O(N__30671),
            .I(N__30665));
    Span4Mux_h I__7175 (
            .O(N__30668),
            .I(N__30662));
    LocalMux I__7174 (
            .O(N__30665),
            .I(N__30659));
    Span4Mux_h I__7173 (
            .O(N__30662),
            .I(N__30655));
    Span12Mux_v I__7172 (
            .O(N__30659),
            .I(N__30652));
    InMux I__7171 (
            .O(N__30658),
            .I(N__30649));
    Odrv4 I__7170 (
            .O(N__30655),
            .I(data_in_10_2));
    Odrv12 I__7169 (
            .O(N__30652),
            .I(data_in_10_2));
    LocalMux I__7168 (
            .O(N__30649),
            .I(data_in_10_2));
    CascadeMux I__7167 (
            .O(N__30642),
            .I(N__30639));
    InMux I__7166 (
            .O(N__30639),
            .I(N__30636));
    LocalMux I__7165 (
            .O(N__30636),
            .I(N__30633));
    Span4Mux_h I__7164 (
            .O(N__30633),
            .I(N__30630));
    Span4Mux_v I__7163 (
            .O(N__30630),
            .I(N__30625));
    InMux I__7162 (
            .O(N__30629),
            .I(N__30620));
    InMux I__7161 (
            .O(N__30628),
            .I(N__30620));
    Odrv4 I__7160 (
            .O(N__30625),
            .I(data_in_4_6));
    LocalMux I__7159 (
            .O(N__30620),
            .I(data_in_4_6));
    InMux I__7158 (
            .O(N__30615),
            .I(N__30611));
    InMux I__7157 (
            .O(N__30614),
            .I(N__30608));
    LocalMux I__7156 (
            .O(N__30611),
            .I(N__30600));
    LocalMux I__7155 (
            .O(N__30608),
            .I(N__30600));
    InMux I__7154 (
            .O(N__30607),
            .I(N__30597));
    CascadeMux I__7153 (
            .O(N__30606),
            .I(N__30594));
    InMux I__7152 (
            .O(N__30605),
            .I(N__30590));
    Span12Mux_v I__7151 (
            .O(N__30600),
            .I(N__30585));
    LocalMux I__7150 (
            .O(N__30597),
            .I(N__30585));
    InMux I__7149 (
            .O(N__30594),
            .I(N__30580));
    InMux I__7148 (
            .O(N__30593),
            .I(N__30580));
    LocalMux I__7147 (
            .O(N__30590),
            .I(\c0.data_in_field_38 ));
    Odrv12 I__7146 (
            .O(N__30585),
            .I(\c0.data_in_field_38 ));
    LocalMux I__7145 (
            .O(N__30580),
            .I(\c0.data_in_field_38 ));
    InMux I__7144 (
            .O(N__30573),
            .I(N__30570));
    LocalMux I__7143 (
            .O(N__30570),
            .I(N__30565));
    InMux I__7142 (
            .O(N__30569),
            .I(N__30562));
    InMux I__7141 (
            .O(N__30568),
            .I(N__30557));
    Span12Mux_h I__7140 (
            .O(N__30565),
            .I(N__30554));
    LocalMux I__7139 (
            .O(N__30562),
            .I(N__30551));
    InMux I__7138 (
            .O(N__30561),
            .I(N__30548));
    InMux I__7137 (
            .O(N__30560),
            .I(N__30545));
    LocalMux I__7136 (
            .O(N__30557),
            .I(\c0.data_in_field_136 ));
    Odrv12 I__7135 (
            .O(N__30554),
            .I(\c0.data_in_field_136 ));
    Odrv4 I__7134 (
            .O(N__30551),
            .I(\c0.data_in_field_136 ));
    LocalMux I__7133 (
            .O(N__30548),
            .I(\c0.data_in_field_136 ));
    LocalMux I__7132 (
            .O(N__30545),
            .I(\c0.data_in_field_136 ));
    InMux I__7131 (
            .O(N__30534),
            .I(N__30531));
    LocalMux I__7130 (
            .O(N__30531),
            .I(N__30526));
    InMux I__7129 (
            .O(N__30530),
            .I(N__30523));
    InMux I__7128 (
            .O(N__30529),
            .I(N__30519));
    Span4Mux_v I__7127 (
            .O(N__30526),
            .I(N__30515));
    LocalMux I__7126 (
            .O(N__30523),
            .I(N__30512));
    InMux I__7125 (
            .O(N__30522),
            .I(N__30509));
    LocalMux I__7124 (
            .O(N__30519),
            .I(N__30506));
    InMux I__7123 (
            .O(N__30518),
            .I(N__30503));
    Sp12to4 I__7122 (
            .O(N__30515),
            .I(N__30498));
    Sp12to4 I__7121 (
            .O(N__30512),
            .I(N__30498));
    LocalMux I__7120 (
            .O(N__30509),
            .I(\c0.data_in_field_31 ));
    Odrv12 I__7119 (
            .O(N__30506),
            .I(\c0.data_in_field_31 ));
    LocalMux I__7118 (
            .O(N__30503),
            .I(\c0.data_in_field_31 ));
    Odrv12 I__7117 (
            .O(N__30498),
            .I(\c0.data_in_field_31 ));
    InMux I__7116 (
            .O(N__30489),
            .I(N__30486));
    LocalMux I__7115 (
            .O(N__30486),
            .I(\c0.n2113 ));
    CascadeMux I__7114 (
            .O(N__30483),
            .I(N__30479));
    InMux I__7113 (
            .O(N__30482),
            .I(N__30476));
    InMux I__7112 (
            .O(N__30479),
            .I(N__30473));
    LocalMux I__7111 (
            .O(N__30476),
            .I(N__30470));
    LocalMux I__7110 (
            .O(N__30473),
            .I(N__30466));
    Span4Mux_h I__7109 (
            .O(N__30470),
            .I(N__30463));
    InMux I__7108 (
            .O(N__30469),
            .I(N__30460));
    Odrv4 I__7107 (
            .O(N__30466),
            .I(data_in_11_0));
    Odrv4 I__7106 (
            .O(N__30463),
            .I(data_in_11_0));
    LocalMux I__7105 (
            .O(N__30460),
            .I(data_in_11_0));
    InMux I__7104 (
            .O(N__30453),
            .I(N__30449));
    InMux I__7103 (
            .O(N__30452),
            .I(N__30446));
    LocalMux I__7102 (
            .O(N__30449),
            .I(N__30443));
    LocalMux I__7101 (
            .O(N__30446),
            .I(N__30440));
    Span4Mux_v I__7100 (
            .O(N__30443),
            .I(N__30434));
    Span4Mux_v I__7099 (
            .O(N__30440),
            .I(N__30434));
    InMux I__7098 (
            .O(N__30439),
            .I(N__30431));
    Span4Mux_h I__7097 (
            .O(N__30434),
            .I(N__30428));
    LocalMux I__7096 (
            .O(N__30431),
            .I(data_in_10_0));
    Odrv4 I__7095 (
            .O(N__30428),
            .I(data_in_10_0));
    CascadeMux I__7094 (
            .O(N__30423),
            .I(N__30420));
    InMux I__7093 (
            .O(N__30420),
            .I(N__30416));
    InMux I__7092 (
            .O(N__30419),
            .I(N__30413));
    LocalMux I__7091 (
            .O(N__30416),
            .I(N__30410));
    LocalMux I__7090 (
            .O(N__30413),
            .I(N__30407));
    Span4Mux_h I__7089 (
            .O(N__30410),
            .I(N__30403));
    Span4Mux_h I__7088 (
            .O(N__30407),
            .I(N__30400));
    InMux I__7087 (
            .O(N__30406),
            .I(N__30397));
    Odrv4 I__7086 (
            .O(N__30403),
            .I(data_in_10_4));
    Odrv4 I__7085 (
            .O(N__30400),
            .I(data_in_10_4));
    LocalMux I__7084 (
            .O(N__30397),
            .I(data_in_10_4));
    InMux I__7083 (
            .O(N__30390),
            .I(N__30387));
    LocalMux I__7082 (
            .O(N__30387),
            .I(N__30383));
    InMux I__7081 (
            .O(N__30386),
            .I(N__30380));
    Span4Mux_h I__7080 (
            .O(N__30383),
            .I(N__30377));
    LocalMux I__7079 (
            .O(N__30380),
            .I(N__30374));
    Span4Mux_h I__7078 (
            .O(N__30377),
            .I(N__30371));
    Span4Mux_v I__7077 (
            .O(N__30374),
            .I(N__30368));
    Span4Mux_v I__7076 (
            .O(N__30371),
            .I(N__30364));
    Span4Mux_h I__7075 (
            .O(N__30368),
            .I(N__30361));
    InMux I__7074 (
            .O(N__30367),
            .I(N__30358));
    Odrv4 I__7073 (
            .O(N__30364),
            .I(data_in_9_4));
    Odrv4 I__7072 (
            .O(N__30361),
            .I(data_in_9_4));
    LocalMux I__7071 (
            .O(N__30358),
            .I(data_in_9_4));
    CascadeMux I__7070 (
            .O(N__30351),
            .I(N__30348));
    InMux I__7069 (
            .O(N__30348),
            .I(N__30345));
    LocalMux I__7068 (
            .O(N__30345),
            .I(N__30342));
    Span4Mux_h I__7067 (
            .O(N__30342),
            .I(N__30337));
    InMux I__7066 (
            .O(N__30341),
            .I(N__30334));
    InMux I__7065 (
            .O(N__30340),
            .I(N__30331));
    Odrv4 I__7064 (
            .O(N__30337),
            .I(data_in_16_4));
    LocalMux I__7063 (
            .O(N__30334),
            .I(data_in_16_4));
    LocalMux I__7062 (
            .O(N__30331),
            .I(data_in_16_4));
    CascadeMux I__7061 (
            .O(N__30324),
            .I(N__30321));
    InMux I__7060 (
            .O(N__30321),
            .I(N__30318));
    LocalMux I__7059 (
            .O(N__30318),
            .I(N__30315));
    Span4Mux_h I__7058 (
            .O(N__30315),
            .I(N__30312));
    Span4Mux_h I__7057 (
            .O(N__30312),
            .I(N__30309));
    Span4Mux_h I__7056 (
            .O(N__30309),
            .I(N__30304));
    InMux I__7055 (
            .O(N__30308),
            .I(N__30301));
    InMux I__7054 (
            .O(N__30307),
            .I(N__30298));
    Odrv4 I__7053 (
            .O(N__30304),
            .I(data_in_15_4));
    LocalMux I__7052 (
            .O(N__30301),
            .I(data_in_15_4));
    LocalMux I__7051 (
            .O(N__30298),
            .I(data_in_15_4));
    CascadeMux I__7050 (
            .O(N__30291),
            .I(N__30287));
    CascadeMux I__7049 (
            .O(N__30290),
            .I(N__30284));
    InMux I__7048 (
            .O(N__30287),
            .I(N__30281));
    InMux I__7047 (
            .O(N__30284),
            .I(N__30277));
    LocalMux I__7046 (
            .O(N__30281),
            .I(N__30274));
    InMux I__7045 (
            .O(N__30280),
            .I(N__30271));
    LocalMux I__7044 (
            .O(N__30277),
            .I(data_in_13_4));
    Odrv4 I__7043 (
            .O(N__30274),
            .I(data_in_13_4));
    LocalMux I__7042 (
            .O(N__30271),
            .I(data_in_13_4));
    CascadeMux I__7041 (
            .O(N__30264),
            .I(N__30261));
    InMux I__7040 (
            .O(N__30261),
            .I(N__30257));
    InMux I__7039 (
            .O(N__30260),
            .I(N__30254));
    LocalMux I__7038 (
            .O(N__30257),
            .I(N__30251));
    LocalMux I__7037 (
            .O(N__30254),
            .I(N__30247));
    Span4Mux_v I__7036 (
            .O(N__30251),
            .I(N__30244));
    InMux I__7035 (
            .O(N__30250),
            .I(N__30240));
    Span4Mux_h I__7034 (
            .O(N__30247),
            .I(N__30237));
    Span4Mux_v I__7033 (
            .O(N__30244),
            .I(N__30234));
    InMux I__7032 (
            .O(N__30243),
            .I(N__30231));
    LocalMux I__7031 (
            .O(N__30240),
            .I(N__30225));
    Span4Mux_v I__7030 (
            .O(N__30237),
            .I(N__30225));
    Span4Mux_h I__7029 (
            .O(N__30234),
            .I(N__30220));
    LocalMux I__7028 (
            .O(N__30231),
            .I(N__30220));
    InMux I__7027 (
            .O(N__30230),
            .I(N__30217));
    Odrv4 I__7026 (
            .O(N__30225),
            .I(\c0.data_in_field_108 ));
    Odrv4 I__7025 (
            .O(N__30220),
            .I(\c0.data_in_field_108 ));
    LocalMux I__7024 (
            .O(N__30217),
            .I(\c0.data_in_field_108 ));
    InMux I__7023 (
            .O(N__30210),
            .I(N__30201));
    CascadeMux I__7022 (
            .O(N__30209),
            .I(N__30195));
    CascadeMux I__7021 (
            .O(N__30208),
            .I(N__30190));
    CascadeMux I__7020 (
            .O(N__30207),
            .I(N__30187));
    CascadeMux I__7019 (
            .O(N__30206),
            .I(N__30181));
    CascadeMux I__7018 (
            .O(N__30205),
            .I(N__30177));
    CascadeMux I__7017 (
            .O(N__30204),
            .I(N__30167));
    LocalMux I__7016 (
            .O(N__30201),
            .I(N__30164));
    InMux I__7015 (
            .O(N__30200),
            .I(N__30161));
    InMux I__7014 (
            .O(N__30199),
            .I(N__30154));
    InMux I__7013 (
            .O(N__30198),
            .I(N__30154));
    InMux I__7012 (
            .O(N__30195),
            .I(N__30154));
    CascadeMux I__7011 (
            .O(N__30194),
            .I(N__30150));
    CascadeMux I__7010 (
            .O(N__30193),
            .I(N__30141));
    InMux I__7009 (
            .O(N__30190),
            .I(N__30136));
    InMux I__7008 (
            .O(N__30187),
            .I(N__30136));
    InMux I__7007 (
            .O(N__30186),
            .I(N__30133));
    CascadeMux I__7006 (
            .O(N__30185),
            .I(N__30129));
    CascadeMux I__7005 (
            .O(N__30184),
            .I(N__30122));
    InMux I__7004 (
            .O(N__30181),
            .I(N__30114));
    InMux I__7003 (
            .O(N__30180),
            .I(N__30114));
    InMux I__7002 (
            .O(N__30177),
            .I(N__30114));
    CascadeMux I__7001 (
            .O(N__30176),
            .I(N__30106));
    CascadeMux I__7000 (
            .O(N__30175),
            .I(N__30102));
    CascadeMux I__6999 (
            .O(N__30174),
            .I(N__30097));
    CascadeMux I__6998 (
            .O(N__30173),
            .I(N__30094));
    InMux I__6997 (
            .O(N__30172),
            .I(N__30090));
    CascadeMux I__6996 (
            .O(N__30171),
            .I(N__30086));
    InMux I__6995 (
            .O(N__30170),
            .I(N__30081));
    InMux I__6994 (
            .O(N__30167),
            .I(N__30081));
    Span4Mux_v I__6993 (
            .O(N__30164),
            .I(N__30074));
    LocalMux I__6992 (
            .O(N__30161),
            .I(N__30074));
    LocalMux I__6991 (
            .O(N__30154),
            .I(N__30074));
    CascadeMux I__6990 (
            .O(N__30153),
            .I(N__30071));
    InMux I__6989 (
            .O(N__30150),
            .I(N__30066));
    CascadeMux I__6988 (
            .O(N__30149),
            .I(N__30062));
    CascadeMux I__6987 (
            .O(N__30148),
            .I(N__30056));
    InMux I__6986 (
            .O(N__30147),
            .I(N__30050));
    InMux I__6985 (
            .O(N__30146),
            .I(N__30047));
    InMux I__6984 (
            .O(N__30145),
            .I(N__30040));
    InMux I__6983 (
            .O(N__30144),
            .I(N__30040));
    InMux I__6982 (
            .O(N__30141),
            .I(N__30040));
    LocalMux I__6981 (
            .O(N__30136),
            .I(N__30035));
    LocalMux I__6980 (
            .O(N__30133),
            .I(N__30035));
    InMux I__6979 (
            .O(N__30132),
            .I(N__30030));
    InMux I__6978 (
            .O(N__30129),
            .I(N__30030));
    CascadeMux I__6977 (
            .O(N__30128),
            .I(N__30026));
    CascadeMux I__6976 (
            .O(N__30127),
            .I(N__30022));
    CascadeMux I__6975 (
            .O(N__30126),
            .I(N__30019));
    InMux I__6974 (
            .O(N__30125),
            .I(N__30009));
    InMux I__6973 (
            .O(N__30122),
            .I(N__30009));
    InMux I__6972 (
            .O(N__30121),
            .I(N__30009));
    LocalMux I__6971 (
            .O(N__30114),
            .I(N__30006));
    InMux I__6970 (
            .O(N__30113),
            .I(N__30003));
    CascadeMux I__6969 (
            .O(N__30112),
            .I(N__30000));
    InMux I__6968 (
            .O(N__30111),
            .I(N__29994));
    InMux I__6967 (
            .O(N__30110),
            .I(N__29994));
    InMux I__6966 (
            .O(N__30109),
            .I(N__29989));
    InMux I__6965 (
            .O(N__30106),
            .I(N__29989));
    InMux I__6964 (
            .O(N__30105),
            .I(N__29986));
    InMux I__6963 (
            .O(N__30102),
            .I(N__29981));
    InMux I__6962 (
            .O(N__30101),
            .I(N__29981));
    InMux I__6961 (
            .O(N__30100),
            .I(N__29978));
    InMux I__6960 (
            .O(N__30097),
            .I(N__29975));
    InMux I__6959 (
            .O(N__30094),
            .I(N__29972));
    CascadeMux I__6958 (
            .O(N__30093),
            .I(N__29967));
    LocalMux I__6957 (
            .O(N__30090),
            .I(N__29964));
    InMux I__6956 (
            .O(N__30089),
            .I(N__29959));
    InMux I__6955 (
            .O(N__30086),
            .I(N__29959));
    LocalMux I__6954 (
            .O(N__30081),
            .I(N__29956));
    Span4Mux_h I__6953 (
            .O(N__30074),
            .I(N__29953));
    InMux I__6952 (
            .O(N__30071),
            .I(N__29950));
    CascadeMux I__6951 (
            .O(N__30070),
            .I(N__29944));
    CascadeMux I__6950 (
            .O(N__30069),
            .I(N__29940));
    LocalMux I__6949 (
            .O(N__30066),
            .I(N__29935));
    InMux I__6948 (
            .O(N__30065),
            .I(N__29930));
    InMux I__6947 (
            .O(N__30062),
            .I(N__29930));
    CascadeMux I__6946 (
            .O(N__30061),
            .I(N__29926));
    CascadeMux I__6945 (
            .O(N__30060),
            .I(N__29921));
    CascadeMux I__6944 (
            .O(N__30059),
            .I(N__29918));
    InMux I__6943 (
            .O(N__30056),
            .I(N__29911));
    InMux I__6942 (
            .O(N__30055),
            .I(N__29911));
    InMux I__6941 (
            .O(N__30054),
            .I(N__29911));
    InMux I__6940 (
            .O(N__30053),
            .I(N__29908));
    LocalMux I__6939 (
            .O(N__30050),
            .I(N__29897));
    LocalMux I__6938 (
            .O(N__30047),
            .I(N__29897));
    LocalMux I__6937 (
            .O(N__30040),
            .I(N__29897));
    Span4Mux_h I__6936 (
            .O(N__30035),
            .I(N__29897));
    LocalMux I__6935 (
            .O(N__30030),
            .I(N__29897));
    InMux I__6934 (
            .O(N__30029),
            .I(N__29892));
    InMux I__6933 (
            .O(N__30026),
            .I(N__29892));
    InMux I__6932 (
            .O(N__30025),
            .I(N__29883));
    InMux I__6931 (
            .O(N__30022),
            .I(N__29883));
    InMux I__6930 (
            .O(N__30019),
            .I(N__29883));
    InMux I__6929 (
            .O(N__30018),
            .I(N__29883));
    InMux I__6928 (
            .O(N__30017),
            .I(N__29878));
    InMux I__6927 (
            .O(N__30016),
            .I(N__29878));
    LocalMux I__6926 (
            .O(N__30009),
            .I(N__29875));
    Span4Mux_v I__6925 (
            .O(N__30006),
            .I(N__29870));
    LocalMux I__6924 (
            .O(N__30003),
            .I(N__29870));
    InMux I__6923 (
            .O(N__30000),
            .I(N__29867));
    InMux I__6922 (
            .O(N__29999),
            .I(N__29864));
    LocalMux I__6921 (
            .O(N__29994),
            .I(N__29857));
    LocalMux I__6920 (
            .O(N__29989),
            .I(N__29857));
    LocalMux I__6919 (
            .O(N__29986),
            .I(N__29857));
    LocalMux I__6918 (
            .O(N__29981),
            .I(N__29854));
    LocalMux I__6917 (
            .O(N__29978),
            .I(N__29847));
    LocalMux I__6916 (
            .O(N__29975),
            .I(N__29847));
    LocalMux I__6915 (
            .O(N__29972),
            .I(N__29847));
    InMux I__6914 (
            .O(N__29971),
            .I(N__29842));
    InMux I__6913 (
            .O(N__29970),
            .I(N__29842));
    InMux I__6912 (
            .O(N__29967),
            .I(N__29839));
    Span4Mux_v I__6911 (
            .O(N__29964),
            .I(N__29828));
    LocalMux I__6910 (
            .O(N__29959),
            .I(N__29828));
    Span4Mux_v I__6909 (
            .O(N__29956),
            .I(N__29828));
    Span4Mux_h I__6908 (
            .O(N__29953),
            .I(N__29828));
    LocalMux I__6907 (
            .O(N__29950),
            .I(N__29828));
    InMux I__6906 (
            .O(N__29949),
            .I(N__29818));
    InMux I__6905 (
            .O(N__29948),
            .I(N__29818));
    InMux I__6904 (
            .O(N__29947),
            .I(N__29813));
    InMux I__6903 (
            .O(N__29944),
            .I(N__29813));
    InMux I__6902 (
            .O(N__29943),
            .I(N__29810));
    InMux I__6901 (
            .O(N__29940),
            .I(N__29807));
    InMux I__6900 (
            .O(N__29939),
            .I(N__29804));
    CascadeMux I__6899 (
            .O(N__29938),
            .I(N__29799));
    Span4Mux_h I__6898 (
            .O(N__29935),
            .I(N__29796));
    LocalMux I__6897 (
            .O(N__29930),
            .I(N__29793));
    InMux I__6896 (
            .O(N__29929),
            .I(N__29787));
    InMux I__6895 (
            .O(N__29926),
            .I(N__29787));
    CascadeMux I__6894 (
            .O(N__29925),
            .I(N__29783));
    CascadeMux I__6893 (
            .O(N__29924),
            .I(N__29779));
    InMux I__6892 (
            .O(N__29921),
            .I(N__29776));
    InMux I__6891 (
            .O(N__29918),
            .I(N__29773));
    LocalMux I__6890 (
            .O(N__29911),
            .I(N__29770));
    LocalMux I__6889 (
            .O(N__29908),
            .I(N__29765));
    Span4Mux_v I__6888 (
            .O(N__29897),
            .I(N__29765));
    LocalMux I__6887 (
            .O(N__29892),
            .I(N__29752));
    LocalMux I__6886 (
            .O(N__29883),
            .I(N__29752));
    LocalMux I__6885 (
            .O(N__29878),
            .I(N__29752));
    Span4Mux_v I__6884 (
            .O(N__29875),
            .I(N__29752));
    Span4Mux_h I__6883 (
            .O(N__29870),
            .I(N__29752));
    LocalMux I__6882 (
            .O(N__29867),
            .I(N__29752));
    LocalMux I__6881 (
            .O(N__29864),
            .I(N__29745));
    Span4Mux_v I__6880 (
            .O(N__29857),
            .I(N__29745));
    Span4Mux_v I__6879 (
            .O(N__29854),
            .I(N__29745));
    Span4Mux_v I__6878 (
            .O(N__29847),
            .I(N__29742));
    LocalMux I__6877 (
            .O(N__29842),
            .I(N__29735));
    LocalMux I__6876 (
            .O(N__29839),
            .I(N__29735));
    Span4Mux_v I__6875 (
            .O(N__29828),
            .I(N__29735));
    InMux I__6874 (
            .O(N__29827),
            .I(N__29732));
    InMux I__6873 (
            .O(N__29826),
            .I(N__29723));
    InMux I__6872 (
            .O(N__29825),
            .I(N__29723));
    InMux I__6871 (
            .O(N__29824),
            .I(N__29723));
    InMux I__6870 (
            .O(N__29823),
            .I(N__29723));
    LocalMux I__6869 (
            .O(N__29818),
            .I(N__29718));
    LocalMux I__6868 (
            .O(N__29813),
            .I(N__29718));
    LocalMux I__6867 (
            .O(N__29810),
            .I(N__29713));
    LocalMux I__6866 (
            .O(N__29807),
            .I(N__29713));
    LocalMux I__6865 (
            .O(N__29804),
            .I(N__29710));
    InMux I__6864 (
            .O(N__29803),
            .I(N__29703));
    InMux I__6863 (
            .O(N__29802),
            .I(N__29703));
    InMux I__6862 (
            .O(N__29799),
            .I(N__29703));
    Span4Mux_h I__6861 (
            .O(N__29796),
            .I(N__29698));
    Span4Mux_v I__6860 (
            .O(N__29793),
            .I(N__29698));
    InMux I__6859 (
            .O(N__29792),
            .I(N__29695));
    LocalMux I__6858 (
            .O(N__29787),
            .I(N__29692));
    InMux I__6857 (
            .O(N__29786),
            .I(N__29689));
    InMux I__6856 (
            .O(N__29783),
            .I(N__29686));
    InMux I__6855 (
            .O(N__29782),
            .I(N__29683));
    InMux I__6854 (
            .O(N__29779),
            .I(N__29680));
    LocalMux I__6853 (
            .O(N__29776),
            .I(N__29675));
    LocalMux I__6852 (
            .O(N__29773),
            .I(N__29675));
    Span4Mux_s2_h I__6851 (
            .O(N__29770),
            .I(N__29668));
    Span4Mux_v I__6850 (
            .O(N__29765),
            .I(N__29668));
    Span4Mux_h I__6849 (
            .O(N__29752),
            .I(N__29668));
    Span4Mux_v I__6848 (
            .O(N__29745),
            .I(N__29661));
    Span4Mux_h I__6847 (
            .O(N__29742),
            .I(N__29661));
    Span4Mux_v I__6846 (
            .O(N__29735),
            .I(N__29661));
    LocalMux I__6845 (
            .O(N__29732),
            .I(N__29646));
    LocalMux I__6844 (
            .O(N__29723),
            .I(N__29646));
    Span4Mux_s2_h I__6843 (
            .O(N__29718),
            .I(N__29646));
    Span4Mux_v I__6842 (
            .O(N__29713),
            .I(N__29646));
    Span4Mux_h I__6841 (
            .O(N__29710),
            .I(N__29646));
    LocalMux I__6840 (
            .O(N__29703),
            .I(N__29646));
    Span4Mux_h I__6839 (
            .O(N__29698),
            .I(N__29646));
    LocalMux I__6838 (
            .O(N__29695),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__6837 (
            .O(N__29692),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__6836 (
            .O(N__29689),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__6835 (
            .O(N__29686),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__6834 (
            .O(N__29683),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__6833 (
            .O(N__29680),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv12 I__6832 (
            .O(N__29675),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__6831 (
            .O(N__29668),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__6830 (
            .O(N__29661),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__6829 (
            .O(N__29646),
            .I(\c0.byte_transmit_counter2_1 ));
    CascadeMux I__6828 (
            .O(N__29625),
            .I(N__29622));
    InMux I__6827 (
            .O(N__29622),
            .I(N__29619));
    LocalMux I__6826 (
            .O(N__29619),
            .I(N__29616));
    Span4Mux_h I__6825 (
            .O(N__29616),
            .I(N__29613));
    Span4Mux_h I__6824 (
            .O(N__29613),
            .I(N__29609));
    InMux I__6823 (
            .O(N__29612),
            .I(N__29604));
    Span4Mux_h I__6822 (
            .O(N__29609),
            .I(N__29601));
    InMux I__6821 (
            .O(N__29608),
            .I(N__29598));
    InMux I__6820 (
            .O(N__29607),
            .I(N__29595));
    LocalMux I__6819 (
            .O(N__29604),
            .I(\c0.data_in_field_47 ));
    Odrv4 I__6818 (
            .O(N__29601),
            .I(\c0.data_in_field_47 ));
    LocalMux I__6817 (
            .O(N__29598),
            .I(\c0.data_in_field_47 ));
    LocalMux I__6816 (
            .O(N__29595),
            .I(\c0.data_in_field_47 ));
    InMux I__6815 (
            .O(N__29586),
            .I(N__29583));
    LocalMux I__6814 (
            .O(N__29583),
            .I(\c0.n5997 ));
    InMux I__6813 (
            .O(N__29580),
            .I(N__29577));
    LocalMux I__6812 (
            .O(N__29577),
            .I(N__29574));
    Span4Mux_v I__6811 (
            .O(N__29574),
            .I(N__29571));
    Span4Mux_h I__6810 (
            .O(N__29571),
            .I(N__29568));
    Span4Mux_h I__6809 (
            .O(N__29568),
            .I(N__29565));
    Odrv4 I__6808 (
            .O(N__29565),
            .I(\c0.n6000 ));
    InMux I__6807 (
            .O(N__29562),
            .I(N__29559));
    LocalMux I__6806 (
            .O(N__29559),
            .I(N__29555));
    InMux I__6805 (
            .O(N__29558),
            .I(N__29552));
    Span4Mux_v I__6804 (
            .O(N__29555),
            .I(N__29549));
    LocalMux I__6803 (
            .O(N__29552),
            .I(N__29546));
    Span4Mux_h I__6802 (
            .O(N__29549),
            .I(N__29543));
    Span4Mux_v I__6801 (
            .O(N__29546),
            .I(N__29539));
    Span4Mux_h I__6800 (
            .O(N__29543),
            .I(N__29536));
    InMux I__6799 (
            .O(N__29542),
            .I(N__29532));
    Span4Mux_h I__6798 (
            .O(N__29539),
            .I(N__29529));
    Span4Mux_v I__6797 (
            .O(N__29536),
            .I(N__29526));
    InMux I__6796 (
            .O(N__29535),
            .I(N__29523));
    LocalMux I__6795 (
            .O(N__29532),
            .I(\c0.data_in_field_84 ));
    Odrv4 I__6794 (
            .O(N__29529),
            .I(\c0.data_in_field_84 ));
    Odrv4 I__6793 (
            .O(N__29526),
            .I(\c0.data_in_field_84 ));
    LocalMux I__6792 (
            .O(N__29523),
            .I(\c0.data_in_field_84 ));
    InMux I__6791 (
            .O(N__29514),
            .I(N__29510));
    InMux I__6790 (
            .O(N__29513),
            .I(N__29507));
    LocalMux I__6789 (
            .O(N__29510),
            .I(N__29504));
    LocalMux I__6788 (
            .O(N__29507),
            .I(N__29500));
    Span4Mux_h I__6787 (
            .O(N__29504),
            .I(N__29497));
    InMux I__6786 (
            .O(N__29503),
            .I(N__29494));
    Sp12to4 I__6785 (
            .O(N__29500),
            .I(N__29491));
    Span4Mux_h I__6784 (
            .O(N__29497),
            .I(N__29488));
    LocalMux I__6783 (
            .O(N__29494),
            .I(N__29485));
    Span12Mux_v I__6782 (
            .O(N__29491),
            .I(N__29480));
    Span4Mux_h I__6781 (
            .O(N__29488),
            .I(N__29477));
    Span4Mux_h I__6780 (
            .O(N__29485),
            .I(N__29474));
    InMux I__6779 (
            .O(N__29484),
            .I(N__29469));
    InMux I__6778 (
            .O(N__29483),
            .I(N__29469));
    Odrv12 I__6777 (
            .O(N__29480),
            .I(\c0.data_in_field_70 ));
    Odrv4 I__6776 (
            .O(N__29477),
            .I(\c0.data_in_field_70 ));
    Odrv4 I__6775 (
            .O(N__29474),
            .I(\c0.data_in_field_70 ));
    LocalMux I__6774 (
            .O(N__29469),
            .I(\c0.data_in_field_70 ));
    InMux I__6773 (
            .O(N__29460),
            .I(N__29455));
    InMux I__6772 (
            .O(N__29459),
            .I(N__29450));
    InMux I__6771 (
            .O(N__29458),
            .I(N__29450));
    LocalMux I__6770 (
            .O(N__29455),
            .I(\c0.data_in_field_56 ));
    LocalMux I__6769 (
            .O(N__29450),
            .I(\c0.data_in_field_56 ));
    InMux I__6768 (
            .O(N__29445),
            .I(N__29442));
    LocalMux I__6767 (
            .O(N__29442),
            .I(N__29439));
    Span4Mux_h I__6766 (
            .O(N__29439),
            .I(N__29436));
    Odrv4 I__6765 (
            .O(N__29436),
            .I(\c0.n5494 ));
    InMux I__6764 (
            .O(N__29433),
            .I(N__29430));
    LocalMux I__6763 (
            .O(N__29430),
            .I(N__29426));
    InMux I__6762 (
            .O(N__29429),
            .I(N__29423));
    Span4Mux_s3_h I__6761 (
            .O(N__29426),
            .I(N__29420));
    LocalMux I__6760 (
            .O(N__29423),
            .I(N__29417));
    Odrv4 I__6759 (
            .O(N__29420),
            .I(\c0.n5554 ));
    Odrv12 I__6758 (
            .O(N__29417),
            .I(\c0.n5554 ));
    InMux I__6757 (
            .O(N__29412),
            .I(N__29409));
    LocalMux I__6756 (
            .O(N__29409),
            .I(N__29405));
    InMux I__6755 (
            .O(N__29408),
            .I(N__29402));
    Span4Mux_h I__6754 (
            .O(N__29405),
            .I(N__29399));
    LocalMux I__6753 (
            .O(N__29402),
            .I(N__29396));
    Span4Mux_v I__6752 (
            .O(N__29399),
            .I(N__29393));
    Span4Mux_v I__6751 (
            .O(N__29396),
            .I(N__29388));
    Span4Mux_h I__6750 (
            .O(N__29393),
            .I(N__29388));
    Odrv4 I__6749 (
            .O(N__29388),
            .I(\c0.n5524 ));
    CascadeMux I__6748 (
            .O(N__29385),
            .I(\c0.n5494_cascade_ ));
    InMux I__6747 (
            .O(N__29382),
            .I(N__29379));
    LocalMux I__6746 (
            .O(N__29379),
            .I(N__29375));
    InMux I__6745 (
            .O(N__29378),
            .I(N__29372));
    Span4Mux_v I__6744 (
            .O(N__29375),
            .I(N__29369));
    LocalMux I__6743 (
            .O(N__29372),
            .I(N__29366));
    Odrv4 I__6742 (
            .O(N__29369),
            .I(\c0.n5391 ));
    Odrv12 I__6741 (
            .O(N__29366),
            .I(\c0.n5391 ));
    InMux I__6740 (
            .O(N__29361),
            .I(N__29358));
    LocalMux I__6739 (
            .O(N__29358),
            .I(\c0.n26_adj_1927 ));
    InMux I__6738 (
            .O(N__29355),
            .I(N__29349));
    InMux I__6737 (
            .O(N__29354),
            .I(N__29349));
    LocalMux I__6736 (
            .O(N__29349),
            .I(r_Tx_Data_3));
    InMux I__6735 (
            .O(N__29346),
            .I(N__29342));
    InMux I__6734 (
            .O(N__29345),
            .I(N__29339));
    LocalMux I__6733 (
            .O(N__29342),
            .I(r_Tx_Data_2));
    LocalMux I__6732 (
            .O(N__29339),
            .I(r_Tx_Data_2));
    InMux I__6731 (
            .O(N__29334),
            .I(N__29328));
    InMux I__6730 (
            .O(N__29333),
            .I(N__29328));
    LocalMux I__6729 (
            .O(N__29328),
            .I(N__29322));
    InMux I__6728 (
            .O(N__29327),
            .I(N__29318));
    InMux I__6727 (
            .O(N__29326),
            .I(N__29312));
    InMux I__6726 (
            .O(N__29325),
            .I(N__29312));
    Span4Mux_h I__6725 (
            .O(N__29322),
            .I(N__29309));
    InMux I__6724 (
            .O(N__29321),
            .I(N__29306));
    LocalMux I__6723 (
            .O(N__29318),
            .I(N__29303));
    InMux I__6722 (
            .O(N__29317),
            .I(N__29300));
    LocalMux I__6721 (
            .O(N__29312),
            .I(N__29297));
    Odrv4 I__6720 (
            .O(N__29309),
            .I(\c0.tx.r_Bit_Index_0 ));
    LocalMux I__6719 (
            .O(N__29306),
            .I(\c0.tx.r_Bit_Index_0 ));
    Odrv12 I__6718 (
            .O(N__29303),
            .I(\c0.tx.r_Bit_Index_0 ));
    LocalMux I__6717 (
            .O(N__29300),
            .I(\c0.tx.r_Bit_Index_0 ));
    Odrv4 I__6716 (
            .O(N__29297),
            .I(\c0.tx.r_Bit_Index_0 ));
    InMux I__6715 (
            .O(N__29286),
            .I(N__29283));
    LocalMux I__6714 (
            .O(N__29283),
            .I(N__29279));
    InMux I__6713 (
            .O(N__29282),
            .I(N__29276));
    Span4Mux_h I__6712 (
            .O(N__29279),
            .I(N__29273));
    LocalMux I__6711 (
            .O(N__29276),
            .I(\c0.tx.r_Tx_Data_0 ));
    Odrv4 I__6710 (
            .O(N__29273),
            .I(\c0.tx.r_Tx_Data_0 ));
    CascadeMux I__6709 (
            .O(N__29268),
            .I(\c0.tx.n6051_cascade_ ));
    InMux I__6708 (
            .O(N__29265),
            .I(N__29261));
    InMux I__6707 (
            .O(N__29264),
            .I(N__29258));
    LocalMux I__6706 (
            .O(N__29261),
            .I(r_Tx_Data_1));
    LocalMux I__6705 (
            .O(N__29258),
            .I(r_Tx_Data_1));
    CascadeMux I__6704 (
            .O(N__29253),
            .I(N__29249));
    InMux I__6703 (
            .O(N__29252),
            .I(N__29246));
    InMux I__6702 (
            .O(N__29249),
            .I(N__29243));
    LocalMux I__6701 (
            .O(N__29246),
            .I(N__29240));
    LocalMux I__6700 (
            .O(N__29243),
            .I(N__29235));
    Span4Mux_h I__6699 (
            .O(N__29240),
            .I(N__29232));
    InMux I__6698 (
            .O(N__29239),
            .I(N__29229));
    InMux I__6697 (
            .O(N__29238),
            .I(N__29226));
    Span4Mux_v I__6696 (
            .O(N__29235),
            .I(N__29223));
    Span4Mux_h I__6695 (
            .O(N__29232),
            .I(N__29220));
    LocalMux I__6694 (
            .O(N__29229),
            .I(\c0.tx.r_Bit_Index_2 ));
    LocalMux I__6693 (
            .O(N__29226),
            .I(\c0.tx.r_Bit_Index_2 ));
    Odrv4 I__6692 (
            .O(N__29223),
            .I(\c0.tx.r_Bit_Index_2 ));
    Odrv4 I__6691 (
            .O(N__29220),
            .I(\c0.tx.r_Bit_Index_2 ));
    InMux I__6690 (
            .O(N__29211),
            .I(N__29208));
    LocalMux I__6689 (
            .O(N__29208),
            .I(\c0.tx.n6054 ));
    InMux I__6688 (
            .O(N__29205),
            .I(N__29193));
    InMux I__6687 (
            .O(N__29204),
            .I(N__29193));
    InMux I__6686 (
            .O(N__29203),
            .I(N__29190));
    InMux I__6685 (
            .O(N__29202),
            .I(N__29185));
    InMux I__6684 (
            .O(N__29201),
            .I(N__29185));
    InMux I__6683 (
            .O(N__29200),
            .I(N__29182));
    InMux I__6682 (
            .O(N__29199),
            .I(N__29179));
    InMux I__6681 (
            .O(N__29198),
            .I(N__29176));
    LocalMux I__6680 (
            .O(N__29193),
            .I(N__29170));
    LocalMux I__6679 (
            .O(N__29190),
            .I(N__29167));
    LocalMux I__6678 (
            .O(N__29185),
            .I(N__29164));
    LocalMux I__6677 (
            .O(N__29182),
            .I(N__29161));
    LocalMux I__6676 (
            .O(N__29179),
            .I(N__29156));
    LocalMux I__6675 (
            .O(N__29176),
            .I(N__29156));
    InMux I__6674 (
            .O(N__29175),
            .I(N__29153));
    InMux I__6673 (
            .O(N__29174),
            .I(N__29150));
    InMux I__6672 (
            .O(N__29173),
            .I(N__29147));
    Span4Mux_v I__6671 (
            .O(N__29170),
            .I(N__29138));
    Span4Mux_v I__6670 (
            .O(N__29167),
            .I(N__29138));
    Span4Mux_v I__6669 (
            .O(N__29164),
            .I(N__29138));
    Span4Mux_h I__6668 (
            .O(N__29161),
            .I(N__29138));
    Span4Mux_h I__6667 (
            .O(N__29156),
            .I(N__29135));
    LocalMux I__6666 (
            .O(N__29153),
            .I(r_SM_Main_0));
    LocalMux I__6665 (
            .O(N__29150),
            .I(r_SM_Main_0));
    LocalMux I__6664 (
            .O(N__29147),
            .I(r_SM_Main_0));
    Odrv4 I__6663 (
            .O(N__29138),
            .I(r_SM_Main_0));
    Odrv4 I__6662 (
            .O(N__29135),
            .I(r_SM_Main_0));
    CascadeMux I__6661 (
            .O(N__29124),
            .I(\c0.tx.o_Tx_Serial_N_1798_cascade_ ));
    InMux I__6660 (
            .O(N__29121),
            .I(N__29118));
    LocalMux I__6659 (
            .O(N__29118),
            .I(N__29109));
    InMux I__6658 (
            .O(N__29117),
            .I(N__29106));
    InMux I__6657 (
            .O(N__29116),
            .I(N__29101));
    InMux I__6656 (
            .O(N__29115),
            .I(N__29101));
    InMux I__6655 (
            .O(N__29114),
            .I(N__29098));
    InMux I__6654 (
            .O(N__29113),
            .I(N__29093));
    InMux I__6653 (
            .O(N__29112),
            .I(N__29093));
    Span4Mux_h I__6652 (
            .O(N__29109),
            .I(N__29082));
    LocalMux I__6651 (
            .O(N__29106),
            .I(N__29082));
    LocalMux I__6650 (
            .O(N__29101),
            .I(N__29079));
    LocalMux I__6649 (
            .O(N__29098),
            .I(N__29074));
    LocalMux I__6648 (
            .O(N__29093),
            .I(N__29074));
    InMux I__6647 (
            .O(N__29092),
            .I(N__29071));
    InMux I__6646 (
            .O(N__29091),
            .I(N__29067));
    InMux I__6645 (
            .O(N__29090),
            .I(N__29064));
    InMux I__6644 (
            .O(N__29089),
            .I(N__29061));
    InMux I__6643 (
            .O(N__29088),
            .I(N__29056));
    InMux I__6642 (
            .O(N__29087),
            .I(N__29056));
    Span4Mux_h I__6641 (
            .O(N__29082),
            .I(N__29053));
    Span4Mux_h I__6640 (
            .O(N__29079),
            .I(N__29050));
    Span4Mux_h I__6639 (
            .O(N__29074),
            .I(N__29045));
    LocalMux I__6638 (
            .O(N__29071),
            .I(N__29045));
    InMux I__6637 (
            .O(N__29070),
            .I(N__29042));
    LocalMux I__6636 (
            .O(N__29067),
            .I(r_SM_Main_1));
    LocalMux I__6635 (
            .O(N__29064),
            .I(r_SM_Main_1));
    LocalMux I__6634 (
            .O(N__29061),
            .I(r_SM_Main_1));
    LocalMux I__6633 (
            .O(N__29056),
            .I(r_SM_Main_1));
    Odrv4 I__6632 (
            .O(N__29053),
            .I(r_SM_Main_1));
    Odrv4 I__6631 (
            .O(N__29050),
            .I(r_SM_Main_1));
    Odrv4 I__6630 (
            .O(N__29045),
            .I(r_SM_Main_1));
    LocalMux I__6629 (
            .O(N__29042),
            .I(r_SM_Main_1));
    CascadeMux I__6628 (
            .O(N__29025),
            .I(\c0.tx.n12_cascade_ ));
    CascadeMux I__6627 (
            .O(N__29022),
            .I(N__29018));
    CascadeMux I__6626 (
            .O(N__29021),
            .I(N__29012));
    InMux I__6625 (
            .O(N__29018),
            .I(N__29006));
    InMux I__6624 (
            .O(N__29017),
            .I(N__29001));
    InMux I__6623 (
            .O(N__29016),
            .I(N__28998));
    InMux I__6622 (
            .O(N__29015),
            .I(N__28993));
    InMux I__6621 (
            .O(N__29012),
            .I(N__28993));
    InMux I__6620 (
            .O(N__29011),
            .I(N__28986));
    InMux I__6619 (
            .O(N__29010),
            .I(N__28986));
    InMux I__6618 (
            .O(N__29009),
            .I(N__28986));
    LocalMux I__6617 (
            .O(N__29006),
            .I(N__28983));
    InMux I__6616 (
            .O(N__29005),
            .I(N__28980));
    CascadeMux I__6615 (
            .O(N__29004),
            .I(N__28970));
    LocalMux I__6614 (
            .O(N__29001),
            .I(N__28965));
    LocalMux I__6613 (
            .O(N__28998),
            .I(N__28962));
    LocalMux I__6612 (
            .O(N__28993),
            .I(N__28959));
    LocalMux I__6611 (
            .O(N__28986),
            .I(N__28949));
    Span4Mux_v I__6610 (
            .O(N__28983),
            .I(N__28949));
    LocalMux I__6609 (
            .O(N__28980),
            .I(N__28949));
    InMux I__6608 (
            .O(N__28979),
            .I(N__28946));
    InMux I__6607 (
            .O(N__28978),
            .I(N__28937));
    InMux I__6606 (
            .O(N__28977),
            .I(N__28937));
    InMux I__6605 (
            .O(N__28976),
            .I(N__28937));
    InMux I__6604 (
            .O(N__28975),
            .I(N__28937));
    InMux I__6603 (
            .O(N__28974),
            .I(N__28934));
    InMux I__6602 (
            .O(N__28973),
            .I(N__28925));
    InMux I__6601 (
            .O(N__28970),
            .I(N__28925));
    InMux I__6600 (
            .O(N__28969),
            .I(N__28925));
    InMux I__6599 (
            .O(N__28968),
            .I(N__28925));
    Span4Mux_h I__6598 (
            .O(N__28965),
            .I(N__28922));
    Span4Mux_h I__6597 (
            .O(N__28962),
            .I(N__28917));
    Span4Mux_v I__6596 (
            .O(N__28959),
            .I(N__28917));
    InMux I__6595 (
            .O(N__28958),
            .I(N__28910));
    InMux I__6594 (
            .O(N__28957),
            .I(N__28910));
    InMux I__6593 (
            .O(N__28956),
            .I(N__28910));
    Span4Mux_h I__6592 (
            .O(N__28949),
            .I(N__28907));
    LocalMux I__6591 (
            .O(N__28946),
            .I(r_SM_Main_2));
    LocalMux I__6590 (
            .O(N__28937),
            .I(r_SM_Main_2));
    LocalMux I__6589 (
            .O(N__28934),
            .I(r_SM_Main_2));
    LocalMux I__6588 (
            .O(N__28925),
            .I(r_SM_Main_2));
    Odrv4 I__6587 (
            .O(N__28922),
            .I(r_SM_Main_2));
    Odrv4 I__6586 (
            .O(N__28917),
            .I(r_SM_Main_2));
    LocalMux I__6585 (
            .O(N__28910),
            .I(r_SM_Main_2));
    Odrv4 I__6584 (
            .O(N__28907),
            .I(r_SM_Main_2));
    IoInMux I__6583 (
            .O(N__28890),
            .I(N__28887));
    LocalMux I__6582 (
            .O(N__28887),
            .I(N__28884));
    IoSpan4Mux I__6581 (
            .O(N__28884),
            .I(N__28880));
    InMux I__6580 (
            .O(N__28883),
            .I(N__28877));
    Span4Mux_s0_v I__6579 (
            .O(N__28880),
            .I(N__28872));
    LocalMux I__6578 (
            .O(N__28877),
            .I(N__28872));
    Span4Mux_v I__6577 (
            .O(N__28872),
            .I(N__28869));
    Span4Mux_h I__6576 (
            .O(N__28869),
            .I(N__28865));
    InMux I__6575 (
            .O(N__28868),
            .I(N__28862));
    Odrv4 I__6574 (
            .O(N__28865),
            .I(tx_o));
    LocalMux I__6573 (
            .O(N__28862),
            .I(tx_o));
    CascadeMux I__6572 (
            .O(N__28857),
            .I(N__28854));
    InMux I__6571 (
            .O(N__28854),
            .I(N__28851));
    LocalMux I__6570 (
            .O(N__28851),
            .I(N__28848));
    Span4Mux_h I__6569 (
            .O(N__28848),
            .I(N__28845));
    Span4Mux_h I__6568 (
            .O(N__28845),
            .I(N__28842));
    Span4Mux_v I__6567 (
            .O(N__28842),
            .I(N__28837));
    InMux I__6566 (
            .O(N__28841),
            .I(N__28834));
    InMux I__6565 (
            .O(N__28840),
            .I(N__28831));
    Odrv4 I__6564 (
            .O(N__28837),
            .I(data_in_10_5));
    LocalMux I__6563 (
            .O(N__28834),
            .I(data_in_10_5));
    LocalMux I__6562 (
            .O(N__28831),
            .I(data_in_10_5));
    CascadeMux I__6561 (
            .O(N__28824),
            .I(N__28821));
    InMux I__6560 (
            .O(N__28821),
            .I(N__28818));
    LocalMux I__6559 (
            .O(N__28818),
            .I(N__28813));
    InMux I__6558 (
            .O(N__28817),
            .I(N__28810));
    InMux I__6557 (
            .O(N__28816),
            .I(N__28807));
    Odrv12 I__6556 (
            .O(N__28813),
            .I(data_in_9_5));
    LocalMux I__6555 (
            .O(N__28810),
            .I(data_in_9_5));
    LocalMux I__6554 (
            .O(N__28807),
            .I(data_in_9_5));
    InMux I__6553 (
            .O(N__28800),
            .I(N__28796));
    InMux I__6552 (
            .O(N__28799),
            .I(N__28793));
    LocalMux I__6551 (
            .O(N__28796),
            .I(N__28790));
    LocalMux I__6550 (
            .O(N__28793),
            .I(N__28787));
    Span4Mux_v I__6549 (
            .O(N__28790),
            .I(N__28782));
    Span4Mux_v I__6548 (
            .O(N__28787),
            .I(N__28782));
    Span4Mux_h I__6547 (
            .O(N__28782),
            .I(N__28778));
    InMux I__6546 (
            .O(N__28781),
            .I(N__28775));
    Odrv4 I__6545 (
            .O(N__28778),
            .I(data_in_6_0));
    LocalMux I__6544 (
            .O(N__28775),
            .I(data_in_6_0));
    CascadeMux I__6543 (
            .O(N__28770),
            .I(N__28767));
    InMux I__6542 (
            .O(N__28767),
            .I(N__28764));
    LocalMux I__6541 (
            .O(N__28764),
            .I(N__28761));
    Odrv4 I__6540 (
            .O(N__28761),
            .I(\c0.n9 ));
    InMux I__6539 (
            .O(N__28758),
            .I(N__28755));
    LocalMux I__6538 (
            .O(N__28755),
            .I(N__28752));
    Span4Mux_h I__6537 (
            .O(N__28752),
            .I(N__28749));
    Odrv4 I__6536 (
            .O(N__28749),
            .I(n8_adj_1987));
    InMux I__6535 (
            .O(N__28746),
            .I(N__28740));
    InMux I__6534 (
            .O(N__28745),
            .I(N__28740));
    LocalMux I__6533 (
            .O(N__28740),
            .I(N__28737));
    Odrv4 I__6532 (
            .O(N__28737),
            .I(n5400));
    InMux I__6531 (
            .O(N__28734),
            .I(N__28731));
    LocalMux I__6530 (
            .O(N__28731),
            .I(N__28728));
    Odrv4 I__6529 (
            .O(N__28728),
            .I(tx_data_2_N_keep));
    InMux I__6528 (
            .O(N__28725),
            .I(N__28722));
    LocalMux I__6527 (
            .O(N__28722),
            .I(N__28719));
    Span4Mux_h I__6526 (
            .O(N__28719),
            .I(N__28716));
    Odrv4 I__6525 (
            .O(N__28716),
            .I(n5364));
    CascadeMux I__6524 (
            .O(N__28713),
            .I(N__28710));
    InMux I__6523 (
            .O(N__28710),
            .I(N__28706));
    InMux I__6522 (
            .O(N__28709),
            .I(N__28703));
    LocalMux I__6521 (
            .O(N__28706),
            .I(N__28700));
    LocalMux I__6520 (
            .O(N__28703),
            .I(N__28697));
    Odrv12 I__6519 (
            .O(N__28700),
            .I(n5482));
    Odrv4 I__6518 (
            .O(N__28697),
            .I(n5482));
    InMux I__6517 (
            .O(N__28692),
            .I(N__28689));
    LocalMux I__6516 (
            .O(N__28689),
            .I(N__28685));
    InMux I__6515 (
            .O(N__28688),
            .I(N__28682));
    Odrv4 I__6514 (
            .O(N__28685),
            .I(n1768));
    LocalMux I__6513 (
            .O(N__28682),
            .I(n1768));
    CascadeMux I__6512 (
            .O(N__28677),
            .I(n5364_cascade_));
    CascadeMux I__6511 (
            .O(N__28674),
            .I(N__28671));
    InMux I__6510 (
            .O(N__28671),
            .I(N__28668));
    LocalMux I__6509 (
            .O(N__28668),
            .I(n5871));
    InMux I__6508 (
            .O(N__28665),
            .I(N__28662));
    LocalMux I__6507 (
            .O(N__28662),
            .I(\c0.n6312 ));
    CascadeMux I__6506 (
            .O(N__28659),
            .I(N__28656));
    InMux I__6505 (
            .O(N__28656),
            .I(N__28653));
    LocalMux I__6504 (
            .O(N__28653),
            .I(tx_data_3_N_keep));
    CascadeMux I__6503 (
            .O(N__28650),
            .I(N__28647));
    InMux I__6502 (
            .O(N__28647),
            .I(N__28644));
    LocalMux I__6501 (
            .O(N__28644),
            .I(\c0.n5853 ));
    InMux I__6500 (
            .O(N__28641),
            .I(N__28629));
    InMux I__6499 (
            .O(N__28640),
            .I(N__28629));
    InMux I__6498 (
            .O(N__28639),
            .I(N__28629));
    InMux I__6497 (
            .O(N__28638),
            .I(N__28622));
    InMux I__6496 (
            .O(N__28637),
            .I(N__28622));
    InMux I__6495 (
            .O(N__28636),
            .I(N__28622));
    LocalMux I__6494 (
            .O(N__28629),
            .I(tx_active));
    LocalMux I__6493 (
            .O(N__28622),
            .I(tx_active));
    CascadeMux I__6492 (
            .O(N__28617),
            .I(N__28614));
    InMux I__6491 (
            .O(N__28614),
            .I(N__28610));
    InMux I__6490 (
            .O(N__28613),
            .I(N__28605));
    LocalMux I__6489 (
            .O(N__28610),
            .I(N__28602));
    InMux I__6488 (
            .O(N__28609),
            .I(N__28599));
    CascadeMux I__6487 (
            .O(N__28608),
            .I(N__28594));
    LocalMux I__6486 (
            .O(N__28605),
            .I(N__28587));
    Span4Mux_h I__6485 (
            .O(N__28602),
            .I(N__28587));
    LocalMux I__6484 (
            .O(N__28599),
            .I(N__28587));
    CascadeMux I__6483 (
            .O(N__28598),
            .I(N__28584));
    CascadeMux I__6482 (
            .O(N__28597),
            .I(N__28580));
    InMux I__6481 (
            .O(N__28594),
            .I(N__28577));
    Span4Mux_v I__6480 (
            .O(N__28587),
            .I(N__28574));
    InMux I__6479 (
            .O(N__28584),
            .I(N__28567));
    InMux I__6478 (
            .O(N__28583),
            .I(N__28567));
    InMux I__6477 (
            .O(N__28580),
            .I(N__28567));
    LocalMux I__6476 (
            .O(N__28577),
            .I(\c0.tx_transmit ));
    Odrv4 I__6475 (
            .O(N__28574),
            .I(\c0.tx_transmit ));
    LocalMux I__6474 (
            .O(N__28567),
            .I(\c0.tx_transmit ));
    InMux I__6473 (
            .O(N__28560),
            .I(N__28557));
    LocalMux I__6472 (
            .O(N__28557),
            .I(N__28554));
    Odrv4 I__6471 (
            .O(N__28554),
            .I(n135));
    CascadeMux I__6470 (
            .O(N__28551),
            .I(n4_adj_1986_cascade_));
    InMux I__6469 (
            .O(N__28548),
            .I(N__28544));
    InMux I__6468 (
            .O(N__28547),
            .I(N__28541));
    LocalMux I__6467 (
            .O(N__28544),
            .I(N__28538));
    LocalMux I__6466 (
            .O(N__28541),
            .I(data_out_19_6));
    Odrv12 I__6465 (
            .O(N__28538),
            .I(data_out_19_6));
    CascadeMux I__6464 (
            .O(N__28533),
            .I(N__28529));
    InMux I__6463 (
            .O(N__28532),
            .I(N__28526));
    InMux I__6462 (
            .O(N__28529),
            .I(N__28523));
    LocalMux I__6461 (
            .O(N__28526),
            .I(data_out_19_5));
    LocalMux I__6460 (
            .O(N__28523),
            .I(data_out_19_5));
    CascadeMux I__6459 (
            .O(N__28518),
            .I(N__28514));
    InMux I__6458 (
            .O(N__28517),
            .I(N__28509));
    InMux I__6457 (
            .O(N__28514),
            .I(N__28509));
    LocalMux I__6456 (
            .O(N__28509),
            .I(n5440));
    CascadeMux I__6455 (
            .O(N__28506),
            .I(n5_cascade_));
    InMux I__6454 (
            .O(N__28503),
            .I(N__28500));
    LocalMux I__6453 (
            .O(N__28500),
            .I(\c0.tx_active_prev ));
    InMux I__6452 (
            .O(N__28497),
            .I(N__28490));
    InMux I__6451 (
            .O(N__28496),
            .I(N__28490));
    InMux I__6450 (
            .O(N__28495),
            .I(N__28487));
    LocalMux I__6449 (
            .O(N__28490),
            .I(N__28482));
    LocalMux I__6448 (
            .O(N__28487),
            .I(N__28479));
    InMux I__6447 (
            .O(N__28486),
            .I(N__28472));
    InMux I__6446 (
            .O(N__28485),
            .I(N__28472));
    Span4Mux_h I__6445 (
            .O(N__28482),
            .I(N__28469));
    Span4Mux_h I__6444 (
            .O(N__28479),
            .I(N__28466));
    InMux I__6443 (
            .O(N__28478),
            .I(N__28461));
    InMux I__6442 (
            .O(N__28477),
            .I(N__28461));
    LocalMux I__6441 (
            .O(N__28472),
            .I(\c0.tx.r_SM_Main_2_N_1767_1 ));
    Odrv4 I__6440 (
            .O(N__28469),
            .I(\c0.tx.r_SM_Main_2_N_1767_1 ));
    Odrv4 I__6439 (
            .O(N__28466),
            .I(\c0.tx.r_SM_Main_2_N_1767_1 ));
    LocalMux I__6438 (
            .O(N__28461),
            .I(\c0.tx.r_SM_Main_2_N_1767_1 ));
    InMux I__6437 (
            .O(N__28452),
            .I(N__28449));
    LocalMux I__6436 (
            .O(N__28449),
            .I(N__28446));
    Odrv4 I__6435 (
            .O(N__28446),
            .I(\c0.tx.n2177 ));
    CascadeMux I__6434 (
            .O(N__28443),
            .I(n4333_cascade_));
    CascadeMux I__6433 (
            .O(N__28440),
            .I(\c0.n81_adj_1872_cascade_ ));
    InMux I__6432 (
            .O(N__28437),
            .I(N__28434));
    LocalMux I__6431 (
            .O(N__28434),
            .I(N__28429));
    InMux I__6430 (
            .O(N__28433),
            .I(N__28426));
    InMux I__6429 (
            .O(N__28432),
            .I(N__28423));
    Span4Mux_v I__6428 (
            .O(N__28429),
            .I(N__28420));
    LocalMux I__6427 (
            .O(N__28426),
            .I(N__28416));
    LocalMux I__6426 (
            .O(N__28423),
            .I(N__28413));
    Span4Mux_h I__6425 (
            .O(N__28420),
            .I(N__28410));
    InMux I__6424 (
            .O(N__28419),
            .I(N__28407));
    Span4Mux_v I__6423 (
            .O(N__28416),
            .I(N__28402));
    Span4Mux_v I__6422 (
            .O(N__28413),
            .I(N__28402));
    Odrv4 I__6421 (
            .O(N__28410),
            .I(data_in_2_0));
    LocalMux I__6420 (
            .O(N__28407),
            .I(data_in_2_0));
    Odrv4 I__6419 (
            .O(N__28402),
            .I(data_in_2_0));
    CascadeMux I__6418 (
            .O(N__28395),
            .I(N__28392));
    InMux I__6417 (
            .O(N__28392),
            .I(N__28388));
    InMux I__6416 (
            .O(N__28391),
            .I(N__28385));
    LocalMux I__6415 (
            .O(N__28388),
            .I(N__28382));
    LocalMux I__6414 (
            .O(N__28385),
            .I(N__28379));
    Span4Mux_v I__6413 (
            .O(N__28382),
            .I(N__28376));
    Span4Mux_h I__6412 (
            .O(N__28379),
            .I(N__28373));
    Span4Mux_h I__6411 (
            .O(N__28376),
            .I(N__28368));
    Span4Mux_h I__6410 (
            .O(N__28373),
            .I(N__28368));
    Span4Mux_h I__6409 (
            .O(N__28368),
            .I(N__28364));
    InMux I__6408 (
            .O(N__28367),
            .I(N__28361));
    Odrv4 I__6407 (
            .O(N__28364),
            .I(data_in_13_2));
    LocalMux I__6406 (
            .O(N__28361),
            .I(data_in_13_2));
    InMux I__6405 (
            .O(N__28356),
            .I(N__28353));
    LocalMux I__6404 (
            .O(N__28353),
            .I(N__28350));
    Span4Mux_v I__6403 (
            .O(N__28350),
            .I(N__28345));
    InMux I__6402 (
            .O(N__28349),
            .I(N__28340));
    InMux I__6401 (
            .O(N__28348),
            .I(N__28340));
    Sp12to4 I__6400 (
            .O(N__28345),
            .I(N__28333));
    LocalMux I__6399 (
            .O(N__28340),
            .I(N__28333));
    InMux I__6398 (
            .O(N__28339),
            .I(N__28329));
    InMux I__6397 (
            .O(N__28338),
            .I(N__28326));
    Span12Mux_s10_h I__6396 (
            .O(N__28333),
            .I(N__28323));
    InMux I__6395 (
            .O(N__28332),
            .I(N__28320));
    LocalMux I__6394 (
            .O(N__28329),
            .I(\c0.data_in_field_88 ));
    LocalMux I__6393 (
            .O(N__28326),
            .I(\c0.data_in_field_88 ));
    Odrv12 I__6392 (
            .O(N__28323),
            .I(\c0.data_in_field_88 ));
    LocalMux I__6391 (
            .O(N__28320),
            .I(\c0.data_in_field_88 ));
    CascadeMux I__6390 (
            .O(N__28311),
            .I(N__28307));
    InMux I__6389 (
            .O(N__28310),
            .I(N__28303));
    InMux I__6388 (
            .O(N__28307),
            .I(N__28300));
    InMux I__6387 (
            .O(N__28306),
            .I(N__28296));
    LocalMux I__6386 (
            .O(N__28303),
            .I(N__28291));
    LocalMux I__6385 (
            .O(N__28300),
            .I(N__28291));
    InMux I__6384 (
            .O(N__28299),
            .I(N__28288));
    LocalMux I__6383 (
            .O(N__28296),
            .I(N__28285));
    Span4Mux_s3_h I__6382 (
            .O(N__28291),
            .I(N__28282));
    LocalMux I__6381 (
            .O(N__28288),
            .I(N__28278));
    Span4Mux_h I__6380 (
            .O(N__28285),
            .I(N__28274));
    Span4Mux_h I__6379 (
            .O(N__28282),
            .I(N__28271));
    InMux I__6378 (
            .O(N__28281),
            .I(N__28267));
    Span4Mux_h I__6377 (
            .O(N__28278),
            .I(N__28264));
    InMux I__6376 (
            .O(N__28277),
            .I(N__28261));
    Span4Mux_h I__6375 (
            .O(N__28274),
            .I(N__28258));
    Span4Mux_h I__6374 (
            .O(N__28271),
            .I(N__28255));
    InMux I__6373 (
            .O(N__28270),
            .I(N__28252));
    LocalMux I__6372 (
            .O(N__28267),
            .I(\c0.data_in_field_98 ));
    Odrv4 I__6371 (
            .O(N__28264),
            .I(\c0.data_in_field_98 ));
    LocalMux I__6370 (
            .O(N__28261),
            .I(\c0.data_in_field_98 ));
    Odrv4 I__6369 (
            .O(N__28258),
            .I(\c0.data_in_field_98 ));
    Odrv4 I__6368 (
            .O(N__28255),
            .I(\c0.data_in_field_98 ));
    LocalMux I__6367 (
            .O(N__28252),
            .I(\c0.data_in_field_98 ));
    InMux I__6366 (
            .O(N__28239),
            .I(N__28235));
    InMux I__6365 (
            .O(N__28238),
            .I(N__28231));
    LocalMux I__6364 (
            .O(N__28235),
            .I(N__28228));
    CascadeMux I__6363 (
            .O(N__28234),
            .I(N__28225));
    LocalMux I__6362 (
            .O(N__28231),
            .I(N__28221));
    Span4Mux_v I__6361 (
            .O(N__28228),
            .I(N__28218));
    InMux I__6360 (
            .O(N__28225),
            .I(N__28215));
    InMux I__6359 (
            .O(N__28224),
            .I(N__28212));
    Span4Mux_v I__6358 (
            .O(N__28221),
            .I(N__28209));
    Span4Mux_h I__6357 (
            .O(N__28218),
            .I(N__28204));
    LocalMux I__6356 (
            .O(N__28215),
            .I(N__28204));
    LocalMux I__6355 (
            .O(N__28212),
            .I(\c0.data_in_field_28 ));
    Odrv4 I__6354 (
            .O(N__28209),
            .I(\c0.data_in_field_28 ));
    Odrv4 I__6353 (
            .O(N__28204),
            .I(\c0.data_in_field_28 ));
    InMux I__6352 (
            .O(N__28197),
            .I(N__28192));
    InMux I__6351 (
            .O(N__28196),
            .I(N__28189));
    InMux I__6350 (
            .O(N__28195),
            .I(N__28185));
    LocalMux I__6349 (
            .O(N__28192),
            .I(N__28182));
    LocalMux I__6348 (
            .O(N__28189),
            .I(N__28179));
    InMux I__6347 (
            .O(N__28188),
            .I(N__28176));
    LocalMux I__6346 (
            .O(N__28185),
            .I(N__28173));
    Span4Mux_v I__6345 (
            .O(N__28182),
            .I(N__28170));
    Span4Mux_h I__6344 (
            .O(N__28179),
            .I(N__28165));
    LocalMux I__6343 (
            .O(N__28176),
            .I(N__28162));
    Span4Mux_v I__6342 (
            .O(N__28173),
            .I(N__28157));
    Span4Mux_h I__6341 (
            .O(N__28170),
            .I(N__28157));
    InMux I__6340 (
            .O(N__28169),
            .I(N__28152));
    InMux I__6339 (
            .O(N__28168),
            .I(N__28152));
    Odrv4 I__6338 (
            .O(N__28165),
            .I(\c0.data_in_field_121 ));
    Odrv4 I__6337 (
            .O(N__28162),
            .I(\c0.data_in_field_121 ));
    Odrv4 I__6336 (
            .O(N__28157),
            .I(\c0.data_in_field_121 ));
    LocalMux I__6335 (
            .O(N__28152),
            .I(\c0.data_in_field_121 ));
    CascadeMux I__6334 (
            .O(N__28143),
            .I(N__28140));
    InMux I__6333 (
            .O(N__28140),
            .I(N__28137));
    LocalMux I__6332 (
            .O(N__28137),
            .I(N__28134));
    Odrv4 I__6331 (
            .O(N__28134),
            .I(\c0.n23_adj_1935 ));
    InMux I__6330 (
            .O(N__28131),
            .I(N__28127));
    InMux I__6329 (
            .O(N__28130),
            .I(N__28123));
    LocalMux I__6328 (
            .O(N__28127),
            .I(N__28118));
    InMux I__6327 (
            .O(N__28126),
            .I(N__28115));
    LocalMux I__6326 (
            .O(N__28123),
            .I(N__28111));
    InMux I__6325 (
            .O(N__28122),
            .I(N__28108));
    CascadeMux I__6324 (
            .O(N__28121),
            .I(N__28105));
    Span4Mux_v I__6323 (
            .O(N__28118),
            .I(N__28100));
    LocalMux I__6322 (
            .O(N__28115),
            .I(N__28100));
    InMux I__6321 (
            .O(N__28114),
            .I(N__28097));
    Span4Mux_h I__6320 (
            .O(N__28111),
            .I(N__28093));
    LocalMux I__6319 (
            .O(N__28108),
            .I(N__28090));
    InMux I__6318 (
            .O(N__28105),
            .I(N__28087));
    Span4Mux_h I__6317 (
            .O(N__28100),
            .I(N__28082));
    LocalMux I__6316 (
            .O(N__28097),
            .I(N__28082));
    InMux I__6315 (
            .O(N__28096),
            .I(N__28079));
    Span4Mux_h I__6314 (
            .O(N__28093),
            .I(N__28074));
    Span4Mux_h I__6313 (
            .O(N__28090),
            .I(N__28074));
    LocalMux I__6312 (
            .O(N__28087),
            .I(\c0.data_in_field_87 ));
    Odrv4 I__6311 (
            .O(N__28082),
            .I(\c0.data_in_field_87 ));
    LocalMux I__6310 (
            .O(N__28079),
            .I(\c0.data_in_field_87 ));
    Odrv4 I__6309 (
            .O(N__28074),
            .I(\c0.data_in_field_87 ));
    InMux I__6308 (
            .O(N__28065),
            .I(N__28062));
    LocalMux I__6307 (
            .O(N__28062),
            .I(N__28059));
    Span4Mux_v I__6306 (
            .O(N__28059),
            .I(N__28055));
    InMux I__6305 (
            .O(N__28058),
            .I(N__28052));
    Sp12to4 I__6304 (
            .O(N__28055),
            .I(N__28049));
    LocalMux I__6303 (
            .O(N__28052),
            .I(N__28046));
    Span12Mux_s10_h I__6302 (
            .O(N__28049),
            .I(N__28040));
    Span4Mux_v I__6301 (
            .O(N__28046),
            .I(N__28037));
    InMux I__6300 (
            .O(N__28045),
            .I(N__28032));
    InMux I__6299 (
            .O(N__28044),
            .I(N__28032));
    InMux I__6298 (
            .O(N__28043),
            .I(N__28029));
    Odrv12 I__6297 (
            .O(N__28040),
            .I(\c0.data_in_field_128 ));
    Odrv4 I__6296 (
            .O(N__28037),
            .I(\c0.data_in_field_128 ));
    LocalMux I__6295 (
            .O(N__28032),
            .I(\c0.data_in_field_128 ));
    LocalMux I__6294 (
            .O(N__28029),
            .I(\c0.data_in_field_128 ));
    InMux I__6293 (
            .O(N__28020),
            .I(N__28017));
    LocalMux I__6292 (
            .O(N__28017),
            .I(N__28013));
    InMux I__6291 (
            .O(N__28016),
            .I(N__28010));
    Odrv12 I__6290 (
            .O(N__28013),
            .I(\c0.n2068 ));
    LocalMux I__6289 (
            .O(N__28010),
            .I(\c0.n2068 ));
    InMux I__6288 (
            .O(N__28005),
            .I(N__28002));
    LocalMux I__6287 (
            .O(N__28002),
            .I(N__27998));
    InMux I__6286 (
            .O(N__28001),
            .I(N__27995));
    Span4Mux_h I__6285 (
            .O(N__27998),
            .I(N__27991));
    LocalMux I__6284 (
            .O(N__27995),
            .I(N__27988));
    InMux I__6283 (
            .O(N__27994),
            .I(N__27983));
    Span4Mux_h I__6282 (
            .O(N__27991),
            .I(N__27980));
    Span4Mux_h I__6281 (
            .O(N__27988),
            .I(N__27977));
    InMux I__6280 (
            .O(N__27987),
            .I(N__27974));
    InMux I__6279 (
            .O(N__27986),
            .I(N__27971));
    LocalMux I__6278 (
            .O(N__27983),
            .I(\c0.data_in_field_46 ));
    Odrv4 I__6277 (
            .O(N__27980),
            .I(\c0.data_in_field_46 ));
    Odrv4 I__6276 (
            .O(N__27977),
            .I(\c0.data_in_field_46 ));
    LocalMux I__6275 (
            .O(N__27974),
            .I(\c0.data_in_field_46 ));
    LocalMux I__6274 (
            .O(N__27971),
            .I(\c0.data_in_field_46 ));
    CascadeMux I__6273 (
            .O(N__27960),
            .I(\c0.n1965_cascade_ ));
    InMux I__6272 (
            .O(N__27957),
            .I(N__27954));
    LocalMux I__6271 (
            .O(N__27954),
            .I(N__27948));
    InMux I__6270 (
            .O(N__27953),
            .I(N__27945));
    InMux I__6269 (
            .O(N__27952),
            .I(N__27942));
    InMux I__6268 (
            .O(N__27951),
            .I(N__27937));
    Span4Mux_h I__6267 (
            .O(N__27948),
            .I(N__27934));
    LocalMux I__6266 (
            .O(N__27945),
            .I(N__27931));
    LocalMux I__6265 (
            .O(N__27942),
            .I(N__27928));
    InMux I__6264 (
            .O(N__27941),
            .I(N__27923));
    InMux I__6263 (
            .O(N__27940),
            .I(N__27923));
    LocalMux I__6262 (
            .O(N__27937),
            .I(N__27916));
    Span4Mux_v I__6261 (
            .O(N__27934),
            .I(N__27916));
    Span4Mux_h I__6260 (
            .O(N__27931),
            .I(N__27916));
    Odrv4 I__6259 (
            .O(N__27928),
            .I(\c0.data_in_field_91 ));
    LocalMux I__6258 (
            .O(N__27923),
            .I(\c0.data_in_field_91 ));
    Odrv4 I__6257 (
            .O(N__27916),
            .I(\c0.data_in_field_91 ));
    InMux I__6256 (
            .O(N__27909),
            .I(N__27906));
    LocalMux I__6255 (
            .O(N__27906),
            .I(N__27903));
    Odrv4 I__6254 (
            .O(N__27903),
            .I(\c0.n24_adj_1930 ));
    CascadeMux I__6253 (
            .O(N__27900),
            .I(N__27897));
    InMux I__6252 (
            .O(N__27897),
            .I(N__27893));
    InMux I__6251 (
            .O(N__27896),
            .I(N__27890));
    LocalMux I__6250 (
            .O(N__27893),
            .I(N__27886));
    LocalMux I__6249 (
            .O(N__27890),
            .I(N__27883));
    InMux I__6248 (
            .O(N__27889),
            .I(N__27879));
    Span4Mux_h I__6247 (
            .O(N__27886),
            .I(N__27876));
    Span12Mux_s10_h I__6246 (
            .O(N__27883),
            .I(N__27873));
    InMux I__6245 (
            .O(N__27882),
            .I(N__27870));
    LocalMux I__6244 (
            .O(N__27879),
            .I(data_in_3_5));
    Odrv4 I__6243 (
            .O(N__27876),
            .I(data_in_3_5));
    Odrv12 I__6242 (
            .O(N__27873),
            .I(data_in_3_5));
    LocalMux I__6241 (
            .O(N__27870),
            .I(data_in_3_5));
    InMux I__6240 (
            .O(N__27861),
            .I(N__27858));
    LocalMux I__6239 (
            .O(N__27858),
            .I(N__27853));
    InMux I__6238 (
            .O(N__27857),
            .I(N__27850));
    InMux I__6237 (
            .O(N__27856),
            .I(N__27847));
    Span4Mux_h I__6236 (
            .O(N__27853),
            .I(N__27844));
    LocalMux I__6235 (
            .O(N__27850),
            .I(N__27840));
    LocalMux I__6234 (
            .O(N__27847),
            .I(N__27837));
    Sp12to4 I__6233 (
            .O(N__27844),
            .I(N__27834));
    InMux I__6232 (
            .O(N__27843),
            .I(N__27831));
    Span4Mux_h I__6231 (
            .O(N__27840),
            .I(N__27828));
    Odrv4 I__6230 (
            .O(N__27837),
            .I(data_in_3_0));
    Odrv12 I__6229 (
            .O(N__27834),
            .I(data_in_3_0));
    LocalMux I__6228 (
            .O(N__27831),
            .I(data_in_3_0));
    Odrv4 I__6227 (
            .O(N__27828),
            .I(data_in_3_0));
    InMux I__6226 (
            .O(N__27819),
            .I(N__27816));
    LocalMux I__6225 (
            .O(N__27816),
            .I(N__27811));
    CascadeMux I__6224 (
            .O(N__27815),
            .I(N__27808));
    InMux I__6223 (
            .O(N__27814),
            .I(N__27805));
    Span4Mux_h I__6222 (
            .O(N__27811),
            .I(N__27802));
    InMux I__6221 (
            .O(N__27808),
            .I(N__27799));
    LocalMux I__6220 (
            .O(N__27805),
            .I(N__27796));
    Span4Mux_v I__6219 (
            .O(N__27802),
            .I(N__27792));
    LocalMux I__6218 (
            .O(N__27799),
            .I(N__27787));
    Span4Mux_h I__6217 (
            .O(N__27796),
            .I(N__27787));
    InMux I__6216 (
            .O(N__27795),
            .I(N__27784));
    Span4Mux_v I__6215 (
            .O(N__27792),
            .I(N__27781));
    Span4Mux_h I__6214 (
            .O(N__27787),
            .I(N__27778));
    LocalMux I__6213 (
            .O(N__27784),
            .I(data_in_2_6));
    Odrv4 I__6212 (
            .O(N__27781),
            .I(data_in_2_6));
    Odrv4 I__6211 (
            .O(N__27778),
            .I(data_in_2_6));
    InMux I__6210 (
            .O(N__27771),
            .I(N__27768));
    LocalMux I__6209 (
            .O(N__27768),
            .I(N__27765));
    Span4Mux_v I__6208 (
            .O(N__27765),
            .I(N__27762));
    Span4Mux_h I__6207 (
            .O(N__27762),
            .I(N__27759));
    Odrv4 I__6206 (
            .O(N__27759),
            .I(\c0.n28_adj_1925 ));
    InMux I__6205 (
            .O(N__27756),
            .I(N__27750));
    InMux I__6204 (
            .O(N__27755),
            .I(N__27738));
    InMux I__6203 (
            .O(N__27754),
            .I(N__27738));
    InMux I__6202 (
            .O(N__27753),
            .I(N__27735));
    LocalMux I__6201 (
            .O(N__27750),
            .I(N__27732));
    InMux I__6200 (
            .O(N__27749),
            .I(N__27729));
    InMux I__6199 (
            .O(N__27748),
            .I(N__27726));
    InMux I__6198 (
            .O(N__27747),
            .I(N__27721));
    InMux I__6197 (
            .O(N__27746),
            .I(N__27721));
    InMux I__6196 (
            .O(N__27745),
            .I(N__27713));
    InMux I__6195 (
            .O(N__27744),
            .I(N__27710));
    InMux I__6194 (
            .O(N__27743),
            .I(N__27707));
    LocalMux I__6193 (
            .O(N__27738),
            .I(N__27704));
    LocalMux I__6192 (
            .O(N__27735),
            .I(N__27691));
    Span4Mux_s2_h I__6191 (
            .O(N__27732),
            .I(N__27691));
    LocalMux I__6190 (
            .O(N__27729),
            .I(N__27691));
    LocalMux I__6189 (
            .O(N__27726),
            .I(N__27691));
    LocalMux I__6188 (
            .O(N__27721),
            .I(N__27691));
    InMux I__6187 (
            .O(N__27720),
            .I(N__27688));
    InMux I__6186 (
            .O(N__27719),
            .I(N__27680));
    InMux I__6185 (
            .O(N__27718),
            .I(N__27677));
    InMux I__6184 (
            .O(N__27717),
            .I(N__27674));
    InMux I__6183 (
            .O(N__27716),
            .I(N__27671));
    LocalMux I__6182 (
            .O(N__27713),
            .I(N__27668));
    LocalMux I__6181 (
            .O(N__27710),
            .I(N__27658));
    LocalMux I__6180 (
            .O(N__27707),
            .I(N__27658));
    Span4Mux_v I__6179 (
            .O(N__27704),
            .I(N__27655));
    InMux I__6178 (
            .O(N__27703),
            .I(N__27652));
    CascadeMux I__6177 (
            .O(N__27702),
            .I(N__27649));
    Span4Mux_v I__6176 (
            .O(N__27691),
            .I(N__27641));
    LocalMux I__6175 (
            .O(N__27688),
            .I(N__27641));
    InMux I__6174 (
            .O(N__27687),
            .I(N__27636));
    InMux I__6173 (
            .O(N__27686),
            .I(N__27636));
    InMux I__6172 (
            .O(N__27685),
            .I(N__27629));
    InMux I__6171 (
            .O(N__27684),
            .I(N__27624));
    InMux I__6170 (
            .O(N__27683),
            .I(N__27624));
    LocalMux I__6169 (
            .O(N__27680),
            .I(N__27621));
    LocalMux I__6168 (
            .O(N__27677),
            .I(N__27614));
    LocalMux I__6167 (
            .O(N__27674),
            .I(N__27614));
    LocalMux I__6166 (
            .O(N__27671),
            .I(N__27614));
    Span4Mux_v I__6165 (
            .O(N__27668),
            .I(N__27609));
    InMux I__6164 (
            .O(N__27667),
            .I(N__27604));
    InMux I__6163 (
            .O(N__27666),
            .I(N__27601));
    InMux I__6162 (
            .O(N__27665),
            .I(N__27598));
    InMux I__6161 (
            .O(N__27664),
            .I(N__27595));
    InMux I__6160 (
            .O(N__27663),
            .I(N__27592));
    Span4Mux_v I__6159 (
            .O(N__27658),
            .I(N__27585));
    Span4Mux_v I__6158 (
            .O(N__27655),
            .I(N__27585));
    LocalMux I__6157 (
            .O(N__27652),
            .I(N__27585));
    InMux I__6156 (
            .O(N__27649),
            .I(N__27582));
    InMux I__6155 (
            .O(N__27648),
            .I(N__27579));
    InMux I__6154 (
            .O(N__27647),
            .I(N__27574));
    InMux I__6153 (
            .O(N__27646),
            .I(N__27574));
    Span4Mux_h I__6152 (
            .O(N__27641),
            .I(N__27569));
    LocalMux I__6151 (
            .O(N__27636),
            .I(N__27569));
    InMux I__6150 (
            .O(N__27635),
            .I(N__27565));
    InMux I__6149 (
            .O(N__27634),
            .I(N__27558));
    InMux I__6148 (
            .O(N__27633),
            .I(N__27558));
    InMux I__6147 (
            .O(N__27632),
            .I(N__27558));
    LocalMux I__6146 (
            .O(N__27629),
            .I(N__27554));
    LocalMux I__6145 (
            .O(N__27624),
            .I(N__27547));
    Span4Mux_v I__6144 (
            .O(N__27621),
            .I(N__27547));
    Span4Mux_v I__6143 (
            .O(N__27614),
            .I(N__27547));
    InMux I__6142 (
            .O(N__27613),
            .I(N__27543));
    InMux I__6141 (
            .O(N__27612),
            .I(N__27540));
    Sp12to4 I__6140 (
            .O(N__27609),
            .I(N__27537));
    InMux I__6139 (
            .O(N__27608),
            .I(N__27534));
    InMux I__6138 (
            .O(N__27607),
            .I(N__27531));
    LocalMux I__6137 (
            .O(N__27604),
            .I(N__27528));
    LocalMux I__6136 (
            .O(N__27601),
            .I(N__27517));
    LocalMux I__6135 (
            .O(N__27598),
            .I(N__27517));
    LocalMux I__6134 (
            .O(N__27595),
            .I(N__27517));
    LocalMux I__6133 (
            .O(N__27592),
            .I(N__27517));
    Span4Mux_h I__6132 (
            .O(N__27585),
            .I(N__27517));
    LocalMux I__6131 (
            .O(N__27582),
            .I(N__27514));
    LocalMux I__6130 (
            .O(N__27579),
            .I(N__27507));
    LocalMux I__6129 (
            .O(N__27574),
            .I(N__27507));
    Span4Mux_v I__6128 (
            .O(N__27569),
            .I(N__27507));
    InMux I__6127 (
            .O(N__27568),
            .I(N__27504));
    LocalMux I__6126 (
            .O(N__27565),
            .I(N__27501));
    LocalMux I__6125 (
            .O(N__27558),
            .I(N__27498));
    InMux I__6124 (
            .O(N__27557),
            .I(N__27495));
    Span4Mux_v I__6123 (
            .O(N__27554),
            .I(N__27490));
    Span4Mux_v I__6122 (
            .O(N__27547),
            .I(N__27490));
    InMux I__6121 (
            .O(N__27546),
            .I(N__27487));
    LocalMux I__6120 (
            .O(N__27543),
            .I(N__27482));
    LocalMux I__6119 (
            .O(N__27540),
            .I(N__27482));
    Span12Mux_h I__6118 (
            .O(N__27537),
            .I(N__27477));
    LocalMux I__6117 (
            .O(N__27534),
            .I(N__27477));
    LocalMux I__6116 (
            .O(N__27531),
            .I(N__27470));
    Span4Mux_v I__6115 (
            .O(N__27528),
            .I(N__27470));
    Span4Mux_h I__6114 (
            .O(N__27517),
            .I(N__27470));
    Span4Mux_v I__6113 (
            .O(N__27514),
            .I(N__27465));
    Span4Mux_h I__6112 (
            .O(N__27507),
            .I(N__27465));
    LocalMux I__6111 (
            .O(N__27504),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__6110 (
            .O(N__27501),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__6109 (
            .O(N__27498),
            .I(\c0.byte_transmit_counter2_0 ));
    LocalMux I__6108 (
            .O(N__27495),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__6107 (
            .O(N__27490),
            .I(\c0.byte_transmit_counter2_0 ));
    LocalMux I__6106 (
            .O(N__27487),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv12 I__6105 (
            .O(N__27482),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv12 I__6104 (
            .O(N__27477),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__6103 (
            .O(N__27470),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__6102 (
            .O(N__27465),
            .I(\c0.byte_transmit_counter2_0 ));
    InMux I__6101 (
            .O(N__27444),
            .I(N__27439));
    InMux I__6100 (
            .O(N__27443),
            .I(N__27436));
    InMux I__6099 (
            .O(N__27442),
            .I(N__27432));
    LocalMux I__6098 (
            .O(N__27439),
            .I(N__27429));
    LocalMux I__6097 (
            .O(N__27436),
            .I(N__27426));
    InMux I__6096 (
            .O(N__27435),
            .I(N__27423));
    LocalMux I__6095 (
            .O(N__27432),
            .I(\c0.data_in_field_24 ));
    Odrv4 I__6094 (
            .O(N__27429),
            .I(\c0.data_in_field_24 ));
    Odrv4 I__6093 (
            .O(N__27426),
            .I(\c0.data_in_field_24 ));
    LocalMux I__6092 (
            .O(N__27423),
            .I(\c0.data_in_field_24 ));
    CascadeMux I__6091 (
            .O(N__27414),
            .I(N__27411));
    InMux I__6090 (
            .O(N__27411),
            .I(N__27408));
    LocalMux I__6089 (
            .O(N__27408),
            .I(N__27405));
    Span12Mux_s1_h I__6088 (
            .O(N__27405),
            .I(N__27402));
    Odrv12 I__6087 (
            .O(N__27402),
            .I(\c0.n6039 ));
    InMux I__6086 (
            .O(N__27399),
            .I(N__27396));
    LocalMux I__6085 (
            .O(N__27396),
            .I(N__27392));
    CascadeMux I__6084 (
            .O(N__27395),
            .I(N__27389));
    Span4Mux_h I__6083 (
            .O(N__27392),
            .I(N__27386));
    InMux I__6082 (
            .O(N__27389),
            .I(N__27383));
    Span4Mux_v I__6081 (
            .O(N__27386),
            .I(N__27380));
    LocalMux I__6080 (
            .O(N__27383),
            .I(N__27376));
    Span4Mux_h I__6079 (
            .O(N__27380),
            .I(N__27373));
    InMux I__6078 (
            .O(N__27379),
            .I(N__27370));
    Odrv12 I__6077 (
            .O(N__27376),
            .I(data_in_17_4));
    Odrv4 I__6076 (
            .O(N__27373),
            .I(data_in_17_4));
    LocalMux I__6075 (
            .O(N__27370),
            .I(data_in_17_4));
    CascadeMux I__6074 (
            .O(N__27363),
            .I(N__27360));
    InMux I__6073 (
            .O(N__27360),
            .I(N__27357));
    LocalMux I__6072 (
            .O(N__27357),
            .I(N__27353));
    InMux I__6071 (
            .O(N__27356),
            .I(N__27350));
    Span4Mux_v I__6070 (
            .O(N__27353),
            .I(N__27347));
    LocalMux I__6069 (
            .O(N__27350),
            .I(N__27344));
    Span4Mux_h I__6068 (
            .O(N__27347),
            .I(N__27340));
    Span4Mux_h I__6067 (
            .O(N__27344),
            .I(N__27337));
    InMux I__6066 (
            .O(N__27343),
            .I(N__27334));
    Odrv4 I__6065 (
            .O(N__27340),
            .I(data_in_5_4));
    Odrv4 I__6064 (
            .O(N__27337),
            .I(data_in_5_4));
    LocalMux I__6063 (
            .O(N__27334),
            .I(data_in_5_4));
    InMux I__6062 (
            .O(N__27327),
            .I(N__27323));
    InMux I__6061 (
            .O(N__27326),
            .I(N__27320));
    LocalMux I__6060 (
            .O(N__27323),
            .I(N__27317));
    LocalMux I__6059 (
            .O(N__27320),
            .I(N__27314));
    Span4Mux_v I__6058 (
            .O(N__27317),
            .I(N__27311));
    Span4Mux_v I__6057 (
            .O(N__27314),
            .I(N__27306));
    Span4Mux_h I__6056 (
            .O(N__27311),
            .I(N__27306));
    Span4Mux_h I__6055 (
            .O(N__27306),
            .I(N__27303));
    Odrv4 I__6054 (
            .O(N__27303),
            .I(\c0.n5560 ));
    InMux I__6053 (
            .O(N__27300),
            .I(N__27296));
    CascadeMux I__6052 (
            .O(N__27299),
            .I(N__27293));
    LocalMux I__6051 (
            .O(N__27296),
            .I(N__27290));
    InMux I__6050 (
            .O(N__27293),
            .I(N__27287));
    Span4Mux_v I__6049 (
            .O(N__27290),
            .I(N__27281));
    LocalMux I__6048 (
            .O(N__27287),
            .I(N__27278));
    InMux I__6047 (
            .O(N__27286),
            .I(N__27271));
    InMux I__6046 (
            .O(N__27285),
            .I(N__27271));
    InMux I__6045 (
            .O(N__27284),
            .I(N__27271));
    Sp12to4 I__6044 (
            .O(N__27281),
            .I(N__27268));
    Odrv4 I__6043 (
            .O(N__27278),
            .I(\c0.data_in_field_106 ));
    LocalMux I__6042 (
            .O(N__27271),
            .I(\c0.data_in_field_106 ));
    Odrv12 I__6041 (
            .O(N__27268),
            .I(\c0.data_in_field_106 ));
    InMux I__6040 (
            .O(N__27261),
            .I(N__27257));
    CascadeMux I__6039 (
            .O(N__27260),
            .I(N__27254));
    LocalMux I__6038 (
            .O(N__27257),
            .I(N__27251));
    InMux I__6037 (
            .O(N__27254),
            .I(N__27248));
    Span4Mux_v I__6036 (
            .O(N__27251),
            .I(N__27243));
    LocalMux I__6035 (
            .O(N__27248),
            .I(N__27243));
    Span4Mux_h I__6034 (
            .O(N__27243),
            .I(N__27238));
    CascadeMux I__6033 (
            .O(N__27242),
            .I(N__27235));
    InMux I__6032 (
            .O(N__27241),
            .I(N__27231));
    Span4Mux_h I__6031 (
            .O(N__27238),
            .I(N__27228));
    InMux I__6030 (
            .O(N__27235),
            .I(N__27225));
    InMux I__6029 (
            .O(N__27234),
            .I(N__27222));
    LocalMux I__6028 (
            .O(N__27231),
            .I(\c0.data_in_field_2 ));
    Odrv4 I__6027 (
            .O(N__27228),
            .I(\c0.data_in_field_2 ));
    LocalMux I__6026 (
            .O(N__27225),
            .I(\c0.data_in_field_2 ));
    LocalMux I__6025 (
            .O(N__27222),
            .I(\c0.data_in_field_2 ));
    CascadeMux I__6024 (
            .O(N__27213),
            .I(\c0.n5560_cascade_ ));
    InMux I__6023 (
            .O(N__27210),
            .I(N__27207));
    LocalMux I__6022 (
            .O(N__27207),
            .I(N__27204));
    Span4Mux_h I__6021 (
            .O(N__27204),
            .I(N__27201));
    Span4Mux_h I__6020 (
            .O(N__27201),
            .I(N__27198));
    Odrv4 I__6019 (
            .O(N__27198),
            .I(\c0.n34 ));
    InMux I__6018 (
            .O(N__27195),
            .I(N__27192));
    LocalMux I__6017 (
            .O(N__27192),
            .I(N__27189));
    Span4Mux_v I__6016 (
            .O(N__27189),
            .I(N__27185));
    InMux I__6015 (
            .O(N__27188),
            .I(N__27182));
    Span4Mux_h I__6014 (
            .O(N__27185),
            .I(N__27176));
    LocalMux I__6013 (
            .O(N__27182),
            .I(N__27176));
    InMux I__6012 (
            .O(N__27181),
            .I(N__27173));
    Odrv4 I__6011 (
            .O(N__27176),
            .I(data_in_5_7));
    LocalMux I__6010 (
            .O(N__27173),
            .I(data_in_5_7));
    InMux I__6009 (
            .O(N__27168),
            .I(N__27165));
    LocalMux I__6008 (
            .O(N__27165),
            .I(N__27161));
    InMux I__6007 (
            .O(N__27164),
            .I(N__27158));
    Span4Mux_v I__6006 (
            .O(N__27161),
            .I(N__27153));
    LocalMux I__6005 (
            .O(N__27158),
            .I(N__27150));
    InMux I__6004 (
            .O(N__27157),
            .I(N__27145));
    InMux I__6003 (
            .O(N__27156),
            .I(N__27145));
    Odrv4 I__6002 (
            .O(N__27153),
            .I(\c0.data_in_field_133 ));
    Odrv12 I__6001 (
            .O(N__27150),
            .I(\c0.data_in_field_133 ));
    LocalMux I__6000 (
            .O(N__27145),
            .I(\c0.data_in_field_133 ));
    InMux I__5999 (
            .O(N__27138),
            .I(N__27134));
    CascadeMux I__5998 (
            .O(N__27137),
            .I(N__27128));
    LocalMux I__5997 (
            .O(N__27134),
            .I(N__27125));
    InMux I__5996 (
            .O(N__27133),
            .I(N__27120));
    InMux I__5995 (
            .O(N__27132),
            .I(N__27120));
    InMux I__5994 (
            .O(N__27131),
            .I(N__27115));
    InMux I__5993 (
            .O(N__27128),
            .I(N__27115));
    Span4Mux_v I__5992 (
            .O(N__27125),
            .I(N__27112));
    LocalMux I__5991 (
            .O(N__27120),
            .I(N__27109));
    LocalMux I__5990 (
            .O(N__27115),
            .I(N__27104));
    Span4Mux_h I__5989 (
            .O(N__27112),
            .I(N__27104));
    Odrv12 I__5988 (
            .O(N__27109),
            .I(\c0.data_in_field_21 ));
    Odrv4 I__5987 (
            .O(N__27104),
            .I(\c0.data_in_field_21 ));
    InMux I__5986 (
            .O(N__27099),
            .I(N__27094));
    InMux I__5985 (
            .O(N__27098),
            .I(N__27091));
    InMux I__5984 (
            .O(N__27097),
            .I(N__27088));
    LocalMux I__5983 (
            .O(N__27094),
            .I(N__27085));
    LocalMux I__5982 (
            .O(N__27091),
            .I(N__27081));
    LocalMux I__5981 (
            .O(N__27088),
            .I(N__27078));
    Span4Mux_h I__5980 (
            .O(N__27085),
            .I(N__27075));
    InMux I__5979 (
            .O(N__27084),
            .I(N__27072));
    Span4Mux_s3_h I__5978 (
            .O(N__27081),
            .I(N__27067));
    Span4Mux_h I__5977 (
            .O(N__27078),
            .I(N__27064));
    Span4Mux_h I__5976 (
            .O(N__27075),
            .I(N__27061));
    LocalMux I__5975 (
            .O(N__27072),
            .I(N__27058));
    InMux I__5974 (
            .O(N__27071),
            .I(N__27053));
    InMux I__5973 (
            .O(N__27070),
            .I(N__27053));
    Odrv4 I__5972 (
            .O(N__27067),
            .I(\c0.data_in_field_143 ));
    Odrv4 I__5971 (
            .O(N__27064),
            .I(\c0.data_in_field_143 ));
    Odrv4 I__5970 (
            .O(N__27061),
            .I(\c0.data_in_field_143 ));
    Odrv4 I__5969 (
            .O(N__27058),
            .I(\c0.data_in_field_143 ));
    LocalMux I__5968 (
            .O(N__27053),
            .I(\c0.data_in_field_143 ));
    InMux I__5967 (
            .O(N__27042),
            .I(N__27039));
    LocalMux I__5966 (
            .O(N__27039),
            .I(N__27036));
    Span4Mux_h I__5965 (
            .O(N__27036),
            .I(N__27033));
    Span4Mux_h I__5964 (
            .O(N__27033),
            .I(N__27029));
    InMux I__5963 (
            .O(N__27032),
            .I(N__27026));
    Odrv4 I__5962 (
            .O(N__27029),
            .I(\c0.n5378 ));
    LocalMux I__5961 (
            .O(N__27026),
            .I(\c0.n5378 ));
    CascadeMux I__5960 (
            .O(N__27021),
            .I(N__27018));
    InMux I__5959 (
            .O(N__27018),
            .I(N__27015));
    LocalMux I__5958 (
            .O(N__27015),
            .I(N__27011));
    InMux I__5957 (
            .O(N__27014),
            .I(N__27008));
    Span4Mux_v I__5956 (
            .O(N__27011),
            .I(N__27004));
    LocalMux I__5955 (
            .O(N__27008),
            .I(N__27001));
    InMux I__5954 (
            .O(N__27007),
            .I(N__26998));
    Odrv4 I__5953 (
            .O(N__27004),
            .I(data_in_11_5));
    Odrv4 I__5952 (
            .O(N__27001),
            .I(data_in_11_5));
    LocalMux I__5951 (
            .O(N__26998),
            .I(data_in_11_5));
    InMux I__5950 (
            .O(N__26991),
            .I(N__26987));
    CascadeMux I__5949 (
            .O(N__26990),
            .I(N__26983));
    LocalMux I__5948 (
            .O(N__26987),
            .I(N__26979));
    InMux I__5947 (
            .O(N__26986),
            .I(N__26974));
    InMux I__5946 (
            .O(N__26983),
            .I(N__26974));
    InMux I__5945 (
            .O(N__26982),
            .I(N__26971));
    Odrv4 I__5944 (
            .O(N__26979),
            .I(\c0.data_in_field_55 ));
    LocalMux I__5943 (
            .O(N__26974),
            .I(\c0.data_in_field_55 ));
    LocalMux I__5942 (
            .O(N__26971),
            .I(\c0.data_in_field_55 ));
    InMux I__5941 (
            .O(N__26964),
            .I(N__26961));
    LocalMux I__5940 (
            .O(N__26961),
            .I(N__26956));
    InMux I__5939 (
            .O(N__26960),
            .I(N__26953));
    InMux I__5938 (
            .O(N__26959),
            .I(N__26948));
    Span4Mux_v I__5937 (
            .O(N__26956),
            .I(N__26945));
    LocalMux I__5936 (
            .O(N__26953),
            .I(N__26942));
    InMux I__5935 (
            .O(N__26952),
            .I(N__26937));
    InMux I__5934 (
            .O(N__26951),
            .I(N__26937));
    LocalMux I__5933 (
            .O(N__26948),
            .I(N__26934));
    Odrv4 I__5932 (
            .O(N__26945),
            .I(\c0.data_in_field_63 ));
    Odrv4 I__5931 (
            .O(N__26942),
            .I(\c0.data_in_field_63 ));
    LocalMux I__5930 (
            .O(N__26937),
            .I(\c0.data_in_field_63 ));
    Odrv12 I__5929 (
            .O(N__26934),
            .I(\c0.data_in_field_63 ));
    InMux I__5928 (
            .O(N__26925),
            .I(N__26922));
    LocalMux I__5927 (
            .O(N__26922),
            .I(N__26919));
    Span12Mux_s11_h I__5926 (
            .O(N__26919),
            .I(N__26914));
    InMux I__5925 (
            .O(N__26918),
            .I(N__26909));
    InMux I__5924 (
            .O(N__26917),
            .I(N__26909));
    Odrv12 I__5923 (
            .O(N__26914),
            .I(data_in_14_4));
    LocalMux I__5922 (
            .O(N__26909),
            .I(data_in_14_4));
    CascadeMux I__5921 (
            .O(N__26904),
            .I(N__26901));
    InMux I__5920 (
            .O(N__26901),
            .I(N__26898));
    LocalMux I__5919 (
            .O(N__26898),
            .I(N__26894));
    InMux I__5918 (
            .O(N__26897),
            .I(N__26891));
    Span4Mux_h I__5917 (
            .O(N__26894),
            .I(N__26885));
    LocalMux I__5916 (
            .O(N__26891),
            .I(N__26885));
    InMux I__5915 (
            .O(N__26890),
            .I(N__26882));
    Span4Mux_v I__5914 (
            .O(N__26885),
            .I(N__26879));
    LocalMux I__5913 (
            .O(N__26882),
            .I(N__26874));
    Span4Mux_h I__5912 (
            .O(N__26879),
            .I(N__26871));
    InMux I__5911 (
            .O(N__26878),
            .I(N__26866));
    InMux I__5910 (
            .O(N__26877),
            .I(N__26866));
    Odrv12 I__5909 (
            .O(N__26874),
            .I(\c0.data_in_field_48 ));
    Odrv4 I__5908 (
            .O(N__26871),
            .I(\c0.data_in_field_48 ));
    LocalMux I__5907 (
            .O(N__26866),
            .I(\c0.data_in_field_48 ));
    CascadeMux I__5906 (
            .O(N__26859),
            .I(N__26855));
    InMux I__5905 (
            .O(N__26858),
            .I(N__26852));
    InMux I__5904 (
            .O(N__26855),
            .I(N__26849));
    LocalMux I__5903 (
            .O(N__26852),
            .I(N__26845));
    LocalMux I__5902 (
            .O(N__26849),
            .I(N__26842));
    InMux I__5901 (
            .O(N__26848),
            .I(N__26839));
    Span4Mux_h I__5900 (
            .O(N__26845),
            .I(N__26836));
    Span4Mux_v I__5899 (
            .O(N__26842),
            .I(N__26833));
    LocalMux I__5898 (
            .O(N__26839),
            .I(N__26830));
    Span4Mux_h I__5897 (
            .O(N__26836),
            .I(N__26825));
    Span4Mux_h I__5896 (
            .O(N__26833),
            .I(N__26822));
    Span12Mux_s6_h I__5895 (
            .O(N__26830),
            .I(N__26819));
    InMux I__5894 (
            .O(N__26829),
            .I(N__26814));
    InMux I__5893 (
            .O(N__26828),
            .I(N__26814));
    Odrv4 I__5892 (
            .O(N__26825),
            .I(\c0.data_in_field_32 ));
    Odrv4 I__5891 (
            .O(N__26822),
            .I(\c0.data_in_field_32 ));
    Odrv12 I__5890 (
            .O(N__26819),
            .I(\c0.data_in_field_32 ));
    LocalMux I__5889 (
            .O(N__26814),
            .I(\c0.data_in_field_32 ));
    InMux I__5888 (
            .O(N__26805),
            .I(N__26802));
    LocalMux I__5887 (
            .O(N__26802),
            .I(N__26796));
    InMux I__5886 (
            .O(N__26801),
            .I(N__26793));
    InMux I__5885 (
            .O(N__26800),
            .I(N__26790));
    InMux I__5884 (
            .O(N__26799),
            .I(N__26786));
    Span4Mux_h I__5883 (
            .O(N__26796),
            .I(N__26783));
    LocalMux I__5882 (
            .O(N__26793),
            .I(N__26780));
    LocalMux I__5881 (
            .O(N__26790),
            .I(N__26777));
    InMux I__5880 (
            .O(N__26789),
            .I(N__26774));
    LocalMux I__5879 (
            .O(N__26786),
            .I(N__26771));
    Span4Mux_h I__5878 (
            .O(N__26783),
            .I(N__26766));
    Span4Mux_h I__5877 (
            .O(N__26780),
            .I(N__26766));
    Span4Mux_h I__5876 (
            .O(N__26777),
            .I(N__26763));
    LocalMux I__5875 (
            .O(N__26774),
            .I(\c0.data_in_field_40 ));
    Odrv12 I__5874 (
            .O(N__26771),
            .I(\c0.data_in_field_40 ));
    Odrv4 I__5873 (
            .O(N__26766),
            .I(\c0.data_in_field_40 ));
    Odrv4 I__5872 (
            .O(N__26763),
            .I(\c0.data_in_field_40 ));
    CascadeMux I__5871 (
            .O(N__26754),
            .I(\c0.n6033_cascade_ ));
    InMux I__5870 (
            .O(N__26751),
            .I(N__26748));
    LocalMux I__5869 (
            .O(N__26748),
            .I(N__26745));
    Span12Mux_v I__5868 (
            .O(N__26745),
            .I(N__26742));
    Odrv12 I__5867 (
            .O(N__26742),
            .I(\c0.n5791 ));
    InMux I__5866 (
            .O(N__26739),
            .I(N__26736));
    LocalMux I__5865 (
            .O(N__26736),
            .I(N__26733));
    Odrv4 I__5864 (
            .O(N__26733),
            .I(\c0.n1814 ));
    CascadeMux I__5863 (
            .O(N__26730),
            .I(N__26727));
    InMux I__5862 (
            .O(N__26727),
            .I(N__26723));
    InMux I__5861 (
            .O(N__26726),
            .I(N__26720));
    LocalMux I__5860 (
            .O(N__26723),
            .I(N__26717));
    LocalMux I__5859 (
            .O(N__26720),
            .I(N__26714));
    Span4Mux_v I__5858 (
            .O(N__26717),
            .I(N__26711));
    Span4Mux_h I__5857 (
            .O(N__26714),
            .I(N__26707));
    Sp12to4 I__5856 (
            .O(N__26711),
            .I(N__26704));
    InMux I__5855 (
            .O(N__26710),
            .I(N__26701));
    Sp12to4 I__5854 (
            .O(N__26707),
            .I(N__26697));
    Span12Mux_s11_h I__5853 (
            .O(N__26704),
            .I(N__26692));
    LocalMux I__5852 (
            .O(N__26701),
            .I(N__26692));
    InMux I__5851 (
            .O(N__26700),
            .I(N__26689));
    Span12Mux_v I__5850 (
            .O(N__26697),
            .I(N__26686));
    Span12Mux_v I__5849 (
            .O(N__26692),
            .I(N__26683));
    LocalMux I__5848 (
            .O(N__26689),
            .I(data_in_19_1));
    Odrv12 I__5847 (
            .O(N__26686),
            .I(data_in_19_1));
    Odrv12 I__5846 (
            .O(N__26683),
            .I(data_in_19_1));
    InMux I__5845 (
            .O(N__26676),
            .I(N__26672));
    CascadeMux I__5844 (
            .O(N__26675),
            .I(N__26669));
    LocalMux I__5843 (
            .O(N__26672),
            .I(N__26666));
    InMux I__5842 (
            .O(N__26669),
            .I(N__26663));
    Span4Mux_h I__5841 (
            .O(N__26666),
            .I(N__26660));
    LocalMux I__5840 (
            .O(N__26663),
            .I(N__26657));
    Span4Mux_h I__5839 (
            .O(N__26660),
            .I(N__26654));
    Odrv4 I__5838 (
            .O(N__26657),
            .I(\c0.n2143 ));
    Odrv4 I__5837 (
            .O(N__26654),
            .I(\c0.n2143 ));
    CascadeMux I__5836 (
            .O(N__26649),
            .I(\c0.n1814_cascade_ ));
    InMux I__5835 (
            .O(N__26646),
            .I(N__26639));
    CascadeMux I__5834 (
            .O(N__26645),
            .I(N__26636));
    InMux I__5833 (
            .O(N__26644),
            .I(N__26633));
    InMux I__5832 (
            .O(N__26643),
            .I(N__26630));
    InMux I__5831 (
            .O(N__26642),
            .I(N__26627));
    LocalMux I__5830 (
            .O(N__26639),
            .I(N__26624));
    InMux I__5829 (
            .O(N__26636),
            .I(N__26621));
    LocalMux I__5828 (
            .O(N__26633),
            .I(N__26618));
    LocalMux I__5827 (
            .O(N__26630),
            .I(N__26613));
    LocalMux I__5826 (
            .O(N__26627),
            .I(N__26613));
    Span12Mux_v I__5825 (
            .O(N__26624),
            .I(N__26608));
    LocalMux I__5824 (
            .O(N__26621),
            .I(N__26605));
    Span4Mux_h I__5823 (
            .O(N__26618),
            .I(N__26600));
    Span4Mux_v I__5822 (
            .O(N__26613),
            .I(N__26600));
    InMux I__5821 (
            .O(N__26612),
            .I(N__26595));
    InMux I__5820 (
            .O(N__26611),
            .I(N__26595));
    Odrv12 I__5819 (
            .O(N__26608),
            .I(\c0.data_in_field_109 ));
    Odrv4 I__5818 (
            .O(N__26605),
            .I(\c0.data_in_field_109 ));
    Odrv4 I__5817 (
            .O(N__26600),
            .I(\c0.data_in_field_109 ));
    LocalMux I__5816 (
            .O(N__26595),
            .I(\c0.data_in_field_109 ));
    InMux I__5815 (
            .O(N__26586),
            .I(N__26583));
    LocalMux I__5814 (
            .O(N__26583),
            .I(\c0.n32_adj_1901 ));
    InMux I__5813 (
            .O(N__26580),
            .I(N__26576));
    InMux I__5812 (
            .O(N__26579),
            .I(N__26572));
    LocalMux I__5811 (
            .O(N__26576),
            .I(N__26569));
    InMux I__5810 (
            .O(N__26575),
            .I(N__26566));
    LocalMux I__5809 (
            .O(N__26572),
            .I(N__26561));
    Span4Mux_v I__5808 (
            .O(N__26569),
            .I(N__26561));
    LocalMux I__5807 (
            .O(N__26566),
            .I(N__26558));
    Sp12to4 I__5806 (
            .O(N__26561),
            .I(N__26553));
    Span12Mux_s11_h I__5805 (
            .O(N__26558),
            .I(N__26553));
    Odrv12 I__5804 (
            .O(N__26553),
            .I(data_in_8_5));
    CascadeMux I__5803 (
            .O(N__26550),
            .I(N__26547));
    InMux I__5802 (
            .O(N__26547),
            .I(N__26544));
    LocalMux I__5801 (
            .O(N__26544),
            .I(N__26541));
    Odrv4 I__5800 (
            .O(N__26541),
            .I(n318));
    InMux I__5799 (
            .O(N__26538),
            .I(N__26534));
    InMux I__5798 (
            .O(N__26537),
            .I(N__26529));
    LocalMux I__5797 (
            .O(N__26534),
            .I(N__26526));
    InMux I__5796 (
            .O(N__26533),
            .I(N__26523));
    InMux I__5795 (
            .O(N__26532),
            .I(N__26520));
    LocalMux I__5794 (
            .O(N__26529),
            .I(r_Clock_Count_3));
    Odrv4 I__5793 (
            .O(N__26526),
            .I(r_Clock_Count_3));
    LocalMux I__5792 (
            .O(N__26523),
            .I(r_Clock_Count_3));
    LocalMux I__5791 (
            .O(N__26520),
            .I(r_Clock_Count_3));
    CascadeMux I__5790 (
            .O(N__26511),
            .I(N__26508));
    InMux I__5789 (
            .O(N__26508),
            .I(N__26505));
    LocalMux I__5788 (
            .O(N__26505),
            .I(N__26502));
    Odrv4 I__5787 (
            .O(N__26502),
            .I(n321));
    InMux I__5786 (
            .O(N__26499),
            .I(N__26496));
    LocalMux I__5785 (
            .O(N__26496),
            .I(N__26490));
    InMux I__5784 (
            .O(N__26495),
            .I(N__26485));
    InMux I__5783 (
            .O(N__26494),
            .I(N__26485));
    InMux I__5782 (
            .O(N__26493),
            .I(N__26482));
    Odrv4 I__5781 (
            .O(N__26490),
            .I(r_Clock_Count_0));
    LocalMux I__5780 (
            .O(N__26485),
            .I(r_Clock_Count_0));
    LocalMux I__5779 (
            .O(N__26482),
            .I(r_Clock_Count_0));
    InMux I__5778 (
            .O(N__26475),
            .I(N__26471));
    InMux I__5777 (
            .O(N__26474),
            .I(N__26468));
    LocalMux I__5776 (
            .O(N__26471),
            .I(N__26465));
    LocalMux I__5775 (
            .O(N__26468),
            .I(data_out_18_5));
    Odrv12 I__5774 (
            .O(N__26465),
            .I(data_out_18_5));
    InMux I__5773 (
            .O(N__26460),
            .I(N__26451));
    InMux I__5772 (
            .O(N__26459),
            .I(N__26451));
    InMux I__5771 (
            .O(N__26458),
            .I(N__26446));
    InMux I__5770 (
            .O(N__26457),
            .I(N__26446));
    InMux I__5769 (
            .O(N__26456),
            .I(N__26443));
    LocalMux I__5768 (
            .O(N__26451),
            .I(n782));
    LocalMux I__5767 (
            .O(N__26446),
            .I(n782));
    LocalMux I__5766 (
            .O(N__26443),
            .I(n782));
    CascadeMux I__5765 (
            .O(N__26436),
            .I(N__26433));
    InMux I__5764 (
            .O(N__26433),
            .I(N__26430));
    LocalMux I__5763 (
            .O(N__26430),
            .I(N__26427));
    Span4Mux_h I__5762 (
            .O(N__26427),
            .I(N__26424));
    Odrv4 I__5761 (
            .O(N__26424),
            .I(n320));
    InMux I__5760 (
            .O(N__26421),
            .I(N__26418));
    LocalMux I__5759 (
            .O(N__26418),
            .I(N__26414));
    InMux I__5758 (
            .O(N__26417),
            .I(N__26409));
    Span4Mux_v I__5757 (
            .O(N__26414),
            .I(N__26406));
    InMux I__5756 (
            .O(N__26413),
            .I(N__26403));
    InMux I__5755 (
            .O(N__26412),
            .I(N__26400));
    LocalMux I__5754 (
            .O(N__26409),
            .I(r_Clock_Count_1));
    Odrv4 I__5753 (
            .O(N__26406),
            .I(r_Clock_Count_1));
    LocalMux I__5752 (
            .O(N__26403),
            .I(r_Clock_Count_1));
    LocalMux I__5751 (
            .O(N__26400),
            .I(r_Clock_Count_1));
    InMux I__5750 (
            .O(N__26391),
            .I(N__26387));
    CascadeMux I__5749 (
            .O(N__26390),
            .I(N__26384));
    LocalMux I__5748 (
            .O(N__26387),
            .I(N__26381));
    InMux I__5747 (
            .O(N__26384),
            .I(N__26378));
    Odrv12 I__5746 (
            .O(N__26381),
            .I(rx_data_1));
    LocalMux I__5745 (
            .O(N__26378),
            .I(rx_data_1));
    CascadeMux I__5744 (
            .O(N__26373),
            .I(N__26370));
    InMux I__5743 (
            .O(N__26370),
            .I(N__26367));
    LocalMux I__5742 (
            .O(N__26367),
            .I(N__26363));
    InMux I__5741 (
            .O(N__26366),
            .I(N__26360));
    Span4Mux_v I__5740 (
            .O(N__26363),
            .I(N__26357));
    LocalMux I__5739 (
            .O(N__26360),
            .I(N__26354));
    Span4Mux_h I__5738 (
            .O(N__26357),
            .I(N__26350));
    Span12Mux_h I__5737 (
            .O(N__26354),
            .I(N__26347));
    InMux I__5736 (
            .O(N__26353),
            .I(N__26344));
    Odrv4 I__5735 (
            .O(N__26350),
            .I(data_in_14_3));
    Odrv12 I__5734 (
            .O(N__26347),
            .I(data_in_14_3));
    LocalMux I__5733 (
            .O(N__26344),
            .I(data_in_14_3));
    CascadeMux I__5732 (
            .O(N__26337),
            .I(N__26334));
    InMux I__5731 (
            .O(N__26334),
            .I(N__26330));
    InMux I__5730 (
            .O(N__26333),
            .I(N__26327));
    LocalMux I__5729 (
            .O(N__26330),
            .I(N__26322));
    LocalMux I__5728 (
            .O(N__26327),
            .I(N__26322));
    Span4Mux_h I__5727 (
            .O(N__26322),
            .I(N__26318));
    InMux I__5726 (
            .O(N__26321),
            .I(N__26315));
    Span4Mux_h I__5725 (
            .O(N__26318),
            .I(N__26312));
    LocalMux I__5724 (
            .O(N__26315),
            .I(data_in_13_3));
    Odrv4 I__5723 (
            .O(N__26312),
            .I(data_in_13_3));
    CascadeMux I__5722 (
            .O(N__26307),
            .I(\c0.n6309_cascade_ ));
    InMux I__5721 (
            .O(N__26304),
            .I(N__26298));
    InMux I__5720 (
            .O(N__26303),
            .I(N__26298));
    LocalMux I__5719 (
            .O(N__26298),
            .I(data_out_18_2));
    InMux I__5718 (
            .O(N__26295),
            .I(N__26292));
    LocalMux I__5717 (
            .O(N__26292),
            .I(\c0.n1249 ));
    InMux I__5716 (
            .O(N__26289),
            .I(N__26286));
    LocalMux I__5715 (
            .O(N__26286),
            .I(N__26283));
    Odrv12 I__5714 (
            .O(N__26283),
            .I(tx_data_4_N_keep));
    InMux I__5713 (
            .O(N__26280),
            .I(N__26277));
    LocalMux I__5712 (
            .O(N__26277),
            .I(\c0.tx.n3644 ));
    InMux I__5711 (
            .O(N__26274),
            .I(N__26271));
    LocalMux I__5710 (
            .O(N__26271),
            .I(n11_adj_1979));
    CascadeMux I__5709 (
            .O(N__26268),
            .I(n5818_cascade_));
    InMux I__5708 (
            .O(N__26265),
            .I(N__26262));
    LocalMux I__5707 (
            .O(N__26262),
            .I(N__26259));
    Odrv4 I__5706 (
            .O(N__26259),
            .I(n4155));
    CascadeMux I__5705 (
            .O(N__26256),
            .I(n4334_cascade_));
    InMux I__5704 (
            .O(N__26253),
            .I(N__26250));
    LocalMux I__5703 (
            .O(N__26250),
            .I(n1991));
    InMux I__5702 (
            .O(N__26247),
            .I(N__26243));
    InMux I__5701 (
            .O(N__26246),
            .I(N__26240));
    LocalMux I__5700 (
            .O(N__26243),
            .I(data_out_19_7));
    LocalMux I__5699 (
            .O(N__26240),
            .I(data_out_19_7));
    InMux I__5698 (
            .O(N__26235),
            .I(N__26232));
    LocalMux I__5697 (
            .O(N__26232),
            .I(\c0.n17_adj_1950 ));
    InMux I__5696 (
            .O(N__26229),
            .I(N__26226));
    LocalMux I__5695 (
            .O(N__26226),
            .I(n4_adj_1982));
    CascadeMux I__5694 (
            .O(N__26223),
            .I(N__26220));
    InMux I__5693 (
            .O(N__26220),
            .I(N__26217));
    LocalMux I__5692 (
            .O(N__26217),
            .I(\c0.n17_adj_1908 ));
    InMux I__5691 (
            .O(N__26214),
            .I(N__26210));
    InMux I__5690 (
            .O(N__26213),
            .I(N__26207));
    LocalMux I__5689 (
            .O(N__26210),
            .I(data_out_18_7));
    LocalMux I__5688 (
            .O(N__26207),
            .I(data_out_18_7));
    InMux I__5687 (
            .O(N__26202),
            .I(N__26195));
    InMux I__5686 (
            .O(N__26201),
            .I(N__26195));
    InMux I__5685 (
            .O(N__26200),
            .I(N__26192));
    LocalMux I__5684 (
            .O(N__26195),
            .I(\c0.n1508 ));
    LocalMux I__5683 (
            .O(N__26192),
            .I(\c0.n1508 ));
    InMux I__5682 (
            .O(N__26187),
            .I(N__26183));
    InMux I__5681 (
            .O(N__26186),
            .I(N__26180));
    LocalMux I__5680 (
            .O(N__26183),
            .I(N__26177));
    LocalMux I__5679 (
            .O(N__26180),
            .I(data_out_19_2));
    Odrv4 I__5678 (
            .O(N__26177),
            .I(data_out_19_2));
    CascadeMux I__5677 (
            .O(N__26172),
            .I(\c0.n1508_cascade_ ));
    InMux I__5676 (
            .O(N__26169),
            .I(N__26166));
    LocalMux I__5675 (
            .O(N__26166),
            .I(\c0.n5840 ));
    InMux I__5674 (
            .O(N__26163),
            .I(N__26159));
    InMux I__5673 (
            .O(N__26162),
            .I(N__26155));
    LocalMux I__5672 (
            .O(N__26159),
            .I(N__26152));
    InMux I__5671 (
            .O(N__26158),
            .I(N__26149));
    LocalMux I__5670 (
            .O(N__26155),
            .I(N__26146));
    Span4Mux_v I__5669 (
            .O(N__26152),
            .I(N__26143));
    LocalMux I__5668 (
            .O(N__26149),
            .I(data_in_11_7));
    Odrv12 I__5667 (
            .O(N__26146),
            .I(data_in_11_7));
    Odrv4 I__5666 (
            .O(N__26143),
            .I(data_in_11_7));
    CascadeMux I__5665 (
            .O(N__26136),
            .I(n5448_cascade_));
    InMux I__5664 (
            .O(N__26133),
            .I(N__26130));
    LocalMux I__5663 (
            .O(N__26130),
            .I(N__26127));
    Odrv4 I__5662 (
            .O(N__26127),
            .I(n4_adj_1975));
    InMux I__5661 (
            .O(N__26124),
            .I(N__26120));
    InMux I__5660 (
            .O(N__26123),
            .I(N__26117));
    LocalMux I__5659 (
            .O(N__26120),
            .I(data_out_19_4));
    LocalMux I__5658 (
            .O(N__26117),
            .I(data_out_19_4));
    InMux I__5657 (
            .O(N__26112),
            .I(N__26106));
    InMux I__5656 (
            .O(N__26111),
            .I(N__26106));
    LocalMux I__5655 (
            .O(N__26106),
            .I(data_out_18_4));
    InMux I__5654 (
            .O(N__26103),
            .I(N__26100));
    LocalMux I__5653 (
            .O(N__26100),
            .I(N__26096));
    InMux I__5652 (
            .O(N__26099),
            .I(N__26093));
    Span4Mux_h I__5651 (
            .O(N__26096),
            .I(N__26090));
    LocalMux I__5650 (
            .O(N__26093),
            .I(\c0.delay_counter_3 ));
    Odrv4 I__5649 (
            .O(N__26090),
            .I(\c0.delay_counter_3 ));
    InMux I__5648 (
            .O(N__26085),
            .I(N__26082));
    LocalMux I__5647 (
            .O(N__26082),
            .I(N__26078));
    InMux I__5646 (
            .O(N__26081),
            .I(N__26075));
    Span4Mux_h I__5645 (
            .O(N__26078),
            .I(N__26072));
    LocalMux I__5644 (
            .O(N__26075),
            .I(\c0.delay_counter_6 ));
    Odrv4 I__5643 (
            .O(N__26072),
            .I(\c0.delay_counter_6 ));
    CascadeMux I__5642 (
            .O(N__26067),
            .I(N__26064));
    InMux I__5641 (
            .O(N__26064),
            .I(N__26060));
    InMux I__5640 (
            .O(N__26063),
            .I(N__26057));
    LocalMux I__5639 (
            .O(N__26060),
            .I(N__26054));
    LocalMux I__5638 (
            .O(N__26057),
            .I(\c0.delay_counter_10 ));
    Odrv4 I__5637 (
            .O(N__26054),
            .I(\c0.delay_counter_10 ));
    InMux I__5636 (
            .O(N__26049),
            .I(N__26046));
    LocalMux I__5635 (
            .O(N__26046),
            .I(\c0.n18_adj_1919 ));
    InMux I__5634 (
            .O(N__26043),
            .I(N__26040));
    LocalMux I__5633 (
            .O(N__26040),
            .I(N__26036));
    InMux I__5632 (
            .O(N__26039),
            .I(N__26033));
    Span4Mux_h I__5631 (
            .O(N__26036),
            .I(N__26030));
    LocalMux I__5630 (
            .O(N__26033),
            .I(\c0.delay_counter_8 ));
    Odrv4 I__5629 (
            .O(N__26030),
            .I(\c0.delay_counter_8 ));
    InMux I__5628 (
            .O(N__26025),
            .I(N__26022));
    LocalMux I__5627 (
            .O(N__26022),
            .I(N__26018));
    InMux I__5626 (
            .O(N__26021),
            .I(N__26015));
    Span4Mux_v I__5625 (
            .O(N__26018),
            .I(N__26012));
    LocalMux I__5624 (
            .O(N__26015),
            .I(\c0.delay_counter_4 ));
    Odrv4 I__5623 (
            .O(N__26012),
            .I(\c0.delay_counter_4 ));
    CascadeMux I__5622 (
            .O(N__26007),
            .I(\c0.n20_adj_1922_cascade_ ));
    InMux I__5621 (
            .O(N__26004),
            .I(N__26001));
    LocalMux I__5620 (
            .O(N__26001),
            .I(N__25998));
    Odrv4 I__5619 (
            .O(N__25998),
            .I(\c0.n16_adj_1921 ));
    InMux I__5618 (
            .O(N__25995),
            .I(N__25991));
    InMux I__5617 (
            .O(N__25994),
            .I(N__25988));
    LocalMux I__5616 (
            .O(N__25991),
            .I(N__25985));
    LocalMux I__5615 (
            .O(N__25988),
            .I(N__25979));
    Span4Mux_v I__5614 (
            .O(N__25985),
            .I(N__25976));
    CascadeMux I__5613 (
            .O(N__25984),
            .I(N__25973));
    InMux I__5612 (
            .O(N__25983),
            .I(N__25970));
    InMux I__5611 (
            .O(N__25982),
            .I(N__25967));
    Span4Mux_v I__5610 (
            .O(N__25979),
            .I(N__25962));
    Span4Mux_h I__5609 (
            .O(N__25976),
            .I(N__25962));
    InMux I__5608 (
            .O(N__25973),
            .I(N__25959));
    LocalMux I__5607 (
            .O(N__25970),
            .I(\c0.data_in_field_77 ));
    LocalMux I__5606 (
            .O(N__25967),
            .I(\c0.data_in_field_77 ));
    Odrv4 I__5605 (
            .O(N__25962),
            .I(\c0.data_in_field_77 ));
    LocalMux I__5604 (
            .O(N__25959),
            .I(\c0.data_in_field_77 ));
    CascadeMux I__5603 (
            .O(N__25950),
            .I(\c0.n6207_cascade_ ));
    InMux I__5602 (
            .O(N__25947),
            .I(N__25943));
    InMux I__5601 (
            .O(N__25946),
            .I(N__25940));
    LocalMux I__5600 (
            .O(N__25943),
            .I(N__25937));
    LocalMux I__5599 (
            .O(N__25940),
            .I(N__25931));
    Span4Mux_h I__5598 (
            .O(N__25937),
            .I(N__25928));
    InMux I__5597 (
            .O(N__25936),
            .I(N__25921));
    InMux I__5596 (
            .O(N__25935),
            .I(N__25921));
    InMux I__5595 (
            .O(N__25934),
            .I(N__25921));
    Odrv4 I__5594 (
            .O(N__25931),
            .I(\c0.data_in_field_69 ));
    Odrv4 I__5593 (
            .O(N__25928),
            .I(\c0.data_in_field_69 ));
    LocalMux I__5592 (
            .O(N__25921),
            .I(\c0.data_in_field_69 ));
    InMux I__5591 (
            .O(N__25914),
            .I(N__25911));
    LocalMux I__5590 (
            .O(N__25911),
            .I(\c0.n5713 ));
    CascadeMux I__5589 (
            .O(N__25908),
            .I(N__25905));
    InMux I__5588 (
            .O(N__25905),
            .I(N__25902));
    LocalMux I__5587 (
            .O(N__25902),
            .I(N__25898));
    CascadeMux I__5586 (
            .O(N__25901),
            .I(N__25895));
    Span4Mux_h I__5585 (
            .O(N__25898),
            .I(N__25890));
    InMux I__5584 (
            .O(N__25895),
            .I(N__25887));
    InMux I__5583 (
            .O(N__25894),
            .I(N__25882));
    InMux I__5582 (
            .O(N__25893),
            .I(N__25882));
    Span4Mux_h I__5581 (
            .O(N__25890),
            .I(N__25879));
    LocalMux I__5580 (
            .O(N__25887),
            .I(N__25876));
    LocalMux I__5579 (
            .O(N__25882),
            .I(data_in_19_2));
    Odrv4 I__5578 (
            .O(N__25879),
            .I(data_in_19_2));
    Odrv12 I__5577 (
            .O(N__25876),
            .I(data_in_19_2));
    InMux I__5576 (
            .O(N__25869),
            .I(N__25865));
    CascadeMux I__5575 (
            .O(N__25868),
            .I(N__25862));
    LocalMux I__5574 (
            .O(N__25865),
            .I(N__25858));
    InMux I__5573 (
            .O(N__25862),
            .I(N__25855));
    InMux I__5572 (
            .O(N__25861),
            .I(N__25852));
    Span4Mux_h I__5571 (
            .O(N__25858),
            .I(N__25849));
    LocalMux I__5570 (
            .O(N__25855),
            .I(data_in_9_0));
    LocalMux I__5569 (
            .O(N__25852),
            .I(data_in_9_0));
    Odrv4 I__5568 (
            .O(N__25849),
            .I(data_in_9_0));
    InMux I__5567 (
            .O(N__25842),
            .I(N__25839));
    LocalMux I__5566 (
            .O(N__25839),
            .I(N__25836));
    Span4Mux_v I__5565 (
            .O(N__25836),
            .I(N__25832));
    InMux I__5564 (
            .O(N__25835),
            .I(N__25829));
    Span4Mux_h I__5563 (
            .O(N__25832),
            .I(N__25825));
    LocalMux I__5562 (
            .O(N__25829),
            .I(N__25822));
    InMux I__5561 (
            .O(N__25828),
            .I(N__25818));
    Span4Mux_h I__5560 (
            .O(N__25825),
            .I(N__25813));
    Span4Mux_v I__5559 (
            .O(N__25822),
            .I(N__25813));
    InMux I__5558 (
            .O(N__25821),
            .I(N__25810));
    LocalMux I__5557 (
            .O(N__25818),
            .I(\c0.data_in_field_42 ));
    Odrv4 I__5556 (
            .O(N__25813),
            .I(\c0.data_in_field_42 ));
    LocalMux I__5555 (
            .O(N__25810),
            .I(\c0.data_in_field_42 ));
    InMux I__5554 (
            .O(N__25803),
            .I(N__25800));
    LocalMux I__5553 (
            .O(N__25800),
            .I(N__25797));
    Span4Mux_s2_h I__5552 (
            .O(N__25797),
            .I(N__25794));
    Span4Mux_h I__5551 (
            .O(N__25794),
            .I(N__25790));
    InMux I__5550 (
            .O(N__25793),
            .I(N__25784));
    Span4Mux_h I__5549 (
            .O(N__25790),
            .I(N__25781));
    InMux I__5548 (
            .O(N__25789),
            .I(N__25776));
    InMux I__5547 (
            .O(N__25788),
            .I(N__25776));
    InMux I__5546 (
            .O(N__25787),
            .I(N__25773));
    LocalMux I__5545 (
            .O(N__25784),
            .I(\c0.data_in_field_72 ));
    Odrv4 I__5544 (
            .O(N__25781),
            .I(\c0.data_in_field_72 ));
    LocalMux I__5543 (
            .O(N__25776),
            .I(\c0.data_in_field_72 ));
    LocalMux I__5542 (
            .O(N__25773),
            .I(\c0.data_in_field_72 ));
    InMux I__5541 (
            .O(N__25764),
            .I(N__25761));
    LocalMux I__5540 (
            .O(N__25761),
            .I(N__25757));
    InMux I__5539 (
            .O(N__25760),
            .I(N__25753));
    Span4Mux_h I__5538 (
            .O(N__25757),
            .I(N__25750));
    InMux I__5537 (
            .O(N__25756),
            .I(N__25747));
    LocalMux I__5536 (
            .O(N__25753),
            .I(N__25744));
    Span4Mux_h I__5535 (
            .O(N__25750),
            .I(N__25741));
    LocalMux I__5534 (
            .O(N__25747),
            .I(data_in_12_0));
    Odrv12 I__5533 (
            .O(N__25744),
            .I(data_in_12_0));
    Odrv4 I__5532 (
            .O(N__25741),
            .I(data_in_12_0));
    InMux I__5531 (
            .O(N__25734),
            .I(N__25731));
    LocalMux I__5530 (
            .O(N__25731),
            .I(N__25728));
    Span4Mux_v I__5529 (
            .O(N__25728),
            .I(N__25724));
    InMux I__5528 (
            .O(N__25727),
            .I(N__25721));
    Span4Mux_h I__5527 (
            .O(N__25724),
            .I(N__25716));
    LocalMux I__5526 (
            .O(N__25721),
            .I(N__25716));
    Span4Mux_v I__5525 (
            .O(N__25716),
            .I(N__25711));
    InMux I__5524 (
            .O(N__25715),
            .I(N__25708));
    InMux I__5523 (
            .O(N__25714),
            .I(N__25705));
    Span4Mux_h I__5522 (
            .O(N__25711),
            .I(N__25702));
    LocalMux I__5521 (
            .O(N__25708),
            .I(data_in_18_2));
    LocalMux I__5520 (
            .O(N__25705),
            .I(data_in_18_2));
    Odrv4 I__5519 (
            .O(N__25702),
            .I(data_in_18_2));
    InMux I__5518 (
            .O(N__25695),
            .I(N__25692));
    LocalMux I__5517 (
            .O(N__25692),
            .I(N__25688));
    InMux I__5516 (
            .O(N__25691),
            .I(N__25685));
    Span4Mux_v I__5515 (
            .O(N__25688),
            .I(N__25682));
    LocalMux I__5514 (
            .O(N__25685),
            .I(N__25679));
    Span4Mux_h I__5513 (
            .O(N__25682),
            .I(N__25674));
    Span4Mux_h I__5512 (
            .O(N__25679),
            .I(N__25674));
    Span4Mux_h I__5511 (
            .O(N__25674),
            .I(N__25670));
    InMux I__5510 (
            .O(N__25673),
            .I(N__25667));
    Odrv4 I__5509 (
            .O(N__25670),
            .I(data_in_17_2));
    LocalMux I__5508 (
            .O(N__25667),
            .I(data_in_17_2));
    CascadeMux I__5507 (
            .O(N__25662),
            .I(N__25658));
    InMux I__5506 (
            .O(N__25661),
            .I(N__25655));
    InMux I__5505 (
            .O(N__25658),
            .I(N__25652));
    LocalMux I__5504 (
            .O(N__25655),
            .I(N__25647));
    LocalMux I__5503 (
            .O(N__25652),
            .I(N__25647));
    Span4Mux_v I__5502 (
            .O(N__25647),
            .I(N__25644));
    Span4Mux_v I__5501 (
            .O(N__25644),
            .I(N__25640));
    InMux I__5500 (
            .O(N__25643),
            .I(N__25637));
    Span4Mux_h I__5499 (
            .O(N__25640),
            .I(N__25634));
    LocalMux I__5498 (
            .O(N__25637),
            .I(data_in_6_2));
    Odrv4 I__5497 (
            .O(N__25634),
            .I(data_in_6_2));
    CascadeMux I__5496 (
            .O(N__25629),
            .I(N__25625));
    InMux I__5495 (
            .O(N__25628),
            .I(N__25622));
    InMux I__5494 (
            .O(N__25625),
            .I(N__25619));
    LocalMux I__5493 (
            .O(N__25622),
            .I(N__25616));
    LocalMux I__5492 (
            .O(N__25619),
            .I(N__25612));
    Span4Mux_h I__5491 (
            .O(N__25616),
            .I(N__25609));
    InMux I__5490 (
            .O(N__25615),
            .I(N__25606));
    Odrv4 I__5489 (
            .O(N__25612),
            .I(data_in_5_2));
    Odrv4 I__5488 (
            .O(N__25609),
            .I(data_in_5_2));
    LocalMux I__5487 (
            .O(N__25606),
            .I(data_in_5_2));
    CascadeMux I__5486 (
            .O(N__25599),
            .I(N__25596));
    InMux I__5485 (
            .O(N__25596),
            .I(N__25592));
    InMux I__5484 (
            .O(N__25595),
            .I(N__25589));
    LocalMux I__5483 (
            .O(N__25592),
            .I(N__25584));
    LocalMux I__5482 (
            .O(N__25589),
            .I(N__25584));
    Span4Mux_v I__5481 (
            .O(N__25584),
            .I(N__25580));
    InMux I__5480 (
            .O(N__25583),
            .I(N__25577));
    Odrv4 I__5479 (
            .O(N__25580),
            .I(data_in_4_5));
    LocalMux I__5478 (
            .O(N__25577),
            .I(data_in_4_5));
    InMux I__5477 (
            .O(N__25572),
            .I(N__25569));
    LocalMux I__5476 (
            .O(N__25569),
            .I(N__25565));
    InMux I__5475 (
            .O(N__25568),
            .I(N__25562));
    Span4Mux_h I__5474 (
            .O(N__25565),
            .I(N__25559));
    LocalMux I__5473 (
            .O(N__25562),
            .I(N__25556));
    Span4Mux_v I__5472 (
            .O(N__25559),
            .I(N__25550));
    Span4Mux_v I__5471 (
            .O(N__25556),
            .I(N__25550));
    InMux I__5470 (
            .O(N__25555),
            .I(N__25547));
    Span4Mux_h I__5469 (
            .O(N__25550),
            .I(N__25544));
    LocalMux I__5468 (
            .O(N__25547),
            .I(N__25539));
    Sp12to4 I__5467 (
            .O(N__25544),
            .I(N__25536));
    InMux I__5466 (
            .O(N__25543),
            .I(N__25531));
    InMux I__5465 (
            .O(N__25542),
            .I(N__25531));
    Odrv12 I__5464 (
            .O(N__25539),
            .I(\c0.data_in_field_120 ));
    Odrv12 I__5463 (
            .O(N__25536),
            .I(\c0.data_in_field_120 ));
    LocalMux I__5462 (
            .O(N__25531),
            .I(\c0.data_in_field_120 ));
    InMux I__5461 (
            .O(N__25524),
            .I(N__25521));
    LocalMux I__5460 (
            .O(N__25521),
            .I(N__25518));
    Span4Mux_h I__5459 (
            .O(N__25518),
            .I(N__25514));
    InMux I__5458 (
            .O(N__25517),
            .I(N__25511));
    Span4Mux_h I__5457 (
            .O(N__25514),
            .I(N__25508));
    LocalMux I__5456 (
            .O(N__25511),
            .I(N__25505));
    Odrv4 I__5455 (
            .O(N__25508),
            .I(\c0.n2107 ));
    Odrv12 I__5454 (
            .O(N__25505),
            .I(\c0.n2107 ));
    InMux I__5453 (
            .O(N__25500),
            .I(N__25497));
    LocalMux I__5452 (
            .O(N__25497),
            .I(N__25493));
    CascadeMux I__5451 (
            .O(N__25496),
            .I(N__25490));
    Span4Mux_h I__5450 (
            .O(N__25493),
            .I(N__25487));
    InMux I__5449 (
            .O(N__25490),
            .I(N__25484));
    Odrv4 I__5448 (
            .O(N__25487),
            .I(rx_data_2));
    LocalMux I__5447 (
            .O(N__25484),
            .I(rx_data_2));
    InMux I__5446 (
            .O(N__25479),
            .I(N__25476));
    LocalMux I__5445 (
            .O(N__25476),
            .I(N__25473));
    Span4Mux_v I__5444 (
            .O(N__25473),
            .I(N__25470));
    Span4Mux_h I__5443 (
            .O(N__25470),
            .I(N__25467));
    Odrv4 I__5442 (
            .O(N__25467),
            .I(\c0.n6201 ));
    InMux I__5441 (
            .O(N__25464),
            .I(N__25459));
    InMux I__5440 (
            .O(N__25463),
            .I(N__25456));
    InMux I__5439 (
            .O(N__25462),
            .I(N__25451));
    LocalMux I__5438 (
            .O(N__25459),
            .I(N__25448));
    LocalMux I__5437 (
            .O(N__25456),
            .I(N__25445));
    CascadeMux I__5436 (
            .O(N__25455),
            .I(N__25442));
    CascadeMux I__5435 (
            .O(N__25454),
            .I(N__25438));
    LocalMux I__5434 (
            .O(N__25451),
            .I(N__25435));
    Span4Mux_v I__5433 (
            .O(N__25448),
            .I(N__25430));
    Span4Mux_h I__5432 (
            .O(N__25445),
            .I(N__25430));
    InMux I__5431 (
            .O(N__25442),
            .I(N__25427));
    InMux I__5430 (
            .O(N__25441),
            .I(N__25422));
    InMux I__5429 (
            .O(N__25438),
            .I(N__25422));
    Odrv4 I__5428 (
            .O(N__25435),
            .I(\c0.data_in_field_101 ));
    Odrv4 I__5427 (
            .O(N__25430),
            .I(\c0.data_in_field_101 ));
    LocalMux I__5426 (
            .O(N__25427),
            .I(\c0.data_in_field_101 ));
    LocalMux I__5425 (
            .O(N__25422),
            .I(\c0.data_in_field_101 ));
    CascadeMux I__5424 (
            .O(N__25413),
            .I(N__25410));
    InMux I__5423 (
            .O(N__25410),
            .I(N__25399));
    InMux I__5422 (
            .O(N__25409),
            .I(N__25396));
    CascadeMux I__5421 (
            .O(N__25408),
            .I(N__25393));
    CascadeMux I__5420 (
            .O(N__25407),
            .I(N__25387));
    InMux I__5419 (
            .O(N__25406),
            .I(N__25383));
    InMux I__5418 (
            .O(N__25405),
            .I(N__25376));
    InMux I__5417 (
            .O(N__25404),
            .I(N__25376));
    InMux I__5416 (
            .O(N__25403),
            .I(N__25373));
    InMux I__5415 (
            .O(N__25402),
            .I(N__25369));
    LocalMux I__5414 (
            .O(N__25399),
            .I(N__25364));
    LocalMux I__5413 (
            .O(N__25396),
            .I(N__25364));
    InMux I__5412 (
            .O(N__25393),
            .I(N__25361));
    InMux I__5411 (
            .O(N__25392),
            .I(N__25358));
    InMux I__5410 (
            .O(N__25391),
            .I(N__25355));
    InMux I__5409 (
            .O(N__25390),
            .I(N__25350));
    InMux I__5408 (
            .O(N__25387),
            .I(N__25350));
    InMux I__5407 (
            .O(N__25386),
            .I(N__25347));
    LocalMux I__5406 (
            .O(N__25383),
            .I(N__25344));
    InMux I__5405 (
            .O(N__25382),
            .I(N__25339));
    InMux I__5404 (
            .O(N__25381),
            .I(N__25339));
    LocalMux I__5403 (
            .O(N__25376),
            .I(N__25336));
    LocalMux I__5402 (
            .O(N__25373),
            .I(N__25333));
    InMux I__5401 (
            .O(N__25372),
            .I(N__25330));
    LocalMux I__5400 (
            .O(N__25369),
            .I(N__25327));
    Span4Mux_h I__5399 (
            .O(N__25364),
            .I(N__25324));
    LocalMux I__5398 (
            .O(N__25361),
            .I(N__25321));
    LocalMux I__5397 (
            .O(N__25358),
            .I(N__25316));
    LocalMux I__5396 (
            .O(N__25355),
            .I(N__25316));
    LocalMux I__5395 (
            .O(N__25350),
            .I(N__25307));
    LocalMux I__5394 (
            .O(N__25347),
            .I(N__25307));
    Span4Mux_v I__5393 (
            .O(N__25344),
            .I(N__25307));
    LocalMux I__5392 (
            .O(N__25339),
            .I(N__25307));
    Span4Mux_v I__5391 (
            .O(N__25336),
            .I(N__25298));
    Span4Mux_s3_h I__5390 (
            .O(N__25333),
            .I(N__25298));
    LocalMux I__5389 (
            .O(N__25330),
            .I(N__25298));
    Span4Mux_v I__5388 (
            .O(N__25327),
            .I(N__25295));
    Span4Mux_v I__5387 (
            .O(N__25324),
            .I(N__25292));
    Span4Mux_h I__5386 (
            .O(N__25321),
            .I(N__25285));
    Span4Mux_s1_h I__5385 (
            .O(N__25316),
            .I(N__25285));
    Span4Mux_v I__5384 (
            .O(N__25307),
            .I(N__25285));
    InMux I__5383 (
            .O(N__25306),
            .I(N__25282));
    InMux I__5382 (
            .O(N__25305),
            .I(N__25279));
    Span4Mux_v I__5381 (
            .O(N__25298),
            .I(N__25276));
    Span4Mux_h I__5380 (
            .O(N__25295),
            .I(N__25269));
    Span4Mux_h I__5379 (
            .O(N__25292),
            .I(N__25269));
    Span4Mux_v I__5378 (
            .O(N__25285),
            .I(N__25269));
    LocalMux I__5377 (
            .O(N__25282),
            .I(\c0.byte_transmit_counter2_3 ));
    LocalMux I__5376 (
            .O(N__25279),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__5375 (
            .O(N__25276),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__5374 (
            .O(N__25269),
            .I(\c0.byte_transmit_counter2_3 ));
    InMux I__5373 (
            .O(N__25260),
            .I(N__25253));
    InMux I__5372 (
            .O(N__25259),
            .I(N__25249));
    InMux I__5371 (
            .O(N__25258),
            .I(N__25244));
    InMux I__5370 (
            .O(N__25257),
            .I(N__25239));
    InMux I__5369 (
            .O(N__25256),
            .I(N__25239));
    LocalMux I__5368 (
            .O(N__25253),
            .I(N__25235));
    InMux I__5367 (
            .O(N__25252),
            .I(N__25232));
    LocalMux I__5366 (
            .O(N__25249),
            .I(N__25228));
    InMux I__5365 (
            .O(N__25248),
            .I(N__25225));
    InMux I__5364 (
            .O(N__25247),
            .I(N__25222));
    LocalMux I__5363 (
            .O(N__25244),
            .I(N__25219));
    LocalMux I__5362 (
            .O(N__25239),
            .I(N__25216));
    InMux I__5361 (
            .O(N__25238),
            .I(N__25213));
    Span4Mux_v I__5360 (
            .O(N__25235),
            .I(N__25210));
    LocalMux I__5359 (
            .O(N__25232),
            .I(N__25207));
    InMux I__5358 (
            .O(N__25231),
            .I(N__25204));
    Span4Mux_h I__5357 (
            .O(N__25228),
            .I(N__25201));
    LocalMux I__5356 (
            .O(N__25225),
            .I(N__25198));
    LocalMux I__5355 (
            .O(N__25222),
            .I(N__25195));
    Span4Mux_v I__5354 (
            .O(N__25219),
            .I(N__25190));
    Span4Mux_s2_h I__5353 (
            .O(N__25216),
            .I(N__25190));
    LocalMux I__5352 (
            .O(N__25213),
            .I(N__25185));
    Span4Mux_v I__5351 (
            .O(N__25210),
            .I(N__25185));
    Span4Mux_h I__5350 (
            .O(N__25207),
            .I(N__25182));
    LocalMux I__5349 (
            .O(N__25204),
            .I(N__25173));
    Span4Mux_h I__5348 (
            .O(N__25201),
            .I(N__25173));
    Span4Mux_v I__5347 (
            .O(N__25198),
            .I(N__25173));
    Span4Mux_s3_h I__5346 (
            .O(N__25195),
            .I(N__25173));
    Span4Mux_v I__5345 (
            .O(N__25190),
            .I(N__25170));
    Odrv4 I__5344 (
            .O(N__25185),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__5343 (
            .O(N__25182),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__5342 (
            .O(N__25173),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__5341 (
            .O(N__25170),
            .I(\c0.byte_transmit_counter2_2 ));
    CascadeMux I__5340 (
            .O(N__25161),
            .I(\c0.n5716_cascade_ ));
    InMux I__5339 (
            .O(N__25158),
            .I(N__25155));
    LocalMux I__5338 (
            .O(N__25155),
            .I(\c0.n6195 ));
    InMux I__5337 (
            .O(N__25152),
            .I(N__25149));
    LocalMux I__5336 (
            .O(N__25149),
            .I(N__25145));
    InMux I__5335 (
            .O(N__25148),
            .I(N__25141));
    Span4Mux_v I__5334 (
            .O(N__25145),
            .I(N__25138));
    InMux I__5333 (
            .O(N__25144),
            .I(N__25135));
    LocalMux I__5332 (
            .O(N__25141),
            .I(N__25131));
    Span4Mux_h I__5331 (
            .O(N__25138),
            .I(N__25126));
    LocalMux I__5330 (
            .O(N__25135),
            .I(N__25126));
    InMux I__5329 (
            .O(N__25134),
            .I(N__25123));
    Span4Mux_v I__5328 (
            .O(N__25131),
            .I(N__25118));
    Span4Mux_h I__5327 (
            .O(N__25126),
            .I(N__25118));
    LocalMux I__5326 (
            .O(N__25123),
            .I(\c0.data_in_field_85 ));
    Odrv4 I__5325 (
            .O(N__25118),
            .I(\c0.data_in_field_85 ));
    InMux I__5324 (
            .O(N__25113),
            .I(N__25109));
    InMux I__5323 (
            .O(N__25112),
            .I(N__25106));
    LocalMux I__5322 (
            .O(N__25109),
            .I(N__25101));
    LocalMux I__5321 (
            .O(N__25106),
            .I(N__25098));
    InMux I__5320 (
            .O(N__25105),
            .I(N__25095));
    InMux I__5319 (
            .O(N__25104),
            .I(N__25091));
    Span4Mux_h I__5318 (
            .O(N__25101),
            .I(N__25088));
    Span12Mux_s3_h I__5317 (
            .O(N__25098),
            .I(N__25085));
    LocalMux I__5316 (
            .O(N__25095),
            .I(N__25082));
    InMux I__5315 (
            .O(N__25094),
            .I(N__25079));
    LocalMux I__5314 (
            .O(N__25091),
            .I(\c0.data_in_field_93 ));
    Odrv4 I__5313 (
            .O(N__25088),
            .I(\c0.data_in_field_93 ));
    Odrv12 I__5312 (
            .O(N__25085),
            .I(\c0.data_in_field_93 ));
    Odrv4 I__5311 (
            .O(N__25082),
            .I(\c0.data_in_field_93 ));
    LocalMux I__5310 (
            .O(N__25079),
            .I(\c0.data_in_field_93 ));
    InMux I__5309 (
            .O(N__25068),
            .I(N__25065));
    LocalMux I__5308 (
            .O(N__25065),
            .I(\c0.n37 ));
    InMux I__5307 (
            .O(N__25062),
            .I(N__25059));
    LocalMux I__5306 (
            .O(N__25059),
            .I(N__25055));
    InMux I__5305 (
            .O(N__25058),
            .I(N__25052));
    Span4Mux_h I__5304 (
            .O(N__25055),
            .I(N__25049));
    LocalMux I__5303 (
            .O(N__25052),
            .I(N__25046));
    Span4Mux_v I__5302 (
            .O(N__25049),
            .I(N__25039));
    Span4Mux_v I__5301 (
            .O(N__25046),
            .I(N__25039));
    InMux I__5300 (
            .O(N__25045),
            .I(N__25036));
    InMux I__5299 (
            .O(N__25044),
            .I(N__25033));
    Odrv4 I__5298 (
            .O(N__25039),
            .I(data_in_1_5));
    LocalMux I__5297 (
            .O(N__25036),
            .I(data_in_1_5));
    LocalMux I__5296 (
            .O(N__25033),
            .I(data_in_1_5));
    CascadeMux I__5295 (
            .O(N__25026),
            .I(N__25022));
    InMux I__5294 (
            .O(N__25025),
            .I(N__25019));
    InMux I__5293 (
            .O(N__25022),
            .I(N__25014));
    LocalMux I__5292 (
            .O(N__25019),
            .I(N__25011));
    InMux I__5291 (
            .O(N__25018),
            .I(N__25006));
    InMux I__5290 (
            .O(N__25017),
            .I(N__25006));
    LocalMux I__5289 (
            .O(N__25014),
            .I(\c0.data_in_field_13 ));
    Odrv4 I__5288 (
            .O(N__25011),
            .I(\c0.data_in_field_13 ));
    LocalMux I__5287 (
            .O(N__25006),
            .I(\c0.data_in_field_13 ));
    CascadeMux I__5286 (
            .O(N__24999),
            .I(N__24996));
    InMux I__5285 (
            .O(N__24996),
            .I(N__24993));
    LocalMux I__5284 (
            .O(N__24993),
            .I(\c0.n6_adj_1939 ));
    CascadeMux I__5283 (
            .O(N__24990),
            .I(N__24987));
    InMux I__5282 (
            .O(N__24987),
            .I(N__24984));
    LocalMux I__5281 (
            .O(N__24984),
            .I(N__24979));
    InMux I__5280 (
            .O(N__24983),
            .I(N__24974));
    InMux I__5279 (
            .O(N__24982),
            .I(N__24974));
    Odrv4 I__5278 (
            .O(N__24979),
            .I(data_in_12_4));
    LocalMux I__5277 (
            .O(N__24974),
            .I(data_in_12_4));
    CascadeMux I__5276 (
            .O(N__24969),
            .I(N__24966));
    InMux I__5275 (
            .O(N__24966),
            .I(N__24963));
    LocalMux I__5274 (
            .O(N__24963),
            .I(N__24960));
    Span4Mux_h I__5273 (
            .O(N__24960),
            .I(N__24955));
    InMux I__5272 (
            .O(N__24959),
            .I(N__24952));
    InMux I__5271 (
            .O(N__24958),
            .I(N__24949));
    Odrv4 I__5270 (
            .O(N__24955),
            .I(data_in_11_4));
    LocalMux I__5269 (
            .O(N__24952),
            .I(data_in_11_4));
    LocalMux I__5268 (
            .O(N__24949),
            .I(data_in_11_4));
    InMux I__5267 (
            .O(N__24942),
            .I(N__24939));
    LocalMux I__5266 (
            .O(N__24939),
            .I(N__24936));
    Span4Mux_h I__5265 (
            .O(N__24936),
            .I(N__24933));
    Span4Mux_h I__5264 (
            .O(N__24933),
            .I(N__24930));
    Odrv4 I__5263 (
            .O(N__24930),
            .I(\c0.n2089 ));
    InMux I__5262 (
            .O(N__24927),
            .I(N__24924));
    LocalMux I__5261 (
            .O(N__24924),
            .I(N__24921));
    Odrv12 I__5260 (
            .O(N__24921),
            .I(\c0.n2074 ));
    InMux I__5259 (
            .O(N__24918),
            .I(N__24915));
    LocalMux I__5258 (
            .O(N__24915),
            .I(N__24911));
    InMux I__5257 (
            .O(N__24914),
            .I(N__24908));
    Span12Mux_s6_h I__5256 (
            .O(N__24911),
            .I(N__24905));
    LocalMux I__5255 (
            .O(N__24908),
            .I(N__24902));
    Odrv12 I__5254 (
            .O(N__24905),
            .I(\c0.n5581 ));
    Odrv4 I__5253 (
            .O(N__24902),
            .I(\c0.n5581 ));
    InMux I__5252 (
            .O(N__24897),
            .I(N__24894));
    LocalMux I__5251 (
            .O(N__24894),
            .I(N__24891));
    Span4Mux_v I__5250 (
            .O(N__24891),
            .I(N__24887));
    InMux I__5249 (
            .O(N__24890),
            .I(N__24883));
    Span4Mux_h I__5248 (
            .O(N__24887),
            .I(N__24880));
    InMux I__5247 (
            .O(N__24886),
            .I(N__24877));
    LocalMux I__5246 (
            .O(N__24883),
            .I(\c0.data_in_field_44 ));
    Odrv4 I__5245 (
            .O(N__24880),
            .I(\c0.data_in_field_44 ));
    LocalMux I__5244 (
            .O(N__24877),
            .I(\c0.data_in_field_44 ));
    InMux I__5243 (
            .O(N__24870),
            .I(N__24865));
    InMux I__5242 (
            .O(N__24869),
            .I(N__24862));
    InMux I__5241 (
            .O(N__24868),
            .I(N__24858));
    LocalMux I__5240 (
            .O(N__24865),
            .I(N__24855));
    LocalMux I__5239 (
            .O(N__24862),
            .I(N__24852));
    InMux I__5238 (
            .O(N__24861),
            .I(N__24849));
    LocalMux I__5237 (
            .O(N__24858),
            .I(N__24846));
    Span4Mux_h I__5236 (
            .O(N__24855),
            .I(N__24842));
    Span4Mux_v I__5235 (
            .O(N__24852),
            .I(N__24839));
    LocalMux I__5234 (
            .O(N__24849),
            .I(N__24836));
    Span4Mux_v I__5233 (
            .O(N__24846),
            .I(N__24833));
    InMux I__5232 (
            .O(N__24845),
            .I(N__24829));
    Span4Mux_h I__5231 (
            .O(N__24842),
            .I(N__24826));
    Span4Mux_v I__5230 (
            .O(N__24839),
            .I(N__24819));
    Span4Mux_v I__5229 (
            .O(N__24836),
            .I(N__24819));
    Span4Mux_h I__5228 (
            .O(N__24833),
            .I(N__24819));
    InMux I__5227 (
            .O(N__24832),
            .I(N__24816));
    LocalMux I__5226 (
            .O(N__24829),
            .I(\c0.data_in_field_100 ));
    Odrv4 I__5225 (
            .O(N__24826),
            .I(\c0.data_in_field_100 ));
    Odrv4 I__5224 (
            .O(N__24819),
            .I(\c0.data_in_field_100 ));
    LocalMux I__5223 (
            .O(N__24816),
            .I(\c0.data_in_field_100 ));
    InMux I__5222 (
            .O(N__24807),
            .I(N__24803));
    InMux I__5221 (
            .O(N__24806),
            .I(N__24799));
    LocalMux I__5220 (
            .O(N__24803),
            .I(N__24796));
    InMux I__5219 (
            .O(N__24802),
            .I(N__24793));
    LocalMux I__5218 (
            .O(N__24799),
            .I(N__24789));
    Span4Mux_h I__5217 (
            .O(N__24796),
            .I(N__24786));
    LocalMux I__5216 (
            .O(N__24793),
            .I(N__24783));
    InMux I__5215 (
            .O(N__24792),
            .I(N__24778));
    Span12Mux_s9_v I__5214 (
            .O(N__24789),
            .I(N__24775));
    Span4Mux_h I__5213 (
            .O(N__24786),
            .I(N__24772));
    Span4Mux_v I__5212 (
            .O(N__24783),
            .I(N__24769));
    InMux I__5211 (
            .O(N__24782),
            .I(N__24766));
    InMux I__5210 (
            .O(N__24781),
            .I(N__24763));
    LocalMux I__5209 (
            .O(N__24778),
            .I(\c0.data_in_field_50 ));
    Odrv12 I__5208 (
            .O(N__24775),
            .I(\c0.data_in_field_50 ));
    Odrv4 I__5207 (
            .O(N__24772),
            .I(\c0.data_in_field_50 ));
    Odrv4 I__5206 (
            .O(N__24769),
            .I(\c0.data_in_field_50 ));
    LocalMux I__5205 (
            .O(N__24766),
            .I(\c0.data_in_field_50 ));
    LocalMux I__5204 (
            .O(N__24763),
            .I(\c0.data_in_field_50 ));
    InMux I__5203 (
            .O(N__24750),
            .I(N__24747));
    LocalMux I__5202 (
            .O(N__24747),
            .I(N__24743));
    InMux I__5201 (
            .O(N__24746),
            .I(N__24740));
    Span4Mux_h I__5200 (
            .O(N__24743),
            .I(N__24737));
    LocalMux I__5199 (
            .O(N__24740),
            .I(\c0.n2053 ));
    Odrv4 I__5198 (
            .O(N__24737),
            .I(\c0.n2053 ));
    CascadeMux I__5197 (
            .O(N__24732),
            .I(N__24729));
    InMux I__5196 (
            .O(N__24729),
            .I(N__24726));
    LocalMux I__5195 (
            .O(N__24726),
            .I(N__24723));
    Span4Mux_h I__5194 (
            .O(N__24723),
            .I(N__24720));
    Span4Mux_h I__5193 (
            .O(N__24720),
            .I(N__24717));
    Odrv4 I__5192 (
            .O(N__24717),
            .I(\c0.n2101 ));
    InMux I__5191 (
            .O(N__24714),
            .I(N__24711));
    LocalMux I__5190 (
            .O(N__24711),
            .I(N__24708));
    Span4Mux_v I__5189 (
            .O(N__24708),
            .I(N__24704));
    InMux I__5188 (
            .O(N__24707),
            .I(N__24701));
    Span4Mux_h I__5187 (
            .O(N__24704),
            .I(N__24696));
    LocalMux I__5186 (
            .O(N__24701),
            .I(N__24696));
    Odrv4 I__5185 (
            .O(N__24696),
            .I(\c0.n2134 ));
    CascadeMux I__5184 (
            .O(N__24693),
            .I(\c0.n31_adj_1900_cascade_ ));
    InMux I__5183 (
            .O(N__24690),
            .I(N__24687));
    LocalMux I__5182 (
            .O(N__24687),
            .I(\c0.n35 ));
    CascadeMux I__5181 (
            .O(N__24684),
            .I(N__24681));
    InMux I__5180 (
            .O(N__24681),
            .I(N__24677));
    CascadeMux I__5179 (
            .O(N__24680),
            .I(N__24674));
    LocalMux I__5178 (
            .O(N__24677),
            .I(N__24671));
    InMux I__5177 (
            .O(N__24674),
            .I(N__24667));
    Span4Mux_h I__5176 (
            .O(N__24671),
            .I(N__24664));
    InMux I__5175 (
            .O(N__24670),
            .I(N__24661));
    LocalMux I__5174 (
            .O(N__24667),
            .I(N__24658));
    Odrv4 I__5173 (
            .O(N__24664),
            .I(data_in_0_2));
    LocalMux I__5172 (
            .O(N__24661),
            .I(data_in_0_2));
    Odrv4 I__5171 (
            .O(N__24658),
            .I(data_in_0_2));
    InMux I__5170 (
            .O(N__24651),
            .I(N__24648));
    LocalMux I__5169 (
            .O(N__24648),
            .I(\c0.n14 ));
    InMux I__5168 (
            .O(N__24645),
            .I(N__24642));
    LocalMux I__5167 (
            .O(N__24642),
            .I(\c0.n5582 ));
    CascadeMux I__5166 (
            .O(N__24639),
            .I(N__24636));
    InMux I__5165 (
            .O(N__24636),
            .I(N__24633));
    LocalMux I__5164 (
            .O(N__24633),
            .I(N__24630));
    Odrv4 I__5163 (
            .O(N__24630),
            .I(\c0.n13_adj_1899 ));
    InMux I__5162 (
            .O(N__24627),
            .I(N__24624));
    LocalMux I__5161 (
            .O(N__24624),
            .I(\c0.n17_adj_1902 ));
    InMux I__5160 (
            .O(N__24621),
            .I(N__24618));
    LocalMux I__5159 (
            .O(N__24618),
            .I(N__24615));
    Odrv12 I__5158 (
            .O(N__24615),
            .I(\c0.n25_adj_1907 ));
    InMux I__5157 (
            .O(N__24612),
            .I(N__24609));
    LocalMux I__5156 (
            .O(N__24609),
            .I(\c0.n4_adj_1920 ));
    InMux I__5155 (
            .O(N__24606),
            .I(N__24600));
    InMux I__5154 (
            .O(N__24605),
            .I(N__24597));
    InMux I__5153 (
            .O(N__24604),
            .I(N__24594));
    CascadeMux I__5152 (
            .O(N__24603),
            .I(N__24591));
    LocalMux I__5151 (
            .O(N__24600),
            .I(N__24588));
    LocalMux I__5150 (
            .O(N__24597),
            .I(N__24585));
    LocalMux I__5149 (
            .O(N__24594),
            .I(N__24582));
    InMux I__5148 (
            .O(N__24591),
            .I(N__24578));
    Span4Mux_h I__5147 (
            .O(N__24588),
            .I(N__24575));
    Span12Mux_v I__5146 (
            .O(N__24585),
            .I(N__24572));
    Span4Mux_h I__5145 (
            .O(N__24582),
            .I(N__24569));
    InMux I__5144 (
            .O(N__24581),
            .I(N__24566));
    LocalMux I__5143 (
            .O(N__24578),
            .I(\c0.data_in_field_122 ));
    Odrv4 I__5142 (
            .O(N__24575),
            .I(\c0.data_in_field_122 ));
    Odrv12 I__5141 (
            .O(N__24572),
            .I(\c0.data_in_field_122 ));
    Odrv4 I__5140 (
            .O(N__24569),
            .I(\c0.data_in_field_122 ));
    LocalMux I__5139 (
            .O(N__24566),
            .I(\c0.data_in_field_122 ));
    InMux I__5138 (
            .O(N__24555),
            .I(N__24552));
    LocalMux I__5137 (
            .O(N__24552),
            .I(N__24549));
    Span4Mux_v I__5136 (
            .O(N__24549),
            .I(N__24546));
    Odrv4 I__5135 (
            .O(N__24546),
            .I(\c0.n5593 ));
    CascadeMux I__5134 (
            .O(N__24543),
            .I(N__24540));
    InMux I__5133 (
            .O(N__24540),
            .I(N__24537));
    LocalMux I__5132 (
            .O(N__24537),
            .I(N__24533));
    InMux I__5131 (
            .O(N__24536),
            .I(N__24530));
    Span4Mux_v I__5130 (
            .O(N__24533),
            .I(N__24522));
    LocalMux I__5129 (
            .O(N__24530),
            .I(N__24522));
    CascadeMux I__5128 (
            .O(N__24529),
            .I(N__24518));
    InMux I__5127 (
            .O(N__24528),
            .I(N__24515));
    InMux I__5126 (
            .O(N__24527),
            .I(N__24512));
    Span4Mux_h I__5125 (
            .O(N__24522),
            .I(N__24509));
    CascadeMux I__5124 (
            .O(N__24521),
            .I(N__24506));
    InMux I__5123 (
            .O(N__24518),
            .I(N__24503));
    LocalMux I__5122 (
            .O(N__24515),
            .I(N__24500));
    LocalMux I__5121 (
            .O(N__24512),
            .I(N__24497));
    Span4Mux_h I__5120 (
            .O(N__24509),
            .I(N__24494));
    InMux I__5119 (
            .O(N__24506),
            .I(N__24491));
    LocalMux I__5118 (
            .O(N__24503),
            .I(\c0.data_in_field_62 ));
    Odrv12 I__5117 (
            .O(N__24500),
            .I(\c0.data_in_field_62 ));
    Odrv4 I__5116 (
            .O(N__24497),
            .I(\c0.data_in_field_62 ));
    Odrv4 I__5115 (
            .O(N__24494),
            .I(\c0.data_in_field_62 ));
    LocalMux I__5114 (
            .O(N__24491),
            .I(\c0.data_in_field_62 ));
    CascadeMux I__5113 (
            .O(N__24480),
            .I(\c0.n5593_cascade_ ));
    InMux I__5112 (
            .O(N__24477),
            .I(N__24474));
    LocalMux I__5111 (
            .O(N__24474),
            .I(\c0.n5430 ));
    InMux I__5110 (
            .O(N__24471),
            .I(N__24468));
    LocalMux I__5109 (
            .O(N__24468),
            .I(\c0.n33 ));
    CascadeMux I__5108 (
            .O(N__24465),
            .I(\c0.n5430_cascade_ ));
    InMux I__5107 (
            .O(N__24462),
            .I(N__24459));
    LocalMux I__5106 (
            .O(N__24459),
            .I(N__24456));
    Odrv12 I__5105 (
            .O(N__24456),
            .I(\c0.n28_adj_1955 ));
    InMux I__5104 (
            .O(N__24453),
            .I(N__24450));
    LocalMux I__5103 (
            .O(N__24450),
            .I(\c0.n5384 ));
    InMux I__5102 (
            .O(N__24447),
            .I(N__24444));
    LocalMux I__5101 (
            .O(N__24444),
            .I(N__24441));
    Span4Mux_h I__5100 (
            .O(N__24441),
            .I(N__24438));
    Span4Mux_h I__5099 (
            .O(N__24438),
            .I(N__24434));
    InMux I__5098 (
            .O(N__24437),
            .I(N__24431));
    Odrv4 I__5097 (
            .O(N__24434),
            .I(\c0.n5476 ));
    LocalMux I__5096 (
            .O(N__24431),
            .I(\c0.n5476 ));
    CascadeMux I__5095 (
            .O(N__24426),
            .I(N__24423));
    InMux I__5094 (
            .O(N__24423),
            .I(N__24420));
    LocalMux I__5093 (
            .O(N__24420),
            .I(N__24417));
    Span4Mux_h I__5092 (
            .O(N__24417),
            .I(N__24414));
    Odrv4 I__5091 (
            .O(N__24414),
            .I(\c0.n5427 ));
    InMux I__5090 (
            .O(N__24411),
            .I(N__24408));
    LocalMux I__5089 (
            .O(N__24408),
            .I(N__24405));
    Span4Mux_h I__5088 (
            .O(N__24405),
            .I(N__24402));
    Span4Mux_h I__5087 (
            .O(N__24402),
            .I(N__24398));
    InMux I__5086 (
            .O(N__24401),
            .I(N__24395));
    Odrv4 I__5085 (
            .O(N__24398),
            .I(\c0.n5521 ));
    LocalMux I__5084 (
            .O(N__24395),
            .I(\c0.n5521 ));
    InMux I__5083 (
            .O(N__24390),
            .I(N__24387));
    LocalMux I__5082 (
            .O(N__24387),
            .I(\c0.n24_adj_1885 ));
    InMux I__5081 (
            .O(N__24384),
            .I(N__24381));
    LocalMux I__5080 (
            .O(N__24381),
            .I(N__24377));
    InMux I__5079 (
            .O(N__24380),
            .I(N__24374));
    Span4Mux_h I__5078 (
            .O(N__24377),
            .I(N__24369));
    LocalMux I__5077 (
            .O(N__24374),
            .I(N__24369));
    Odrv4 I__5076 (
            .O(N__24369),
            .I(\c0.n1866 ));
    InMux I__5075 (
            .O(N__24366),
            .I(N__24362));
    InMux I__5074 (
            .O(N__24365),
            .I(N__24359));
    LocalMux I__5073 (
            .O(N__24362),
            .I(N__24356));
    LocalMux I__5072 (
            .O(N__24359),
            .I(N__24352));
    Span4Mux_v I__5071 (
            .O(N__24356),
            .I(N__24349));
    CascadeMux I__5070 (
            .O(N__24355),
            .I(N__24346));
    Span4Mux_v I__5069 (
            .O(N__24352),
            .I(N__24339));
    Span4Mux_h I__5068 (
            .O(N__24349),
            .I(N__24339));
    InMux I__5067 (
            .O(N__24346),
            .I(N__24336));
    InMux I__5066 (
            .O(N__24345),
            .I(N__24331));
    InMux I__5065 (
            .O(N__24344),
            .I(N__24331));
    Odrv4 I__5064 (
            .O(N__24339),
            .I(\c0.data_in_field_113 ));
    LocalMux I__5063 (
            .O(N__24336),
            .I(\c0.data_in_field_113 ));
    LocalMux I__5062 (
            .O(N__24331),
            .I(\c0.data_in_field_113 ));
    InMux I__5061 (
            .O(N__24324),
            .I(N__24321));
    LocalMux I__5060 (
            .O(N__24321),
            .I(N__24318));
    Span4Mux_v I__5059 (
            .O(N__24318),
            .I(N__24313));
    InMux I__5058 (
            .O(N__24317),
            .I(N__24310));
    InMux I__5057 (
            .O(N__24316),
            .I(N__24306));
    Span4Mux_h I__5056 (
            .O(N__24313),
            .I(N__24303));
    LocalMux I__5055 (
            .O(N__24310),
            .I(N__24300));
    InMux I__5054 (
            .O(N__24309),
            .I(N__24296));
    LocalMux I__5053 (
            .O(N__24306),
            .I(N__24293));
    Span4Mux_h I__5052 (
            .O(N__24303),
            .I(N__24290));
    Span4Mux_h I__5051 (
            .O(N__24300),
            .I(N__24287));
    InMux I__5050 (
            .O(N__24299),
            .I(N__24284));
    LocalMux I__5049 (
            .O(N__24296),
            .I(\c0.data_in_field_57 ));
    Odrv12 I__5048 (
            .O(N__24293),
            .I(\c0.data_in_field_57 ));
    Odrv4 I__5047 (
            .O(N__24290),
            .I(\c0.data_in_field_57 ));
    Odrv4 I__5046 (
            .O(N__24287),
            .I(\c0.data_in_field_57 ));
    LocalMux I__5045 (
            .O(N__24284),
            .I(\c0.data_in_field_57 ));
    CascadeMux I__5044 (
            .O(N__24273),
            .I(\c0.n10_cascade_ ));
    InMux I__5043 (
            .O(N__24270),
            .I(N__24267));
    LocalMux I__5042 (
            .O(N__24267),
            .I(N__24264));
    Span4Mux_v I__5041 (
            .O(N__24264),
            .I(N__24260));
    InMux I__5040 (
            .O(N__24263),
            .I(N__24257));
    Span4Mux_h I__5039 (
            .O(N__24260),
            .I(N__24254));
    LocalMux I__5038 (
            .O(N__24257),
            .I(N__24251));
    Odrv4 I__5037 (
            .O(N__24254),
            .I(\c0.n5466 ));
    Odrv12 I__5036 (
            .O(N__24251),
            .I(\c0.n5466 ));
    InMux I__5035 (
            .O(N__24246),
            .I(N__24243));
    LocalMux I__5034 (
            .O(N__24243),
            .I(\c0.n5519 ));
    InMux I__5033 (
            .O(N__24240),
            .I(N__24236));
    InMux I__5032 (
            .O(N__24239),
            .I(N__24233));
    LocalMux I__5031 (
            .O(N__24236),
            .I(N__24230));
    LocalMux I__5030 (
            .O(N__24233),
            .I(N__24227));
    Span4Mux_v I__5029 (
            .O(N__24230),
            .I(N__24223));
    Span4Mux_h I__5028 (
            .O(N__24227),
            .I(N__24220));
    InMux I__5027 (
            .O(N__24226),
            .I(N__24217));
    Odrv4 I__5026 (
            .O(N__24223),
            .I(data_in_7_6));
    Odrv4 I__5025 (
            .O(N__24220),
            .I(data_in_7_6));
    LocalMux I__5024 (
            .O(N__24217),
            .I(data_in_7_6));
    InMux I__5023 (
            .O(N__24210),
            .I(N__24206));
    InMux I__5022 (
            .O(N__24209),
            .I(N__24203));
    LocalMux I__5021 (
            .O(N__24206),
            .I(N__24199));
    LocalMux I__5020 (
            .O(N__24203),
            .I(N__24196));
    InMux I__5019 (
            .O(N__24202),
            .I(N__24193));
    Span4Mux_h I__5018 (
            .O(N__24199),
            .I(N__24190));
    Span4Mux_h I__5017 (
            .O(N__24196),
            .I(N__24187));
    LocalMux I__5016 (
            .O(N__24193),
            .I(data_in_6_6));
    Odrv4 I__5015 (
            .O(N__24190),
            .I(data_in_6_6));
    Odrv4 I__5014 (
            .O(N__24187),
            .I(data_in_6_6));
    CascadeMux I__5013 (
            .O(N__24180),
            .I(N__24177));
    InMux I__5012 (
            .O(N__24177),
            .I(N__24173));
    InMux I__5011 (
            .O(N__24176),
            .I(N__24170));
    LocalMux I__5010 (
            .O(N__24173),
            .I(N__24165));
    LocalMux I__5009 (
            .O(N__24170),
            .I(N__24162));
    InMux I__5008 (
            .O(N__24169),
            .I(N__24159));
    InMux I__5007 (
            .O(N__24168),
            .I(N__24156));
    Span12Mux_v I__5006 (
            .O(N__24165),
            .I(N__24153));
    Odrv12 I__5005 (
            .O(N__24162),
            .I(data_in_18_0));
    LocalMux I__5004 (
            .O(N__24159),
            .I(data_in_18_0));
    LocalMux I__5003 (
            .O(N__24156),
            .I(data_in_18_0));
    Odrv12 I__5002 (
            .O(N__24153),
            .I(data_in_18_0));
    InMux I__5001 (
            .O(N__24144),
            .I(N__24141));
    LocalMux I__5000 (
            .O(N__24141),
            .I(N__24138));
    Odrv12 I__4999 (
            .O(N__24138),
            .I(\c0.n5548 ));
    InMux I__4998 (
            .O(N__24135),
            .I(N__24131));
    InMux I__4997 (
            .O(N__24134),
            .I(N__24128));
    LocalMux I__4996 (
            .O(N__24131),
            .I(N__24123));
    LocalMux I__4995 (
            .O(N__24128),
            .I(N__24123));
    Odrv12 I__4994 (
            .O(N__24123),
            .I(\c0.n5497 ));
    CascadeMux I__4993 (
            .O(N__24120),
            .I(N__24116));
    InMux I__4992 (
            .O(N__24119),
            .I(N__24113));
    InMux I__4991 (
            .O(N__24116),
            .I(N__24110));
    LocalMux I__4990 (
            .O(N__24113),
            .I(N__24107));
    LocalMux I__4989 (
            .O(N__24110),
            .I(N__24104));
    Odrv12 I__4988 (
            .O(N__24107),
            .I(\c0.n5515 ));
    Odrv4 I__4987 (
            .O(N__24104),
            .I(\c0.n5515 ));
    InMux I__4986 (
            .O(N__24099),
            .I(N__24093));
    InMux I__4985 (
            .O(N__24098),
            .I(N__24086));
    InMux I__4984 (
            .O(N__24097),
            .I(N__24086));
    InMux I__4983 (
            .O(N__24096),
            .I(N__24086));
    LocalMux I__4982 (
            .O(N__24093),
            .I(r_Clock_Count_6));
    LocalMux I__4981 (
            .O(N__24086),
            .I(r_Clock_Count_6));
    CascadeMux I__4980 (
            .O(N__24081),
            .I(N__24078));
    InMux I__4979 (
            .O(N__24078),
            .I(N__24075));
    LocalMux I__4978 (
            .O(N__24075),
            .I(N__24072));
    Odrv4 I__4977 (
            .O(N__24072),
            .I(n317));
    CascadeMux I__4976 (
            .O(N__24069),
            .I(N__24063));
    InMux I__4975 (
            .O(N__24068),
            .I(N__24060));
    InMux I__4974 (
            .O(N__24067),
            .I(N__24055));
    InMux I__4973 (
            .O(N__24066),
            .I(N__24055));
    InMux I__4972 (
            .O(N__24063),
            .I(N__24052));
    LocalMux I__4971 (
            .O(N__24060),
            .I(r_Clock_Count_4));
    LocalMux I__4970 (
            .O(N__24055),
            .I(r_Clock_Count_4));
    LocalMux I__4969 (
            .O(N__24052),
            .I(r_Clock_Count_4));
    InMux I__4968 (
            .O(N__24045),
            .I(N__24042));
    LocalMux I__4967 (
            .O(N__24042),
            .I(\c0.tx.n10_adj_1868 ));
    CascadeMux I__4966 (
            .O(N__24039),
            .I(N__24034));
    InMux I__4965 (
            .O(N__24038),
            .I(N__24030));
    InMux I__4964 (
            .O(N__24037),
            .I(N__24027));
    InMux I__4963 (
            .O(N__24034),
            .I(N__24024));
    InMux I__4962 (
            .O(N__24033),
            .I(N__24021));
    LocalMux I__4961 (
            .O(N__24030),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__4960 (
            .O(N__24027),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__4959 (
            .O(N__24024),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__4958 (
            .O(N__24021),
            .I(\c0.tx.r_Clock_Count_7 ));
    InMux I__4957 (
            .O(N__24012),
            .I(N__24009));
    LocalMux I__4956 (
            .O(N__24009),
            .I(\c0.tx.n5627 ));
    CascadeMux I__4955 (
            .O(N__24006),
            .I(n11_adj_1979_cascade_));
    InMux I__4954 (
            .O(N__24003),
            .I(N__24000));
    LocalMux I__4953 (
            .O(N__24000),
            .I(\c0.tx.n5629 ));
    InMux I__4952 (
            .O(N__23997),
            .I(N__23993));
    InMux I__4951 (
            .O(N__23996),
            .I(N__23990));
    LocalMux I__4950 (
            .O(N__23993),
            .I(\c0.tx.n3120 ));
    LocalMux I__4949 (
            .O(N__23990),
            .I(\c0.tx.n3120 ));
    CascadeMux I__4948 (
            .O(N__23985),
            .I(N__23981));
    CascadeMux I__4947 (
            .O(N__23984),
            .I(N__23974));
    InMux I__4946 (
            .O(N__23981),
            .I(N__23971));
    InMux I__4945 (
            .O(N__23980),
            .I(N__23968));
    InMux I__4944 (
            .O(N__23979),
            .I(N__23963));
    InMux I__4943 (
            .O(N__23978),
            .I(N__23963));
    InMux I__4942 (
            .O(N__23977),
            .I(N__23960));
    InMux I__4941 (
            .O(N__23974),
            .I(N__23957));
    LocalMux I__4940 (
            .O(N__23971),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__4939 (
            .O(N__23968),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__4938 (
            .O(N__23963),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__4937 (
            .O(N__23960),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__4936 (
            .O(N__23957),
            .I(\c0.tx.r_Clock_Count_2 ));
    CascadeMux I__4935 (
            .O(N__23946),
            .I(\c0.tx.n3120_cascade_ ));
    InMux I__4934 (
            .O(N__23943),
            .I(N__23940));
    LocalMux I__4933 (
            .O(N__23940),
            .I(N__23937));
    Odrv4 I__4932 (
            .O(N__23937),
            .I(n313));
    CascadeMux I__4931 (
            .O(N__23934),
            .I(n782_cascade_));
    InMux I__4930 (
            .O(N__23931),
            .I(N__23925));
    InMux I__4929 (
            .O(N__23930),
            .I(N__23922));
    InMux I__4928 (
            .O(N__23929),
            .I(N__23917));
    InMux I__4927 (
            .O(N__23928),
            .I(N__23917));
    LocalMux I__4926 (
            .O(N__23925),
            .I(r_Clock_Count_8));
    LocalMux I__4925 (
            .O(N__23922),
            .I(r_Clock_Count_8));
    LocalMux I__4924 (
            .O(N__23917),
            .I(r_Clock_Count_8));
    CascadeMux I__4923 (
            .O(N__23910),
            .I(N__23907));
    InMux I__4922 (
            .O(N__23907),
            .I(N__23904));
    LocalMux I__4921 (
            .O(N__23904),
            .I(N__23901));
    Span4Mux_v I__4920 (
            .O(N__23901),
            .I(N__23898));
    Span4Mux_v I__4919 (
            .O(N__23898),
            .I(N__23894));
    InMux I__4918 (
            .O(N__23897),
            .I(N__23891));
    Sp12to4 I__4917 (
            .O(N__23894),
            .I(N__23885));
    LocalMux I__4916 (
            .O(N__23891),
            .I(N__23885));
    InMux I__4915 (
            .O(N__23890),
            .I(N__23882));
    Odrv12 I__4914 (
            .O(N__23885),
            .I(data_in_9_2));
    LocalMux I__4913 (
            .O(N__23882),
            .I(data_in_9_2));
    InMux I__4912 (
            .O(N__23877),
            .I(N__23874));
    LocalMux I__4911 (
            .O(N__23874),
            .I(\c0.n5827 ));
    CascadeMux I__4910 (
            .O(N__23871),
            .I(N__23868));
    InMux I__4909 (
            .O(N__23868),
            .I(N__23865));
    LocalMux I__4908 (
            .O(N__23865),
            .I(\c0.n1253 ));
    InMux I__4907 (
            .O(N__23862),
            .I(N__23859));
    LocalMux I__4906 (
            .O(N__23859),
            .I(N__23856));
    Span4Mux_h I__4905 (
            .O(N__23856),
            .I(N__23853));
    Span4Mux_h I__4904 (
            .O(N__23853),
            .I(N__23850));
    Odrv4 I__4903 (
            .O(N__23850),
            .I(tx_data_7_N_keep));
    InMux I__4902 (
            .O(N__23847),
            .I(N__23843));
    InMux I__4901 (
            .O(N__23846),
            .I(N__23840));
    LocalMux I__4900 (
            .O(N__23843),
            .I(data_out_18_0));
    LocalMux I__4899 (
            .O(N__23840),
            .I(data_out_18_0));
    CascadeMux I__4898 (
            .O(N__23835),
            .I(N__23832));
    InMux I__4897 (
            .O(N__23832),
            .I(N__23828));
    InMux I__4896 (
            .O(N__23831),
            .I(N__23825));
    LocalMux I__4895 (
            .O(N__23828),
            .I(N__23822));
    LocalMux I__4894 (
            .O(N__23825),
            .I(data_out_19_0));
    Odrv4 I__4893 (
            .O(N__23822),
            .I(data_out_19_0));
    InMux I__4892 (
            .O(N__23817),
            .I(N__23814));
    LocalMux I__4891 (
            .O(N__23814),
            .I(\c0.n1198 ));
    CascadeMux I__4890 (
            .O(N__23811),
            .I(\c0.n5810_cascade_ ));
    InMux I__4889 (
            .O(N__23808),
            .I(N__23804));
    InMux I__4888 (
            .O(N__23807),
            .I(N__23801));
    LocalMux I__4887 (
            .O(N__23804),
            .I(\c0.tx_data_0_N ));
    LocalMux I__4886 (
            .O(N__23801),
            .I(\c0.tx_data_0_N ));
    CascadeMux I__4885 (
            .O(N__23796),
            .I(\c0.tx.n14_adj_1869_cascade_ ));
    CascadeMux I__4884 (
            .O(N__23793),
            .I(\c0.tx.r_SM_Main_2_N_1767_1_cascade_ ));
    InMux I__4883 (
            .O(N__23790),
            .I(N__23787));
    LocalMux I__4882 (
            .O(N__23787),
            .I(N__23784));
    Odrv4 I__4881 (
            .O(N__23784),
            .I(\c0.tx.n5821 ));
    InMux I__4880 (
            .O(N__23781),
            .I(N__23775));
    InMux I__4879 (
            .O(N__23780),
            .I(N__23768));
    InMux I__4878 (
            .O(N__23779),
            .I(N__23768));
    InMux I__4877 (
            .O(N__23778),
            .I(N__23768));
    LocalMux I__4876 (
            .O(N__23775),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__4875 (
            .O(N__23768),
            .I(\c0.tx.r_Clock_Count_5 ));
    CascadeMux I__4874 (
            .O(N__23763),
            .I(N__23760));
    InMux I__4873 (
            .O(N__23760),
            .I(N__23757));
    LocalMux I__4872 (
            .O(N__23757),
            .I(N__23754));
    Odrv4 I__4871 (
            .O(N__23754),
            .I(n315));
    CascadeMux I__4870 (
            .O(N__23751),
            .I(\c0.n17_adj_1913_cascade_ ));
    InMux I__4869 (
            .O(N__23748),
            .I(N__23745));
    LocalMux I__4868 (
            .O(N__23745),
            .I(\c0.tx.n5883 ));
    CascadeMux I__4867 (
            .O(N__23742),
            .I(\c0.n1253_cascade_ ));
    InMux I__4866 (
            .O(N__23739),
            .I(N__23736));
    LocalMux I__4865 (
            .O(N__23736),
            .I(N__23733));
    Odrv4 I__4864 (
            .O(N__23733),
            .I(\c0.n5830 ));
    CascadeMux I__4863 (
            .O(N__23730),
            .I(\c0.n22_adj_1914_cascade_ ));
    InMux I__4862 (
            .O(N__23727),
            .I(N__23724));
    LocalMux I__4861 (
            .O(N__23724),
            .I(tx_data_6_N_keep));
    CascadeMux I__4860 (
            .O(N__23721),
            .I(n5646_cascade_));
    InMux I__4859 (
            .O(N__23718),
            .I(N__23715));
    LocalMux I__4858 (
            .O(N__23715),
            .I(n5645));
    IoInMux I__4857 (
            .O(N__23712),
            .I(N__23709));
    LocalMux I__4856 (
            .O(N__23709),
            .I(N__23706));
    Span4Mux_s0_v I__4855 (
            .O(N__23706),
            .I(N__23703));
    Span4Mux_h I__4854 (
            .O(N__23703),
            .I(N__23700));
    Span4Mux_v I__4853 (
            .O(N__23700),
            .I(N__23697));
    Span4Mux_v I__4852 (
            .O(N__23697),
            .I(N__23694));
    Odrv4 I__4851 (
            .O(N__23694),
            .I(LED_c));
    InMux I__4850 (
            .O(N__23691),
            .I(N__23688));
    LocalMux I__4849 (
            .O(N__23688),
            .I(N__23685));
    Span4Mux_v I__4848 (
            .O(N__23685),
            .I(N__23681));
    InMux I__4847 (
            .O(N__23684),
            .I(N__23678));
    Span4Mux_h I__4846 (
            .O(N__23681),
            .I(N__23672));
    LocalMux I__4845 (
            .O(N__23678),
            .I(N__23669));
    InMux I__4844 (
            .O(N__23677),
            .I(N__23662));
    InMux I__4843 (
            .O(N__23676),
            .I(N__23662));
    InMux I__4842 (
            .O(N__23675),
            .I(N__23662));
    Odrv4 I__4841 (
            .O(N__23672),
            .I(\c0.data_in_field_110 ));
    Odrv12 I__4840 (
            .O(N__23669),
            .I(\c0.data_in_field_110 ));
    LocalMux I__4839 (
            .O(N__23662),
            .I(\c0.data_in_field_110 ));
    InMux I__4838 (
            .O(N__23655),
            .I(N__23651));
    InMux I__4837 (
            .O(N__23654),
            .I(N__23648));
    LocalMux I__4836 (
            .O(N__23651),
            .I(N__23643));
    LocalMux I__4835 (
            .O(N__23648),
            .I(N__23643));
    Span4Mux_v I__4834 (
            .O(N__23643),
            .I(N__23640));
    Odrv4 I__4833 (
            .O(N__23640),
            .I(\c0.n5533 ));
    CascadeMux I__4832 (
            .O(N__23637),
            .I(N__23634));
    InMux I__4831 (
            .O(N__23634),
            .I(N__23630));
    InMux I__4830 (
            .O(N__23633),
            .I(N__23627));
    LocalMux I__4829 (
            .O(N__23630),
            .I(data_out_18_6));
    LocalMux I__4828 (
            .O(N__23627),
            .I(data_out_18_6));
    InMux I__4827 (
            .O(N__23622),
            .I(N__23619));
    LocalMux I__4826 (
            .O(N__23619),
            .I(N__23616));
    Span4Mux_h I__4825 (
            .O(N__23616),
            .I(N__23613));
    Odrv4 I__4824 (
            .O(N__23613),
            .I(\c0.n2077 ));
    InMux I__4823 (
            .O(N__23610),
            .I(N__23607));
    LocalMux I__4822 (
            .O(N__23607),
            .I(N__23604));
    Span4Mux_v I__4821 (
            .O(N__23604),
            .I(N__23601));
    Odrv4 I__4820 (
            .O(N__23601),
            .I(\c0.n5707 ));
    InMux I__4819 (
            .O(N__23598),
            .I(N__23595));
    LocalMux I__4818 (
            .O(N__23595),
            .I(N__23592));
    Odrv12 I__4817 (
            .O(N__23592),
            .I(\c0.n5710 ));
    InMux I__4816 (
            .O(N__23589),
            .I(N__23586));
    LocalMux I__4815 (
            .O(N__23586),
            .I(N__23583));
    Span4Mux_h I__4814 (
            .O(N__23583),
            .I(N__23580));
    Span4Mux_h I__4813 (
            .O(N__23580),
            .I(N__23577));
    Odrv4 I__4812 (
            .O(N__23577),
            .I(\c0.n6198 ));
    InMux I__4811 (
            .O(N__23574),
            .I(N__23570));
    InMux I__4810 (
            .O(N__23573),
            .I(N__23567));
    LocalMux I__4809 (
            .O(N__23570),
            .I(\c0.delay_counter_9 ));
    LocalMux I__4808 (
            .O(N__23567),
            .I(\c0.delay_counter_9 ));
    InMux I__4807 (
            .O(N__23562),
            .I(N__23558));
    InMux I__4806 (
            .O(N__23561),
            .I(N__23555));
    LocalMux I__4805 (
            .O(N__23558),
            .I(\c0.delay_counter_2 ));
    LocalMux I__4804 (
            .O(N__23555),
            .I(\c0.delay_counter_2 ));
    CascadeMux I__4803 (
            .O(N__23550),
            .I(N__23546));
    InMux I__4802 (
            .O(N__23549),
            .I(N__23543));
    InMux I__4801 (
            .O(N__23546),
            .I(N__23540));
    LocalMux I__4800 (
            .O(N__23543),
            .I(\c0.delay_counter_0 ));
    LocalMux I__4799 (
            .O(N__23540),
            .I(\c0.delay_counter_0 ));
    InMux I__4798 (
            .O(N__23535),
            .I(N__23531));
    InMux I__4797 (
            .O(N__23534),
            .I(N__23528));
    LocalMux I__4796 (
            .O(N__23531),
            .I(\c0.delay_counter_7 ));
    LocalMux I__4795 (
            .O(N__23528),
            .I(\c0.delay_counter_7 ));
    CascadeMux I__4794 (
            .O(N__23523),
            .I(N__23520));
    InMux I__4793 (
            .O(N__23520),
            .I(N__23517));
    LocalMux I__4792 (
            .O(N__23517),
            .I(N__23514));
    Span4Mux_h I__4791 (
            .O(N__23514),
            .I(N__23511));
    Span4Mux_v I__4790 (
            .O(N__23511),
            .I(N__23506));
    InMux I__4789 (
            .O(N__23510),
            .I(N__23501));
    InMux I__4788 (
            .O(N__23509),
            .I(N__23501));
    Odrv4 I__4787 (
            .O(N__23506),
            .I(data_in_5_0));
    LocalMux I__4786 (
            .O(N__23501),
            .I(data_in_5_0));
    InMux I__4785 (
            .O(N__23496),
            .I(N__23493));
    LocalMux I__4784 (
            .O(N__23493),
            .I(N__23489));
    InMux I__4783 (
            .O(N__23492),
            .I(N__23486));
    Span4Mux_v I__4782 (
            .O(N__23489),
            .I(N__23483));
    LocalMux I__4781 (
            .O(N__23486),
            .I(N__23480));
    Span4Mux_v I__4780 (
            .O(N__23483),
            .I(N__23477));
    Span4Mux_h I__4779 (
            .O(N__23480),
            .I(N__23474));
    Sp12to4 I__4778 (
            .O(N__23477),
            .I(N__23470));
    Span4Mux_v I__4777 (
            .O(N__23474),
            .I(N__23467));
    InMux I__4776 (
            .O(N__23473),
            .I(N__23464));
    Odrv12 I__4775 (
            .O(N__23470),
            .I(data_in_4_0));
    Odrv4 I__4774 (
            .O(N__23467),
            .I(data_in_4_0));
    LocalMux I__4773 (
            .O(N__23464),
            .I(data_in_4_0));
    InMux I__4772 (
            .O(N__23457),
            .I(N__23453));
    InMux I__4771 (
            .O(N__23456),
            .I(N__23450));
    LocalMux I__4770 (
            .O(N__23453),
            .I(N__23446));
    LocalMux I__4769 (
            .O(N__23450),
            .I(N__23443));
    InMux I__4768 (
            .O(N__23449),
            .I(N__23440));
    Span4Mux_h I__4767 (
            .O(N__23446),
            .I(N__23437));
    Span4Mux_v I__4766 (
            .O(N__23443),
            .I(N__23434));
    LocalMux I__4765 (
            .O(N__23440),
            .I(data_in_8_4));
    Odrv4 I__4764 (
            .O(N__23437),
            .I(data_in_8_4));
    Odrv4 I__4763 (
            .O(N__23434),
            .I(data_in_8_4));
    CascadeMux I__4762 (
            .O(N__23427),
            .I(N__23424));
    InMux I__4761 (
            .O(N__23424),
            .I(N__23421));
    LocalMux I__4760 (
            .O(N__23421),
            .I(N__23418));
    Span4Mux_h I__4759 (
            .O(N__23418),
            .I(N__23415));
    Span4Mux_v I__4758 (
            .O(N__23415),
            .I(N__23410));
    InMux I__4757 (
            .O(N__23414),
            .I(N__23405));
    InMux I__4756 (
            .O(N__23413),
            .I(N__23405));
    Odrv4 I__4755 (
            .O(N__23410),
            .I(data_in_7_4));
    LocalMux I__4754 (
            .O(N__23405),
            .I(data_in_7_4));
    CascadeMux I__4753 (
            .O(N__23400),
            .I(N__23397));
    InMux I__4752 (
            .O(N__23397),
            .I(N__23393));
    InMux I__4751 (
            .O(N__23396),
            .I(N__23390));
    LocalMux I__4750 (
            .O(N__23393),
            .I(N__23387));
    LocalMux I__4749 (
            .O(N__23390),
            .I(N__23384));
    Span4Mux_v I__4748 (
            .O(N__23387),
            .I(N__23380));
    Span12Mux_v I__4747 (
            .O(N__23384),
            .I(N__23377));
    InMux I__4746 (
            .O(N__23383),
            .I(N__23374));
    Odrv4 I__4745 (
            .O(N__23380),
            .I(data_in_6_4));
    Odrv12 I__4744 (
            .O(N__23377),
            .I(data_in_6_4));
    LocalMux I__4743 (
            .O(N__23374),
            .I(data_in_6_4));
    CascadeMux I__4742 (
            .O(N__23367),
            .I(N__23364));
    InMux I__4741 (
            .O(N__23364),
            .I(N__23361));
    LocalMux I__4740 (
            .O(N__23361),
            .I(N__23358));
    Span4Mux_v I__4739 (
            .O(N__23358),
            .I(N__23355));
    Span4Mux_v I__4738 (
            .O(N__23355),
            .I(N__23350));
    InMux I__4737 (
            .O(N__23354),
            .I(N__23345));
    InMux I__4736 (
            .O(N__23353),
            .I(N__23345));
    Odrv4 I__4735 (
            .O(N__23350),
            .I(data_in_5_6));
    LocalMux I__4734 (
            .O(N__23345),
            .I(data_in_5_6));
    InMux I__4733 (
            .O(N__23340),
            .I(N__23335));
    InMux I__4732 (
            .O(N__23339),
            .I(N__23332));
    InMux I__4731 (
            .O(N__23338),
            .I(N__23328));
    LocalMux I__4730 (
            .O(N__23335),
            .I(N__23325));
    LocalMux I__4729 (
            .O(N__23332),
            .I(N__23322));
    InMux I__4728 (
            .O(N__23331),
            .I(N__23319));
    LocalMux I__4727 (
            .O(N__23328),
            .I(\c0.data_in_field_89 ));
    Odrv12 I__4726 (
            .O(N__23325),
            .I(\c0.data_in_field_89 ));
    Odrv4 I__4725 (
            .O(N__23322),
            .I(\c0.data_in_field_89 ));
    LocalMux I__4724 (
            .O(N__23319),
            .I(\c0.data_in_field_89 ));
    InMux I__4723 (
            .O(N__23310),
            .I(N__23307));
    LocalMux I__4722 (
            .O(N__23307),
            .I(N__23303));
    InMux I__4721 (
            .O(N__23306),
            .I(N__23300));
    Span12Mux_s9_h I__4720 (
            .O(N__23303),
            .I(N__23294));
    LocalMux I__4719 (
            .O(N__23300),
            .I(N__23291));
    InMux I__4718 (
            .O(N__23299),
            .I(N__23284));
    InMux I__4717 (
            .O(N__23298),
            .I(N__23284));
    InMux I__4716 (
            .O(N__23297),
            .I(N__23284));
    Odrv12 I__4715 (
            .O(N__23294),
            .I(\c0.data_in_field_90 ));
    Odrv4 I__4714 (
            .O(N__23291),
            .I(\c0.data_in_field_90 ));
    LocalMux I__4713 (
            .O(N__23284),
            .I(\c0.data_in_field_90 ));
    CascadeMux I__4712 (
            .O(N__23277),
            .I(N__23274));
    InMux I__4711 (
            .O(N__23274),
            .I(N__23271));
    LocalMux I__4710 (
            .O(N__23271),
            .I(N__23268));
    Span4Mux_v I__4709 (
            .O(N__23268),
            .I(N__23264));
    InMux I__4708 (
            .O(N__23267),
            .I(N__23261));
    Span4Mux_h I__4707 (
            .O(N__23264),
            .I(N__23256));
    LocalMux I__4706 (
            .O(N__23261),
            .I(N__23256));
    Span4Mux_h I__4705 (
            .O(N__23256),
            .I(N__23253));
    Span4Mux_h I__4704 (
            .O(N__23253),
            .I(N__23250));
    Span4Mux_v I__4703 (
            .O(N__23250),
            .I(N__23246));
    InMux I__4702 (
            .O(N__23249),
            .I(N__23243));
    Odrv4 I__4701 (
            .O(N__23246),
            .I(data_in_7_7));
    LocalMux I__4700 (
            .O(N__23243),
            .I(data_in_7_7));
    InMux I__4699 (
            .O(N__23238),
            .I(N__23234));
    InMux I__4698 (
            .O(N__23237),
            .I(N__23231));
    LocalMux I__4697 (
            .O(N__23234),
            .I(N__23228));
    LocalMux I__4696 (
            .O(N__23231),
            .I(N__23222));
    Span4Mux_v I__4695 (
            .O(N__23228),
            .I(N__23222));
    InMux I__4694 (
            .O(N__23227),
            .I(N__23218));
    Span4Mux_h I__4693 (
            .O(N__23222),
            .I(N__23215));
    InMux I__4692 (
            .O(N__23221),
            .I(N__23212));
    LocalMux I__4691 (
            .O(N__23218),
            .I(\c0.data_in_field_37 ));
    Odrv4 I__4690 (
            .O(N__23215),
            .I(\c0.data_in_field_37 ));
    LocalMux I__4689 (
            .O(N__23212),
            .I(\c0.data_in_field_37 ));
    InMux I__4688 (
            .O(N__23205),
            .I(N__23202));
    LocalMux I__4687 (
            .O(N__23202),
            .I(N__23199));
    Span4Mux_v I__4686 (
            .O(N__23199),
            .I(N__23196));
    Span4Mux_h I__4685 (
            .O(N__23196),
            .I(N__23192));
    InMux I__4684 (
            .O(N__23195),
            .I(N__23189));
    Span4Mux_h I__4683 (
            .O(N__23192),
            .I(N__23186));
    LocalMux I__4682 (
            .O(N__23189),
            .I(\c0.data_in_frame_18_0 ));
    Odrv4 I__4681 (
            .O(N__23186),
            .I(\c0.data_in_frame_18_0 ));
    InMux I__4680 (
            .O(N__23181),
            .I(N__23177));
    InMux I__4679 (
            .O(N__23180),
            .I(N__23174));
    LocalMux I__4678 (
            .O(N__23177),
            .I(N__23170));
    LocalMux I__4677 (
            .O(N__23174),
            .I(N__23167));
    InMux I__4676 (
            .O(N__23173),
            .I(N__23164));
    Odrv12 I__4675 (
            .O(N__23170),
            .I(data_in_4_1));
    Odrv4 I__4674 (
            .O(N__23167),
            .I(data_in_4_1));
    LocalMux I__4673 (
            .O(N__23164),
            .I(data_in_4_1));
    CascadeMux I__4672 (
            .O(N__23157),
            .I(N__23153));
    CascadeMux I__4671 (
            .O(N__23156),
            .I(N__23150));
    InMux I__4670 (
            .O(N__23153),
            .I(N__23146));
    InMux I__4669 (
            .O(N__23150),
            .I(N__23143));
    InMux I__4668 (
            .O(N__23149),
            .I(N__23140));
    LocalMux I__4667 (
            .O(N__23146),
            .I(N__23137));
    LocalMux I__4666 (
            .O(N__23143),
            .I(N__23133));
    LocalMux I__4665 (
            .O(N__23140),
            .I(N__23130));
    Span4Mux_h I__4664 (
            .O(N__23137),
            .I(N__23127));
    InMux I__4663 (
            .O(N__23136),
            .I(N__23124));
    Span4Mux_v I__4662 (
            .O(N__23133),
            .I(N__23121));
    Span4Mux_h I__4661 (
            .O(N__23130),
            .I(N__23116));
    Span4Mux_v I__4660 (
            .O(N__23127),
            .I(N__23116));
    LocalMux I__4659 (
            .O(N__23124),
            .I(data_in_18_7));
    Odrv4 I__4658 (
            .O(N__23121),
            .I(data_in_18_7));
    Odrv4 I__4657 (
            .O(N__23116),
            .I(data_in_18_7));
    InMux I__4656 (
            .O(N__23109),
            .I(N__23106));
    LocalMux I__4655 (
            .O(N__23106),
            .I(N__23103));
    Span4Mux_v I__4654 (
            .O(N__23103),
            .I(N__23099));
    InMux I__4653 (
            .O(N__23102),
            .I(N__23096));
    Span4Mux_v I__4652 (
            .O(N__23099),
            .I(N__23092));
    LocalMux I__4651 (
            .O(N__23096),
            .I(N__23089));
    InMux I__4650 (
            .O(N__23095),
            .I(N__23086));
    Odrv4 I__4649 (
            .O(N__23092),
            .I(data_in_17_7));
    Odrv4 I__4648 (
            .O(N__23089),
            .I(data_in_17_7));
    LocalMux I__4647 (
            .O(N__23086),
            .I(data_in_17_7));
    InMux I__4646 (
            .O(N__23079),
            .I(N__23076));
    LocalMux I__4645 (
            .O(N__23076),
            .I(N__23073));
    Odrv12 I__4644 (
            .O(N__23073),
            .I(\c0.n6_adj_1918 ));
    InMux I__4643 (
            .O(N__23070),
            .I(N__23066));
    CascadeMux I__4642 (
            .O(N__23069),
            .I(N__23063));
    LocalMux I__4641 (
            .O(N__23066),
            .I(N__23059));
    InMux I__4640 (
            .O(N__23063),
            .I(N__23056));
    InMux I__4639 (
            .O(N__23062),
            .I(N__23053));
    Span4Mux_v I__4638 (
            .O(N__23059),
            .I(N__23048));
    LocalMux I__4637 (
            .O(N__23056),
            .I(N__23048));
    LocalMux I__4636 (
            .O(N__23053),
            .I(N__23044));
    Span4Mux_h I__4635 (
            .O(N__23048),
            .I(N__23041));
    InMux I__4634 (
            .O(N__23047),
            .I(N__23038));
    Span12Mux_s9_h I__4633 (
            .O(N__23044),
            .I(N__23035));
    Span4Mux_v I__4632 (
            .O(N__23041),
            .I(N__23032));
    LocalMux I__4631 (
            .O(N__23038),
            .I(data_in_1_4));
    Odrv12 I__4630 (
            .O(N__23035),
            .I(data_in_1_4));
    Odrv4 I__4629 (
            .O(N__23032),
            .I(data_in_1_4));
    InMux I__4628 (
            .O(N__23025),
            .I(N__23022));
    LocalMux I__4627 (
            .O(N__23022),
            .I(N__23017));
    InMux I__4626 (
            .O(N__23021),
            .I(N__23014));
    CascadeMux I__4625 (
            .O(N__23020),
            .I(N__23010));
    Span4Mux_h I__4624 (
            .O(N__23017),
            .I(N__23007));
    LocalMux I__4623 (
            .O(N__23014),
            .I(N__23004));
    CascadeMux I__4622 (
            .O(N__23013),
            .I(N__23000));
    InMux I__4621 (
            .O(N__23010),
            .I(N__22997));
    Span4Mux_v I__4620 (
            .O(N__23007),
            .I(N__22994));
    Span4Mux_v I__4619 (
            .O(N__23004),
            .I(N__22991));
    InMux I__4618 (
            .O(N__23003),
            .I(N__22986));
    InMux I__4617 (
            .O(N__23000),
            .I(N__22986));
    LocalMux I__4616 (
            .O(N__22997),
            .I(\c0.data_in_field_18 ));
    Odrv4 I__4615 (
            .O(N__22994),
            .I(\c0.data_in_field_18 ));
    Odrv4 I__4614 (
            .O(N__22991),
            .I(\c0.data_in_field_18 ));
    LocalMux I__4613 (
            .O(N__22986),
            .I(\c0.data_in_field_18 ));
    InMux I__4612 (
            .O(N__22977),
            .I(N__22974));
    LocalMux I__4611 (
            .O(N__22974),
            .I(\c0.n5372 ));
    CascadeMux I__4610 (
            .O(N__22971),
            .I(\c0.n2043_cascade_ ));
    InMux I__4609 (
            .O(N__22968),
            .I(N__22963));
    InMux I__4608 (
            .O(N__22967),
            .I(N__22960));
    InMux I__4607 (
            .O(N__22966),
            .I(N__22956));
    LocalMux I__4606 (
            .O(N__22963),
            .I(N__22953));
    LocalMux I__4605 (
            .O(N__22960),
            .I(N__22950));
    InMux I__4604 (
            .O(N__22959),
            .I(N__22946));
    LocalMux I__4603 (
            .O(N__22956),
            .I(N__22943));
    Span4Mux_h I__4602 (
            .O(N__22953),
            .I(N__22940));
    Span4Mux_h I__4601 (
            .O(N__22950),
            .I(N__22937));
    InMux I__4600 (
            .O(N__22949),
            .I(N__22934));
    LocalMux I__4599 (
            .O(N__22946),
            .I(\c0.data_in_field_107 ));
    Odrv12 I__4598 (
            .O(N__22943),
            .I(\c0.data_in_field_107 ));
    Odrv4 I__4597 (
            .O(N__22940),
            .I(\c0.data_in_field_107 ));
    Odrv4 I__4596 (
            .O(N__22937),
            .I(\c0.data_in_field_107 ));
    LocalMux I__4595 (
            .O(N__22934),
            .I(\c0.data_in_field_107 ));
    InMux I__4594 (
            .O(N__22923),
            .I(N__22920));
    LocalMux I__4593 (
            .O(N__22920),
            .I(N__22917));
    Span4Mux_h I__4592 (
            .O(N__22917),
            .I(N__22912));
    InMux I__4591 (
            .O(N__22916),
            .I(N__22909));
    InMux I__4590 (
            .O(N__22915),
            .I(N__22906));
    Span4Mux_v I__4589 (
            .O(N__22912),
            .I(N__22903));
    LocalMux I__4588 (
            .O(N__22909),
            .I(data_in_13_6));
    LocalMux I__4587 (
            .O(N__22906),
            .I(data_in_13_6));
    Odrv4 I__4586 (
            .O(N__22903),
            .I(data_in_13_6));
    InMux I__4585 (
            .O(N__22896),
            .I(N__22892));
    CascadeMux I__4584 (
            .O(N__22895),
            .I(N__22889));
    LocalMux I__4583 (
            .O(N__22892),
            .I(N__22886));
    InMux I__4582 (
            .O(N__22889),
            .I(N__22883));
    Sp12to4 I__4581 (
            .O(N__22886),
            .I(N__22878));
    LocalMux I__4580 (
            .O(N__22883),
            .I(N__22878));
    Span12Mux_s11_v I__4579 (
            .O(N__22878),
            .I(N__22875));
    Odrv12 I__4578 (
            .O(N__22875),
            .I(\c0.n5443 ));
    InMux I__4577 (
            .O(N__22872),
            .I(N__22869));
    LocalMux I__4576 (
            .O(N__22869),
            .I(N__22866));
    Span4Mux_v I__4575 (
            .O(N__22866),
            .I(N__22863));
    Odrv4 I__4574 (
            .O(N__22863),
            .I(\c0.n47_adj_1897 ));
    InMux I__4573 (
            .O(N__22860),
            .I(N__22857));
    LocalMux I__4572 (
            .O(N__22857),
            .I(N__22854));
    Span4Mux_h I__4571 (
            .O(N__22854),
            .I(N__22851));
    Odrv4 I__4570 (
            .O(N__22851),
            .I(\c0.n48_adj_1895 ));
    CascadeMux I__4569 (
            .O(N__22848),
            .I(\c0.n5567_cascade_ ));
    InMux I__4568 (
            .O(N__22845),
            .I(N__22842));
    LocalMux I__4567 (
            .O(N__22842),
            .I(\c0.n49 ));
    CascadeMux I__4566 (
            .O(N__22839),
            .I(N__22836));
    InMux I__4565 (
            .O(N__22836),
            .I(N__22833));
    LocalMux I__4564 (
            .O(N__22833),
            .I(N__22830));
    Span4Mux_v I__4563 (
            .O(N__22830),
            .I(N__22827));
    Odrv4 I__4562 (
            .O(N__22827),
            .I(\c0.n6219 ));
    InMux I__4561 (
            .O(N__22824),
            .I(N__22820));
    CascadeMux I__4560 (
            .O(N__22823),
            .I(N__22817));
    LocalMux I__4559 (
            .O(N__22820),
            .I(N__22814));
    InMux I__4558 (
            .O(N__22817),
            .I(N__22809));
    Span4Mux_v I__4557 (
            .O(N__22814),
            .I(N__22806));
    InMux I__4556 (
            .O(N__22813),
            .I(N__22801));
    InMux I__4555 (
            .O(N__22812),
            .I(N__22801));
    LocalMux I__4554 (
            .O(N__22809),
            .I(\c0.data_in_field_5 ));
    Odrv4 I__4553 (
            .O(N__22806),
            .I(\c0.data_in_field_5 ));
    LocalMux I__4552 (
            .O(N__22801),
            .I(\c0.data_in_field_5 ));
    InMux I__4551 (
            .O(N__22794),
            .I(N__22790));
    InMux I__4550 (
            .O(N__22793),
            .I(N__22787));
    LocalMux I__4549 (
            .O(N__22790),
            .I(N__22784));
    LocalMux I__4548 (
            .O(N__22787),
            .I(N__22781));
    Span4Mux_h I__4547 (
            .O(N__22784),
            .I(N__22778));
    Span4Mux_v I__4546 (
            .O(N__22781),
            .I(N__22773));
    Span4Mux_h I__4545 (
            .O(N__22778),
            .I(N__22773));
    Odrv4 I__4544 (
            .O(N__22773),
            .I(\c0.n1979 ));
    InMux I__4543 (
            .O(N__22770),
            .I(N__22767));
    LocalMux I__4542 (
            .O(N__22767),
            .I(N__22764));
    Span4Mux_h I__4541 (
            .O(N__22764),
            .I(N__22760));
    InMux I__4540 (
            .O(N__22763),
            .I(N__22757));
    Span4Mux_v I__4539 (
            .O(N__22760),
            .I(N__22752));
    LocalMux I__4538 (
            .O(N__22757),
            .I(N__22752));
    Odrv4 I__4537 (
            .O(N__22752),
            .I(\c0.n1958 ));
    InMux I__4536 (
            .O(N__22749),
            .I(N__22746));
    LocalMux I__4535 (
            .O(N__22746),
            .I(N__22743));
    Span4Mux_v I__4534 (
            .O(N__22743),
            .I(N__22739));
    InMux I__4533 (
            .O(N__22742),
            .I(N__22736));
    Span4Mux_h I__4532 (
            .O(N__22739),
            .I(N__22731));
    LocalMux I__4531 (
            .O(N__22736),
            .I(N__22731));
    Span4Mux_h I__4530 (
            .O(N__22731),
            .I(N__22728));
    Odrv4 I__4529 (
            .O(N__22728),
            .I(\c0.n2056 ));
    InMux I__4528 (
            .O(N__22725),
            .I(N__22722));
    LocalMux I__4527 (
            .O(N__22722),
            .I(\c0.n5506 ));
    InMux I__4526 (
            .O(N__22719),
            .I(N__22716));
    LocalMux I__4525 (
            .O(N__22716),
            .I(N__22713));
    Span4Mux_h I__4524 (
            .O(N__22713),
            .I(N__22709));
    InMux I__4523 (
            .O(N__22712),
            .I(N__22706));
    Span4Mux_h I__4522 (
            .O(N__22709),
            .I(N__22701));
    LocalMux I__4521 (
            .O(N__22706),
            .I(N__22701));
    Odrv4 I__4520 (
            .O(N__22701),
            .I(\c0.n5575 ));
    CascadeMux I__4519 (
            .O(N__22698),
            .I(\c0.n5506_cascade_ ));
    InMux I__4518 (
            .O(N__22695),
            .I(N__22692));
    LocalMux I__4517 (
            .O(N__22692),
            .I(N__22688));
    InMux I__4516 (
            .O(N__22691),
            .I(N__22685));
    Span4Mux_h I__4515 (
            .O(N__22688),
            .I(N__22682));
    LocalMux I__4514 (
            .O(N__22685),
            .I(N__22679));
    Odrv4 I__4513 (
            .O(N__22682),
            .I(\c0.n5539 ));
    Odrv4 I__4512 (
            .O(N__22679),
            .I(\c0.n5539 ));
    InMux I__4511 (
            .O(N__22674),
            .I(N__22670));
    InMux I__4510 (
            .O(N__22673),
            .I(N__22667));
    LocalMux I__4509 (
            .O(N__22670),
            .I(N__22664));
    LocalMux I__4508 (
            .O(N__22667),
            .I(N__22661));
    Span4Mux_v I__4507 (
            .O(N__22664),
            .I(N__22658));
    Span4Mux_h I__4506 (
            .O(N__22661),
            .I(N__22655));
    Odrv4 I__4505 (
            .O(N__22658),
            .I(\c0.n1779 ));
    Odrv4 I__4504 (
            .O(N__22655),
            .I(\c0.n1779 ));
    InMux I__4503 (
            .O(N__22650),
            .I(N__22646));
    InMux I__4502 (
            .O(N__22649),
            .I(N__22643));
    LocalMux I__4501 (
            .O(N__22646),
            .I(N__22639));
    LocalMux I__4500 (
            .O(N__22643),
            .I(N__22634));
    InMux I__4499 (
            .O(N__22642),
            .I(N__22631));
    Span4Mux_h I__4498 (
            .O(N__22639),
            .I(N__22628));
    InMux I__4497 (
            .O(N__22638),
            .I(N__22625));
    InMux I__4496 (
            .O(N__22637),
            .I(N__22622));
    Span4Mux_h I__4495 (
            .O(N__22634),
            .I(N__22619));
    LocalMux I__4494 (
            .O(N__22631),
            .I(\c0.data_in_field_60 ));
    Odrv4 I__4493 (
            .O(N__22628),
            .I(\c0.data_in_field_60 ));
    LocalMux I__4492 (
            .O(N__22625),
            .I(\c0.data_in_field_60 ));
    LocalMux I__4491 (
            .O(N__22622),
            .I(\c0.data_in_field_60 ));
    Odrv4 I__4490 (
            .O(N__22619),
            .I(\c0.data_in_field_60 ));
    InMux I__4489 (
            .O(N__22608),
            .I(N__22605));
    LocalMux I__4488 (
            .O(N__22605),
            .I(N__22601));
    InMux I__4487 (
            .O(N__22604),
            .I(N__22598));
    Odrv4 I__4486 (
            .O(N__22601),
            .I(\c0.n5500 ));
    LocalMux I__4485 (
            .O(N__22598),
            .I(\c0.n5500 ));
    InMux I__4484 (
            .O(N__22593),
            .I(N__22590));
    LocalMux I__4483 (
            .O(N__22590),
            .I(N__22586));
    InMux I__4482 (
            .O(N__22589),
            .I(N__22583));
    Span4Mux_h I__4481 (
            .O(N__22586),
            .I(N__22579));
    LocalMux I__4480 (
            .O(N__22583),
            .I(N__22576));
    InMux I__4479 (
            .O(N__22582),
            .I(N__22571));
    Span4Mux_h I__4478 (
            .O(N__22579),
            .I(N__22566));
    Span4Mux_h I__4477 (
            .O(N__22576),
            .I(N__22566));
    InMux I__4476 (
            .O(N__22575),
            .I(N__22563));
    InMux I__4475 (
            .O(N__22574),
            .I(N__22560));
    LocalMux I__4474 (
            .O(N__22571),
            .I(\c0.data_in_field_19 ));
    Odrv4 I__4473 (
            .O(N__22566),
            .I(\c0.data_in_field_19 ));
    LocalMux I__4472 (
            .O(N__22563),
            .I(\c0.data_in_field_19 ));
    LocalMux I__4471 (
            .O(N__22560),
            .I(\c0.data_in_field_19 ));
    InMux I__4470 (
            .O(N__22551),
            .I(N__22548));
    LocalMux I__4469 (
            .O(N__22548),
            .I(N__22545));
    Span4Mux_s3_h I__4468 (
            .O(N__22545),
            .I(N__22541));
    InMux I__4467 (
            .O(N__22544),
            .I(N__22538));
    Span4Mux_h I__4466 (
            .O(N__22541),
            .I(N__22535));
    LocalMux I__4465 (
            .O(N__22538),
            .I(N__22532));
    Span4Mux_v I__4464 (
            .O(N__22535),
            .I(N__22526));
    Span4Mux_h I__4463 (
            .O(N__22532),
            .I(N__22523));
    InMux I__4462 (
            .O(N__22531),
            .I(N__22520));
    InMux I__4461 (
            .O(N__22530),
            .I(N__22515));
    InMux I__4460 (
            .O(N__22529),
            .I(N__22515));
    Odrv4 I__4459 (
            .O(N__22526),
            .I(\c0.data_in_field_139 ));
    Odrv4 I__4458 (
            .O(N__22523),
            .I(\c0.data_in_field_139 ));
    LocalMux I__4457 (
            .O(N__22520),
            .I(\c0.data_in_field_139 ));
    LocalMux I__4456 (
            .O(N__22515),
            .I(\c0.data_in_field_139 ));
    CascadeMux I__4455 (
            .O(N__22506),
            .I(N__22503));
    InMux I__4454 (
            .O(N__22503),
            .I(N__22498));
    InMux I__4453 (
            .O(N__22502),
            .I(N__22495));
    InMux I__4452 (
            .O(N__22501),
            .I(N__22492));
    LocalMux I__4451 (
            .O(N__22498),
            .I(data_in_5_5));
    LocalMux I__4450 (
            .O(N__22495),
            .I(data_in_5_5));
    LocalMux I__4449 (
            .O(N__22492),
            .I(data_in_5_5));
    InMux I__4448 (
            .O(N__22485),
            .I(N__22481));
    CascadeMux I__4447 (
            .O(N__22484),
            .I(N__22478));
    LocalMux I__4446 (
            .O(N__22481),
            .I(N__22475));
    InMux I__4445 (
            .O(N__22478),
            .I(N__22472));
    Span4Mux_v I__4444 (
            .O(N__22475),
            .I(N__22469));
    LocalMux I__4443 (
            .O(N__22472),
            .I(N__22464));
    Span4Mux_h I__4442 (
            .O(N__22469),
            .I(N__22464));
    Span4Mux_h I__4441 (
            .O(N__22464),
            .I(N__22460));
    InMux I__4440 (
            .O(N__22463),
            .I(N__22457));
    Odrv4 I__4439 (
            .O(N__22460),
            .I(data_in_6_1));
    LocalMux I__4438 (
            .O(N__22457),
            .I(data_in_6_1));
    InMux I__4437 (
            .O(N__22452),
            .I(N__22449));
    LocalMux I__4436 (
            .O(N__22449),
            .I(N__22446));
    Span4Mux_v I__4435 (
            .O(N__22446),
            .I(N__22443));
    Span4Mux_h I__4434 (
            .O(N__22443),
            .I(N__22440));
    Span4Mux_h I__4433 (
            .O(N__22440),
            .I(N__22435));
    InMux I__4432 (
            .O(N__22439),
            .I(N__22430));
    InMux I__4431 (
            .O(N__22438),
            .I(N__22430));
    Odrv4 I__4430 (
            .O(N__22435),
            .I(data_in_5_1));
    LocalMux I__4429 (
            .O(N__22430),
            .I(data_in_5_1));
    InMux I__4428 (
            .O(N__22425),
            .I(N__22422));
    LocalMux I__4427 (
            .O(N__22422),
            .I(N__22419));
    Span4Mux_h I__4426 (
            .O(N__22419),
            .I(N__22416));
    Sp12to4 I__4425 (
            .O(N__22416),
            .I(N__22411));
    InMux I__4424 (
            .O(N__22415),
            .I(N__22406));
    InMux I__4423 (
            .O(N__22414),
            .I(N__22406));
    Odrv12 I__4422 (
            .O(N__22411),
            .I(data_in_16_7));
    LocalMux I__4421 (
            .O(N__22406),
            .I(data_in_16_7));
    InMux I__4420 (
            .O(N__22401),
            .I(N__22398));
    LocalMux I__4419 (
            .O(N__22398),
            .I(\c0.n25 ));
    CascadeMux I__4418 (
            .O(N__22395),
            .I(N__22392));
    InMux I__4417 (
            .O(N__22392),
            .I(N__22389));
    LocalMux I__4416 (
            .O(N__22389),
            .I(N__22386));
    Span4Mux_h I__4415 (
            .O(N__22386),
            .I(N__22383));
    Odrv4 I__4414 (
            .O(N__22383),
            .I(\c0.n23 ));
    InMux I__4413 (
            .O(N__22380),
            .I(N__22377));
    LocalMux I__4412 (
            .O(N__22377),
            .I(N__22374));
    Sp12to4 I__4411 (
            .O(N__22374),
            .I(N__22371));
    Span12Mux_v I__4410 (
            .O(N__22371),
            .I(N__22368));
    Odrv12 I__4409 (
            .O(N__22368),
            .I(\c0.n22_adj_1890 ));
    InMux I__4408 (
            .O(N__22365),
            .I(N__22360));
    InMux I__4407 (
            .O(N__22364),
            .I(N__22357));
    InMux I__4406 (
            .O(N__22363),
            .I(N__22354));
    LocalMux I__4405 (
            .O(N__22360),
            .I(N__22351));
    LocalMux I__4404 (
            .O(N__22357),
            .I(N__22347));
    LocalMux I__4403 (
            .O(N__22354),
            .I(N__22342));
    Span4Mux_h I__4402 (
            .O(N__22351),
            .I(N__22339));
    InMux I__4401 (
            .O(N__22350),
            .I(N__22336));
    Span4Mux_h I__4400 (
            .O(N__22347),
            .I(N__22333));
    InMux I__4399 (
            .O(N__22346),
            .I(N__22328));
    InMux I__4398 (
            .O(N__22345),
            .I(N__22328));
    Odrv12 I__4397 (
            .O(N__22342),
            .I(\c0.data_in_field_61 ));
    Odrv4 I__4396 (
            .O(N__22339),
            .I(\c0.data_in_field_61 ));
    LocalMux I__4395 (
            .O(N__22336),
            .I(\c0.data_in_field_61 ));
    Odrv4 I__4394 (
            .O(N__22333),
            .I(\c0.data_in_field_61 ));
    LocalMux I__4393 (
            .O(N__22328),
            .I(\c0.data_in_field_61 ));
    InMux I__4392 (
            .O(N__22317),
            .I(N__22313));
    InMux I__4391 (
            .O(N__22316),
            .I(N__22310));
    LocalMux I__4390 (
            .O(N__22313),
            .I(N__22304));
    LocalMux I__4389 (
            .O(N__22310),
            .I(N__22304));
    InMux I__4388 (
            .O(N__22309),
            .I(N__22301));
    Span4Mux_h I__4387 (
            .O(N__22304),
            .I(N__22297));
    LocalMux I__4386 (
            .O(N__22301),
            .I(N__22294));
    InMux I__4385 (
            .O(N__22300),
            .I(N__22291));
    Span4Mux_h I__4384 (
            .O(N__22297),
            .I(N__22288));
    Span4Mux_h I__4383 (
            .O(N__22294),
            .I(N__22285));
    LocalMux I__4382 (
            .O(N__22291),
            .I(data_in_3_1));
    Odrv4 I__4381 (
            .O(N__22288),
            .I(data_in_3_1));
    Odrv4 I__4380 (
            .O(N__22285),
            .I(data_in_3_1));
    CascadeMux I__4379 (
            .O(N__22278),
            .I(N__22275));
    InMux I__4378 (
            .O(N__22275),
            .I(N__22271));
    InMux I__4377 (
            .O(N__22274),
            .I(N__22268));
    LocalMux I__4376 (
            .O(N__22271),
            .I(N__22265));
    LocalMux I__4375 (
            .O(N__22268),
            .I(N__22261));
    Span4Mux_v I__4374 (
            .O(N__22265),
            .I(N__22258));
    InMux I__4373 (
            .O(N__22264),
            .I(N__22255));
    Span4Mux_v I__4372 (
            .O(N__22261),
            .I(N__22252));
    Span4Mux_h I__4371 (
            .O(N__22258),
            .I(N__22249));
    LocalMux I__4370 (
            .O(N__22255),
            .I(data_in_0_0));
    Odrv4 I__4369 (
            .O(N__22252),
            .I(data_in_0_0));
    Odrv4 I__4368 (
            .O(N__22249),
            .I(data_in_0_0));
    InMux I__4367 (
            .O(N__22242),
            .I(N__22239));
    LocalMux I__4366 (
            .O(N__22239),
            .I(N__22236));
    Span4Mux_s3_h I__4365 (
            .O(N__22236),
            .I(N__22232));
    InMux I__4364 (
            .O(N__22235),
            .I(N__22229));
    Span4Mux_h I__4363 (
            .O(N__22232),
            .I(N__22223));
    LocalMux I__4362 (
            .O(N__22229),
            .I(N__22223));
    InMux I__4361 (
            .O(N__22228),
            .I(N__22219));
    Span4Mux_v I__4360 (
            .O(N__22223),
            .I(N__22216));
    InMux I__4359 (
            .O(N__22222),
            .I(N__22213));
    LocalMux I__4358 (
            .O(N__22219),
            .I(\c0.data_in_field_0 ));
    Odrv4 I__4357 (
            .O(N__22216),
            .I(\c0.data_in_field_0 ));
    LocalMux I__4356 (
            .O(N__22213),
            .I(\c0.data_in_field_0 ));
    InMux I__4355 (
            .O(N__22206),
            .I(N__22203));
    LocalMux I__4354 (
            .O(N__22203),
            .I(N__22199));
    InMux I__4353 (
            .O(N__22202),
            .I(N__22196));
    Span4Mux_v I__4352 (
            .O(N__22199),
            .I(N__22189));
    LocalMux I__4351 (
            .O(N__22196),
            .I(N__22189));
    InMux I__4350 (
            .O(N__22195),
            .I(N__22183));
    InMux I__4349 (
            .O(N__22194),
            .I(N__22183));
    Span4Mux_v I__4348 (
            .O(N__22189),
            .I(N__22180));
    InMux I__4347 (
            .O(N__22188),
            .I(N__22177));
    LocalMux I__4346 (
            .O(N__22183),
            .I(\c0.data_in_field_117 ));
    Odrv4 I__4345 (
            .O(N__22180),
            .I(\c0.data_in_field_117 ));
    LocalMux I__4344 (
            .O(N__22177),
            .I(\c0.data_in_field_117 ));
    InMux I__4343 (
            .O(N__22170),
            .I(N__22167));
    LocalMux I__4342 (
            .O(N__22167),
            .I(N__22163));
    InMux I__4341 (
            .O(N__22166),
            .I(N__22160));
    Odrv4 I__4340 (
            .O(N__22163),
            .I(\c0.n1855 ));
    LocalMux I__4339 (
            .O(N__22160),
            .I(\c0.n1855 ));
    InMux I__4338 (
            .O(N__22155),
            .I(N__22152));
    LocalMux I__4337 (
            .O(N__22152),
            .I(N__22149));
    Span12Mux_v I__4336 (
            .O(N__22149),
            .I(N__22146));
    Odrv12 I__4335 (
            .O(N__22146),
            .I(\c0.n13 ));
    CascadeMux I__4334 (
            .O(N__22143),
            .I(\c0.n12_adj_1898_cascade_ ));
    InMux I__4333 (
            .O(N__22140),
            .I(N__22137));
    LocalMux I__4332 (
            .O(N__22137),
            .I(\c0.tx.n5885 ));
    InMux I__4331 (
            .O(N__22134),
            .I(N__22130));
    InMux I__4330 (
            .O(N__22133),
            .I(N__22127));
    LocalMux I__4329 (
            .O(N__22130),
            .I(\c0.tx.n15 ));
    LocalMux I__4328 (
            .O(N__22127),
            .I(\c0.tx.n15 ));
    InMux I__4327 (
            .O(N__22122),
            .I(N__22119));
    LocalMux I__4326 (
            .O(N__22119),
            .I(\c0.tx.n5884 ));
    InMux I__4325 (
            .O(N__22116),
            .I(N__22112));
    InMux I__4324 (
            .O(N__22115),
            .I(N__22109));
    LocalMux I__4323 (
            .O(N__22112),
            .I(N__22105));
    LocalMux I__4322 (
            .O(N__22109),
            .I(N__22102));
    InMux I__4321 (
            .O(N__22108),
            .I(N__22099));
    Odrv4 I__4320 (
            .O(N__22105),
            .I(data_in_4_3));
    Odrv12 I__4319 (
            .O(N__22102),
            .I(data_in_4_3));
    LocalMux I__4318 (
            .O(N__22099),
            .I(data_in_4_3));
    InMux I__4317 (
            .O(N__22092),
            .I(N__22088));
    InMux I__4316 (
            .O(N__22091),
            .I(N__22084));
    LocalMux I__4315 (
            .O(N__22088),
            .I(N__22081));
    InMux I__4314 (
            .O(N__22087),
            .I(N__22078));
    LocalMux I__4313 (
            .O(N__22084),
            .I(N__22074));
    Span4Mux_v I__4312 (
            .O(N__22081),
            .I(N__22069));
    LocalMux I__4311 (
            .O(N__22078),
            .I(N__22069));
    InMux I__4310 (
            .O(N__22077),
            .I(N__22066));
    Span4Mux_v I__4309 (
            .O(N__22074),
            .I(N__22063));
    Odrv4 I__4308 (
            .O(N__22069),
            .I(data_in_3_3));
    LocalMux I__4307 (
            .O(N__22066),
            .I(data_in_3_3));
    Odrv4 I__4306 (
            .O(N__22063),
            .I(data_in_3_3));
    InMux I__4305 (
            .O(N__22056),
            .I(N__22051));
    InMux I__4304 (
            .O(N__22055),
            .I(N__22048));
    InMux I__4303 (
            .O(N__22054),
            .I(N__22045));
    LocalMux I__4302 (
            .O(N__22051),
            .I(N__22041));
    LocalMux I__4301 (
            .O(N__22048),
            .I(N__22038));
    LocalMux I__4300 (
            .O(N__22045),
            .I(N__22035));
    InMux I__4299 (
            .O(N__22044),
            .I(N__22032));
    Span4Mux_h I__4298 (
            .O(N__22041),
            .I(N__22027));
    Span4Mux_v I__4297 (
            .O(N__22038),
            .I(N__22027));
    Odrv4 I__4296 (
            .O(N__22035),
            .I(data_in_2_2));
    LocalMux I__4295 (
            .O(N__22032),
            .I(data_in_2_2));
    Odrv4 I__4294 (
            .O(N__22027),
            .I(data_in_2_2));
    InMux I__4293 (
            .O(N__22020),
            .I(N__22016));
    InMux I__4292 (
            .O(N__22019),
            .I(N__22013));
    LocalMux I__4291 (
            .O(N__22016),
            .I(N__22010));
    LocalMux I__4290 (
            .O(N__22013),
            .I(N__22007));
    Span4Mux_v I__4289 (
            .O(N__22010),
            .I(N__22002));
    Span4Mux_h I__4288 (
            .O(N__22007),
            .I(N__21999));
    InMux I__4287 (
            .O(N__22006),
            .I(N__21996));
    InMux I__4286 (
            .O(N__22005),
            .I(N__21993));
    Odrv4 I__4285 (
            .O(N__22002),
            .I(data_in_1_2));
    Odrv4 I__4284 (
            .O(N__21999),
            .I(data_in_1_2));
    LocalMux I__4283 (
            .O(N__21996),
            .I(data_in_1_2));
    LocalMux I__4282 (
            .O(N__21993),
            .I(data_in_1_2));
    InMux I__4281 (
            .O(N__21984),
            .I(N__21979));
    InMux I__4280 (
            .O(N__21983),
            .I(N__21976));
    CascadeMux I__4279 (
            .O(N__21982),
            .I(N__21971));
    LocalMux I__4278 (
            .O(N__21979),
            .I(N__21968));
    LocalMux I__4277 (
            .O(N__21976),
            .I(N__21965));
    InMux I__4276 (
            .O(N__21975),
            .I(N__21962));
    InMux I__4275 (
            .O(N__21974),
            .I(N__21959));
    InMux I__4274 (
            .O(N__21971),
            .I(N__21956));
    Span12Mux_s5_h I__4273 (
            .O(N__21968),
            .I(N__21953));
    Span4Mux_h I__4272 (
            .O(N__21965),
            .I(N__21950));
    LocalMux I__4271 (
            .O(N__21962),
            .I(N__21945));
    LocalMux I__4270 (
            .O(N__21959),
            .I(N__21945));
    LocalMux I__4269 (
            .O(N__21956),
            .I(\c0.data_in_field_80 ));
    Odrv12 I__4268 (
            .O(N__21953),
            .I(\c0.data_in_field_80 ));
    Odrv4 I__4267 (
            .O(N__21950),
            .I(\c0.data_in_field_80 ));
    Odrv4 I__4266 (
            .O(N__21945),
            .I(\c0.data_in_field_80 ));
    CascadeMux I__4265 (
            .O(N__21936),
            .I(\c0.n42_cascade_ ));
    InMux I__4264 (
            .O(N__21933),
            .I(N__21930));
    LocalMux I__4263 (
            .O(N__21930),
            .I(N__21927));
    Span4Mux_v I__4262 (
            .O(N__21927),
            .I(N__21924));
    Span4Mux_h I__4261 (
            .O(N__21924),
            .I(N__21921));
    Span4Mux_h I__4260 (
            .O(N__21921),
            .I(N__21918));
    Odrv4 I__4259 (
            .O(N__21918),
            .I(\c0.n48 ));
    CascadeMux I__4258 (
            .O(N__21915),
            .I(N__21911));
    InMux I__4257 (
            .O(N__21914),
            .I(N__21907));
    InMux I__4256 (
            .O(N__21911),
            .I(N__21904));
    InMux I__4255 (
            .O(N__21910),
            .I(N__21901));
    LocalMux I__4254 (
            .O(N__21907),
            .I(N__21896));
    LocalMux I__4253 (
            .O(N__21904),
            .I(N__21896));
    LocalMux I__4252 (
            .O(N__21901),
            .I(N__21892));
    Span4Mux_v I__4251 (
            .O(N__21896),
            .I(N__21889));
    InMux I__4250 (
            .O(N__21895),
            .I(N__21886));
    Span4Mux_h I__4249 (
            .O(N__21892),
            .I(N__21881));
    Span4Mux_v I__4248 (
            .O(N__21889),
            .I(N__21881));
    LocalMux I__4247 (
            .O(N__21886),
            .I(data_in_19_0));
    Odrv4 I__4246 (
            .O(N__21881),
            .I(data_in_19_0));
    CascadeMux I__4245 (
            .O(N__21876),
            .I(N__21873));
    InMux I__4244 (
            .O(N__21873),
            .I(N__21869));
    InMux I__4243 (
            .O(N__21872),
            .I(N__21866));
    LocalMux I__4242 (
            .O(N__21869),
            .I(N__21863));
    LocalMux I__4241 (
            .O(N__21866),
            .I(N__21860));
    Span4Mux_v I__4240 (
            .O(N__21863),
            .I(N__21857));
    Span4Mux_s3_h I__4239 (
            .O(N__21860),
            .I(N__21854));
    Span4Mux_v I__4238 (
            .O(N__21857),
            .I(N__21848));
    Span4Mux_h I__4237 (
            .O(N__21854),
            .I(N__21848));
    InMux I__4236 (
            .O(N__21853),
            .I(N__21845));
    Odrv4 I__4235 (
            .O(N__21848),
            .I(data_in_15_7));
    LocalMux I__4234 (
            .O(N__21845),
            .I(data_in_15_7));
    InMux I__4233 (
            .O(N__21840),
            .I(bfn_9_27_0_));
    InMux I__4232 (
            .O(N__21837),
            .I(\c0.tx.n4764 ));
    InMux I__4231 (
            .O(N__21834),
            .I(\c0.tx.n4765 ));
    InMux I__4230 (
            .O(N__21831),
            .I(\c0.tx.n4766 ));
    InMux I__4229 (
            .O(N__21828),
            .I(\c0.tx.n4767 ));
    InMux I__4228 (
            .O(N__21825),
            .I(\c0.tx.n4768 ));
    InMux I__4227 (
            .O(N__21822),
            .I(\c0.tx.n4769 ));
    InMux I__4226 (
            .O(N__21819),
            .I(\c0.tx.n4770 ));
    InMux I__4225 (
            .O(N__21816),
            .I(bfn_9_28_0_));
    InMux I__4224 (
            .O(N__21813),
            .I(N__21810));
    LocalMux I__4223 (
            .O(N__21810),
            .I(N__21805));
    InMux I__4222 (
            .O(N__21809),
            .I(N__21802));
    InMux I__4221 (
            .O(N__21808),
            .I(N__21799));
    Span4Mux_v I__4220 (
            .O(N__21805),
            .I(N__21790));
    LocalMux I__4219 (
            .O(N__21802),
            .I(N__21790));
    LocalMux I__4218 (
            .O(N__21799),
            .I(N__21790));
    CascadeMux I__4217 (
            .O(N__21798),
            .I(N__21787));
    InMux I__4216 (
            .O(N__21797),
            .I(N__21784));
    Span4Mux_v I__4215 (
            .O(N__21790),
            .I(N__21781));
    InMux I__4214 (
            .O(N__21787),
            .I(N__21778));
    LocalMux I__4213 (
            .O(N__21784),
            .I(\c0.data_in_field_4 ));
    Odrv4 I__4212 (
            .O(N__21781),
            .I(\c0.data_in_field_4 ));
    LocalMux I__4211 (
            .O(N__21778),
            .I(\c0.data_in_field_4 ));
    InMux I__4210 (
            .O(N__21771),
            .I(N__21766));
    InMux I__4209 (
            .O(N__21770),
            .I(N__21762));
    InMux I__4208 (
            .O(N__21769),
            .I(N__21759));
    LocalMux I__4207 (
            .O(N__21766),
            .I(N__21756));
    CascadeMux I__4206 (
            .O(N__21765),
            .I(N__21753));
    LocalMux I__4205 (
            .O(N__21762),
            .I(N__21750));
    LocalMux I__4204 (
            .O(N__21759),
            .I(N__21747));
    Span4Mux_h I__4203 (
            .O(N__21756),
            .I(N__21744));
    InMux I__4202 (
            .O(N__21753),
            .I(N__21740));
    Span4Mux_v I__4201 (
            .O(N__21750),
            .I(N__21737));
    Span4Mux_v I__4200 (
            .O(N__21747),
            .I(N__21734));
    Span4Mux_h I__4199 (
            .O(N__21744),
            .I(N__21731));
    InMux I__4198 (
            .O(N__21743),
            .I(N__21728));
    LocalMux I__4197 (
            .O(N__21740),
            .I(\c0.data_in_field_12 ));
    Odrv4 I__4196 (
            .O(N__21737),
            .I(\c0.data_in_field_12 ));
    Odrv4 I__4195 (
            .O(N__21734),
            .I(\c0.data_in_field_12 ));
    Odrv4 I__4194 (
            .O(N__21731),
            .I(\c0.data_in_field_12 ));
    LocalMux I__4193 (
            .O(N__21728),
            .I(\c0.data_in_field_12 ));
    InMux I__4192 (
            .O(N__21717),
            .I(N__21714));
    LocalMux I__4191 (
            .O(N__21714),
            .I(N__21711));
    Span4Mux_h I__4190 (
            .O(N__21711),
            .I(N__21708));
    Span4Mux_h I__4189 (
            .O(N__21708),
            .I(N__21705));
    Odrv4 I__4188 (
            .O(N__21705),
            .I(\c0.n5722 ));
    CascadeMux I__4187 (
            .O(N__21702),
            .I(\c0.tx.n3631_cascade_ ));
    InMux I__4186 (
            .O(N__21699),
            .I(N__21694));
    CascadeMux I__4185 (
            .O(N__21698),
            .I(N__21690));
    InMux I__4184 (
            .O(N__21697),
            .I(N__21687));
    LocalMux I__4183 (
            .O(N__21694),
            .I(N__21684));
    InMux I__4182 (
            .O(N__21693),
            .I(N__21681));
    InMux I__4181 (
            .O(N__21690),
            .I(N__21677));
    LocalMux I__4180 (
            .O(N__21687),
            .I(N__21674));
    Span4Mux_v I__4179 (
            .O(N__21684),
            .I(N__21669));
    LocalMux I__4178 (
            .O(N__21681),
            .I(N__21669));
    InMux I__4177 (
            .O(N__21680),
            .I(N__21666));
    LocalMux I__4176 (
            .O(N__21677),
            .I(\c0.data_in_field_20 ));
    Odrv12 I__4175 (
            .O(N__21674),
            .I(\c0.data_in_field_20 ));
    Odrv4 I__4174 (
            .O(N__21669),
            .I(\c0.data_in_field_20 ));
    LocalMux I__4173 (
            .O(N__21666),
            .I(\c0.data_in_field_20 ));
    CascadeMux I__4172 (
            .O(N__21657),
            .I(N__21654));
    InMux I__4171 (
            .O(N__21654),
            .I(N__21651));
    LocalMux I__4170 (
            .O(N__21651),
            .I(\c0.n6189 ));
    CascadeMux I__4169 (
            .O(N__21648),
            .I(\c0.tx.n5812_cascade_ ));
    CascadeMux I__4168 (
            .O(N__21645),
            .I(\c0.tx.n14_cascade_ ));
    InMux I__4167 (
            .O(N__21642),
            .I(N__21639));
    LocalMux I__4166 (
            .O(N__21639),
            .I(N__21635));
    InMux I__4165 (
            .O(N__21638),
            .I(N__21632));
    Span4Mux_h I__4164 (
            .O(N__21635),
            .I(N__21629));
    LocalMux I__4163 (
            .O(N__21632),
            .I(r_Tx_Data_7));
    Odrv4 I__4162 (
            .O(N__21629),
            .I(r_Tx_Data_7));
    InMux I__4161 (
            .O(N__21624),
            .I(N__21620));
    InMux I__4160 (
            .O(N__21623),
            .I(N__21617));
    LocalMux I__4159 (
            .O(N__21620),
            .I(r_Tx_Data_6));
    LocalMux I__4158 (
            .O(N__21617),
            .I(r_Tx_Data_6));
    InMux I__4157 (
            .O(N__21612),
            .I(\c0.n4759 ));
    InMux I__4156 (
            .O(N__21609),
            .I(\c0.n4760 ));
    InMux I__4155 (
            .O(N__21606),
            .I(bfn_9_24_0_));
    InMux I__4154 (
            .O(N__21603),
            .I(\c0.n4762 ));
    InMux I__4153 (
            .O(N__21600),
            .I(\c0.n4763 ));
    InMux I__4152 (
            .O(N__21597),
            .I(N__21593));
    InMux I__4151 (
            .O(N__21596),
            .I(N__21590));
    LocalMux I__4150 (
            .O(N__21593),
            .I(\c0.delay_counter_1 ));
    LocalMux I__4149 (
            .O(N__21590),
            .I(\c0.delay_counter_1 ));
    InMux I__4148 (
            .O(N__21585),
            .I(N__21581));
    InMux I__4147 (
            .O(N__21584),
            .I(N__21578));
    LocalMux I__4146 (
            .O(N__21581),
            .I(\c0.delay_counter_5 ));
    LocalMux I__4145 (
            .O(N__21578),
            .I(\c0.delay_counter_5 ));
    InMux I__4144 (
            .O(N__21573),
            .I(N__21569));
    CascadeMux I__4143 (
            .O(N__21572),
            .I(N__21565));
    LocalMux I__4142 (
            .O(N__21569),
            .I(N__21562));
    CascadeMux I__4141 (
            .O(N__21568),
            .I(N__21559));
    InMux I__4140 (
            .O(N__21565),
            .I(N__21556));
    Span4Mux_h I__4139 (
            .O(N__21562),
            .I(N__21553));
    InMux I__4138 (
            .O(N__21559),
            .I(N__21550));
    LocalMux I__4137 (
            .O(N__21556),
            .I(\c0.data_in_field_116 ));
    Odrv4 I__4136 (
            .O(N__21553),
            .I(\c0.data_in_field_116 ));
    LocalMux I__4135 (
            .O(N__21550),
            .I(\c0.data_in_field_116 ));
    InMux I__4134 (
            .O(N__21543),
            .I(N__21540));
    LocalMux I__4133 (
            .O(N__21540),
            .I(N__21534));
    InMux I__4132 (
            .O(N__21539),
            .I(N__21529));
    InMux I__4131 (
            .O(N__21538),
            .I(N__21529));
    InMux I__4130 (
            .O(N__21537),
            .I(N__21524));
    Span4Mux_h I__4129 (
            .O(N__21534),
            .I(N__21521));
    LocalMux I__4128 (
            .O(N__21529),
            .I(N__21518));
    InMux I__4127 (
            .O(N__21528),
            .I(N__21513));
    InMux I__4126 (
            .O(N__21527),
            .I(N__21513));
    LocalMux I__4125 (
            .O(N__21524),
            .I(\c0.data_in_field_124 ));
    Odrv4 I__4124 (
            .O(N__21521),
            .I(\c0.data_in_field_124 ));
    Odrv12 I__4123 (
            .O(N__21518),
            .I(\c0.data_in_field_124 ));
    LocalMux I__4122 (
            .O(N__21513),
            .I(\c0.data_in_field_124 ));
    CascadeMux I__4121 (
            .O(N__21504),
            .I(\c0.n6171_cascade_ ));
    InMux I__4120 (
            .O(N__21501),
            .I(N__21498));
    LocalMux I__4119 (
            .O(N__21498),
            .I(N__21495));
    Span4Mux_h I__4118 (
            .O(N__21495),
            .I(N__21492));
    Span4Mux_h I__4117 (
            .O(N__21492),
            .I(N__21489));
    Odrv4 I__4116 (
            .O(N__21489),
            .I(\c0.n5731 ));
    InMux I__4115 (
            .O(N__21486),
            .I(N__21482));
    InMux I__4114 (
            .O(N__21485),
            .I(N__21479));
    LocalMux I__4113 (
            .O(N__21482),
            .I(N__21475));
    LocalMux I__4112 (
            .O(N__21479),
            .I(N__21472));
    InMux I__4111 (
            .O(N__21478),
            .I(N__21468));
    Span4Mux_h I__4110 (
            .O(N__21475),
            .I(N__21465));
    Span4Mux_v I__4109 (
            .O(N__21472),
            .I(N__21462));
    InMux I__4108 (
            .O(N__21471),
            .I(N__21459));
    LocalMux I__4107 (
            .O(N__21468),
            .I(N__21456));
    Odrv4 I__4106 (
            .O(N__21465),
            .I(data_in_3_2));
    Odrv4 I__4105 (
            .O(N__21462),
            .I(data_in_3_2));
    LocalMux I__4104 (
            .O(N__21459),
            .I(data_in_3_2));
    Odrv4 I__4103 (
            .O(N__21456),
            .I(data_in_3_2));
    InMux I__4102 (
            .O(N__21447),
            .I(N__21444));
    LocalMux I__4101 (
            .O(N__21444),
            .I(N__21441));
    Span4Mux_h I__4100 (
            .O(N__21441),
            .I(N__21437));
    InMux I__4099 (
            .O(N__21440),
            .I(N__21434));
    Span4Mux_h I__4098 (
            .O(N__21437),
            .I(N__21431));
    LocalMux I__4097 (
            .O(N__21434),
            .I(N__21428));
    Odrv4 I__4096 (
            .O(N__21431),
            .I(\c0.n1955 ));
    Odrv4 I__4095 (
            .O(N__21428),
            .I(\c0.n1955 ));
    CascadeMux I__4094 (
            .O(N__21423),
            .I(N__21420));
    InMux I__4093 (
            .O(N__21420),
            .I(N__21417));
    LocalMux I__4092 (
            .O(N__21417),
            .I(N__21414));
    Span4Mux_v I__4091 (
            .O(N__21414),
            .I(N__21409));
    InMux I__4090 (
            .O(N__21413),
            .I(N__21404));
    InMux I__4089 (
            .O(N__21412),
            .I(N__21404));
    Odrv4 I__4088 (
            .O(N__21409),
            .I(data_in_4_2));
    LocalMux I__4087 (
            .O(N__21404),
            .I(data_in_4_2));
    CascadeMux I__4086 (
            .O(N__21399),
            .I(N__21396));
    InMux I__4085 (
            .O(N__21396),
            .I(N__21392));
    InMux I__4084 (
            .O(N__21395),
            .I(N__21388));
    LocalMux I__4083 (
            .O(N__21392),
            .I(N__21385));
    InMux I__4082 (
            .O(N__21391),
            .I(N__21382));
    LocalMux I__4081 (
            .O(N__21388),
            .I(N__21378));
    Span4Mux_v I__4080 (
            .O(N__21385),
            .I(N__21375));
    LocalMux I__4079 (
            .O(N__21382),
            .I(N__21372));
    InMux I__4078 (
            .O(N__21381),
            .I(N__21369));
    Span4Mux_h I__4077 (
            .O(N__21378),
            .I(N__21366));
    Sp12to4 I__4076 (
            .O(N__21375),
            .I(N__21361));
    Span12Mux_v I__4075 (
            .O(N__21372),
            .I(N__21361));
    LocalMux I__4074 (
            .O(N__21369),
            .I(data_in_18_5));
    Odrv4 I__4073 (
            .O(N__21366),
            .I(data_in_18_5));
    Odrv12 I__4072 (
            .O(N__21361),
            .I(data_in_18_5));
    CascadeMux I__4071 (
            .O(N__21354),
            .I(N__21351));
    InMux I__4070 (
            .O(N__21351),
            .I(N__21348));
    LocalMux I__4069 (
            .O(N__21348),
            .I(N__21344));
    InMux I__4068 (
            .O(N__21347),
            .I(N__21341));
    Span4Mux_v I__4067 (
            .O(N__21344),
            .I(N__21337));
    LocalMux I__4066 (
            .O(N__21341),
            .I(N__21334));
    InMux I__4065 (
            .O(N__21340),
            .I(N__21331));
    Odrv4 I__4064 (
            .O(N__21337),
            .I(data_in_17_5));
    Odrv12 I__4063 (
            .O(N__21334),
            .I(data_in_17_5));
    LocalMux I__4062 (
            .O(N__21331),
            .I(data_in_17_5));
    InMux I__4061 (
            .O(N__21324),
            .I(\c0.n4754 ));
    InMux I__4060 (
            .O(N__21321),
            .I(\c0.n4755 ));
    InMux I__4059 (
            .O(N__21318),
            .I(\c0.n4756 ));
    InMux I__4058 (
            .O(N__21315),
            .I(\c0.n4757 ));
    InMux I__4057 (
            .O(N__21312),
            .I(\c0.n4758 ));
    InMux I__4056 (
            .O(N__21309),
            .I(N__21305));
    InMux I__4055 (
            .O(N__21308),
            .I(N__21302));
    LocalMux I__4054 (
            .O(N__21305),
            .I(N__21299));
    LocalMux I__4053 (
            .O(N__21302),
            .I(N__21296));
    Span4Mux_v I__4052 (
            .O(N__21299),
            .I(N__21293));
    Span4Mux_v I__4051 (
            .O(N__21296),
            .I(N__21290));
    Span4Mux_h I__4050 (
            .O(N__21293),
            .I(N__21286));
    Span4Mux_v I__4049 (
            .O(N__21290),
            .I(N__21283));
    InMux I__4048 (
            .O(N__21289),
            .I(N__21280));
    Odrv4 I__4047 (
            .O(N__21286),
            .I(data_in_15_5));
    Odrv4 I__4046 (
            .O(N__21283),
            .I(data_in_15_5));
    LocalMux I__4045 (
            .O(N__21280),
            .I(data_in_15_5));
    InMux I__4044 (
            .O(N__21273),
            .I(N__21270));
    LocalMux I__4043 (
            .O(N__21270),
            .I(\c0.n6414 ));
    InMux I__4042 (
            .O(N__21267),
            .I(N__21264));
    LocalMux I__4041 (
            .O(N__21264),
            .I(N__21261));
    Odrv4 I__4040 (
            .O(N__21261),
            .I(\c0.n5563 ));
    CascadeMux I__4039 (
            .O(N__21258),
            .I(N__21255));
    InMux I__4038 (
            .O(N__21255),
            .I(N__21252));
    LocalMux I__4037 (
            .O(N__21252),
            .I(N__21249));
    Span4Mux_v I__4036 (
            .O(N__21249),
            .I(N__21245));
    InMux I__4035 (
            .O(N__21248),
            .I(N__21242));
    Span4Mux_h I__4034 (
            .O(N__21245),
            .I(N__21236));
    LocalMux I__4033 (
            .O(N__21242),
            .I(N__21236));
    InMux I__4032 (
            .O(N__21241),
            .I(N__21233));
    Odrv4 I__4031 (
            .O(N__21236),
            .I(data_in_11_1));
    LocalMux I__4030 (
            .O(N__21233),
            .I(data_in_11_1));
    InMux I__4029 (
            .O(N__21228),
            .I(N__21224));
    CascadeMux I__4028 (
            .O(N__21227),
            .I(N__21221));
    LocalMux I__4027 (
            .O(N__21224),
            .I(N__21218));
    InMux I__4026 (
            .O(N__21221),
            .I(N__21215));
    Span4Mux_v I__4025 (
            .O(N__21218),
            .I(N__21212));
    LocalMux I__4024 (
            .O(N__21215),
            .I(N__21206));
    Span4Mux_h I__4023 (
            .O(N__21212),
            .I(N__21203));
    InMux I__4022 (
            .O(N__21211),
            .I(N__21200));
    InMux I__4021 (
            .O(N__21210),
            .I(N__21195));
    InMux I__4020 (
            .O(N__21209),
            .I(N__21195));
    Span4Mux_h I__4019 (
            .O(N__21206),
            .I(N__21192));
    Odrv4 I__4018 (
            .O(N__21203),
            .I(\c0.data_in_field_45 ));
    LocalMux I__4017 (
            .O(N__21200),
            .I(\c0.data_in_field_45 ));
    LocalMux I__4016 (
            .O(N__21195),
            .I(\c0.data_in_field_45 ));
    Odrv4 I__4015 (
            .O(N__21192),
            .I(\c0.data_in_field_45 ));
    InMux I__4014 (
            .O(N__21183),
            .I(N__21180));
    LocalMux I__4013 (
            .O(N__21180),
            .I(N__21175));
    InMux I__4012 (
            .O(N__21179),
            .I(N__21172));
    InMux I__4011 (
            .O(N__21178),
            .I(N__21169));
    Span4Mux_v I__4010 (
            .O(N__21175),
            .I(N__21164));
    LocalMux I__4009 (
            .O(N__21172),
            .I(N__21164));
    LocalMux I__4008 (
            .O(N__21169),
            .I(N__21161));
    Odrv4 I__4007 (
            .O(N__21164),
            .I(\c0.n2065 ));
    Odrv4 I__4006 (
            .O(N__21161),
            .I(\c0.n2065 ));
    InMux I__4005 (
            .O(N__21156),
            .I(N__21153));
    LocalMux I__4004 (
            .O(N__21153),
            .I(\c0.n18 ));
    CascadeMux I__4003 (
            .O(N__21150),
            .I(\c0.n2149_cascade_ ));
    InMux I__4002 (
            .O(N__21147),
            .I(N__21144));
    LocalMux I__4001 (
            .O(N__21144),
            .I(N__21141));
    Span12Mux_v I__4000 (
            .O(N__21141),
            .I(N__21138));
    Odrv12 I__3999 (
            .O(N__21138),
            .I(\c0.n21 ));
    CascadeMux I__3998 (
            .O(N__21135),
            .I(N__21132));
    InMux I__3997 (
            .O(N__21132),
            .I(N__21129));
    LocalMux I__3996 (
            .O(N__21129),
            .I(N__21124));
    InMux I__3995 (
            .O(N__21128),
            .I(N__21121));
    InMux I__3994 (
            .O(N__21127),
            .I(N__21118));
    Odrv12 I__3993 (
            .O(N__21124),
            .I(data_in_17_3));
    LocalMux I__3992 (
            .O(N__21121),
            .I(data_in_17_3));
    LocalMux I__3991 (
            .O(N__21118),
            .I(data_in_17_3));
    CascadeMux I__3990 (
            .O(N__21111),
            .I(N__21108));
    InMux I__3989 (
            .O(N__21108),
            .I(N__21105));
    LocalMux I__3988 (
            .O(N__21105),
            .I(N__21102));
    Span4Mux_v I__3987 (
            .O(N__21102),
            .I(N__21096));
    InMux I__3986 (
            .O(N__21101),
            .I(N__21093));
    InMux I__3985 (
            .O(N__21100),
            .I(N__21088));
    InMux I__3984 (
            .O(N__21099),
            .I(N__21088));
    Odrv4 I__3983 (
            .O(N__21096),
            .I(data_in_2_3));
    LocalMux I__3982 (
            .O(N__21093),
            .I(data_in_2_3));
    LocalMux I__3981 (
            .O(N__21088),
            .I(data_in_2_3));
    InMux I__3980 (
            .O(N__21081),
            .I(N__21077));
    CascadeMux I__3979 (
            .O(N__21080),
            .I(N__21074));
    LocalMux I__3978 (
            .O(N__21077),
            .I(N__21071));
    InMux I__3977 (
            .O(N__21074),
            .I(N__21067));
    Span4Mux_v I__3976 (
            .O(N__21071),
            .I(N__21064));
    InMux I__3975 (
            .O(N__21070),
            .I(N__21061));
    LocalMux I__3974 (
            .O(N__21067),
            .I(N__21056));
    Span4Mux_h I__3973 (
            .O(N__21064),
            .I(N__21056));
    LocalMux I__3972 (
            .O(N__21061),
            .I(data_in_6_7));
    Odrv4 I__3971 (
            .O(N__21056),
            .I(data_in_6_7));
    CascadeMux I__3970 (
            .O(N__21051),
            .I(N__21048));
    InMux I__3969 (
            .O(N__21048),
            .I(N__21045));
    LocalMux I__3968 (
            .O(N__21045),
            .I(N__21041));
    InMux I__3967 (
            .O(N__21044),
            .I(N__21038));
    Span4Mux_v I__3966 (
            .O(N__21041),
            .I(N__21033));
    LocalMux I__3965 (
            .O(N__21038),
            .I(N__21033));
    Span4Mux_h I__3964 (
            .O(N__21033),
            .I(N__21029));
    CascadeMux I__3963 (
            .O(N__21032),
            .I(N__21026));
    Span4Mux_h I__3962 (
            .O(N__21029),
            .I(N__21023));
    InMux I__3961 (
            .O(N__21026),
            .I(N__21020));
    Odrv4 I__3960 (
            .O(N__21023),
            .I(data_in_6_5));
    LocalMux I__3959 (
            .O(N__21020),
            .I(data_in_6_5));
    InMux I__3958 (
            .O(N__21015),
            .I(N__21012));
    LocalMux I__3957 (
            .O(N__21012),
            .I(N__21009));
    Span4Mux_h I__3956 (
            .O(N__21009),
            .I(N__21006));
    Odrv4 I__3955 (
            .O(N__21006),
            .I(\c0.n25_adj_1948 ));
    InMux I__3954 (
            .O(N__21003),
            .I(N__20997));
    InMux I__3953 (
            .O(N__21002),
            .I(N__20994));
    InMux I__3952 (
            .O(N__21001),
            .I(N__20991));
    InMux I__3951 (
            .O(N__21000),
            .I(N__20988));
    LocalMux I__3950 (
            .O(N__20997),
            .I(N__20985));
    LocalMux I__3949 (
            .O(N__20994),
            .I(N__20982));
    LocalMux I__3948 (
            .O(N__20991),
            .I(N__20979));
    LocalMux I__3947 (
            .O(N__20988),
            .I(N__20968));
    Span4Mux_v I__3946 (
            .O(N__20985),
            .I(N__20968));
    Span4Mux_v I__3945 (
            .O(N__20982),
            .I(N__20968));
    Span4Mux_h I__3944 (
            .O(N__20979),
            .I(N__20968));
    InMux I__3943 (
            .O(N__20978),
            .I(N__20963));
    InMux I__3942 (
            .O(N__20977),
            .I(N__20963));
    Odrv4 I__3941 (
            .O(N__20968),
            .I(\c0.data_in_field_94 ));
    LocalMux I__3940 (
            .O(N__20963),
            .I(\c0.data_in_field_94 ));
    InMux I__3939 (
            .O(N__20958),
            .I(N__20955));
    LocalMux I__3938 (
            .O(N__20955),
            .I(N__20952));
    Span4Mux_v I__3937 (
            .O(N__20952),
            .I(N__20947));
    InMux I__3936 (
            .O(N__20951),
            .I(N__20944));
    InMux I__3935 (
            .O(N__20950),
            .I(N__20940));
    Span4Mux_h I__3934 (
            .O(N__20947),
            .I(N__20935));
    LocalMux I__3933 (
            .O(N__20944),
            .I(N__20935));
    InMux I__3932 (
            .O(N__20943),
            .I(N__20932));
    LocalMux I__3931 (
            .O(N__20940),
            .I(\c0.data_in_field_66 ));
    Odrv4 I__3930 (
            .O(N__20935),
            .I(\c0.data_in_field_66 ));
    LocalMux I__3929 (
            .O(N__20932),
            .I(\c0.data_in_field_66 ));
    CascadeMux I__3928 (
            .O(N__20925),
            .I(N__20920));
    InMux I__3927 (
            .O(N__20924),
            .I(N__20917));
    InMux I__3926 (
            .O(N__20923),
            .I(N__20914));
    InMux I__3925 (
            .O(N__20920),
            .I(N__20910));
    LocalMux I__3924 (
            .O(N__20917),
            .I(N__20907));
    LocalMux I__3923 (
            .O(N__20914),
            .I(N__20904));
    InMux I__3922 (
            .O(N__20913),
            .I(N__20901));
    LocalMux I__3921 (
            .O(N__20910),
            .I(\c0.data_in_field_79 ));
    Odrv4 I__3920 (
            .O(N__20907),
            .I(\c0.data_in_field_79 ));
    Odrv12 I__3919 (
            .O(N__20904),
            .I(\c0.data_in_field_79 ));
    LocalMux I__3918 (
            .O(N__20901),
            .I(\c0.data_in_field_79 ));
    InMux I__3917 (
            .O(N__20892),
            .I(N__20888));
    InMux I__3916 (
            .O(N__20891),
            .I(N__20885));
    LocalMux I__3915 (
            .O(N__20888),
            .I(N__20882));
    LocalMux I__3914 (
            .O(N__20885),
            .I(N__20879));
    Odrv12 I__3913 (
            .O(N__20882),
            .I(\c0.n5545 ));
    Odrv4 I__3912 (
            .O(N__20879),
            .I(\c0.n5545 ));
    InMux I__3911 (
            .O(N__20874),
            .I(N__20871));
    LocalMux I__3910 (
            .O(N__20871),
            .I(N__20868));
    Span4Mux_h I__3909 (
            .O(N__20868),
            .I(N__20865));
    Span4Mux_h I__3908 (
            .O(N__20865),
            .I(N__20862));
    Odrv4 I__3907 (
            .O(N__20862),
            .I(\c0.n46 ));
    CascadeMux I__3906 (
            .O(N__20859),
            .I(N__20854));
    InMux I__3905 (
            .O(N__20858),
            .I(N__20851));
    InMux I__3904 (
            .O(N__20857),
            .I(N__20848));
    InMux I__3903 (
            .O(N__20854),
            .I(N__20844));
    LocalMux I__3902 (
            .O(N__20851),
            .I(N__20839));
    LocalMux I__3901 (
            .O(N__20848),
            .I(N__20836));
    InMux I__3900 (
            .O(N__20847),
            .I(N__20833));
    LocalMux I__3899 (
            .O(N__20844),
            .I(N__20830));
    InMux I__3898 (
            .O(N__20843),
            .I(N__20825));
    InMux I__3897 (
            .O(N__20842),
            .I(N__20825));
    Span4Mux_h I__3896 (
            .O(N__20839),
            .I(N__20818));
    Span4Mux_v I__3895 (
            .O(N__20836),
            .I(N__20818));
    LocalMux I__3894 (
            .O(N__20833),
            .I(N__20818));
    Odrv12 I__3893 (
            .O(N__20830),
            .I(\c0.data_in_field_95 ));
    LocalMux I__3892 (
            .O(N__20825),
            .I(\c0.data_in_field_95 ));
    Odrv4 I__3891 (
            .O(N__20818),
            .I(\c0.data_in_field_95 ));
    InMux I__3890 (
            .O(N__20811),
            .I(N__20806));
    InMux I__3889 (
            .O(N__20810),
            .I(N__20803));
    InMux I__3888 (
            .O(N__20809),
            .I(N__20799));
    LocalMux I__3887 (
            .O(N__20806),
            .I(N__20796));
    LocalMux I__3886 (
            .O(N__20803),
            .I(N__20793));
    CascadeMux I__3885 (
            .O(N__20802),
            .I(N__20790));
    LocalMux I__3884 (
            .O(N__20799),
            .I(N__20787));
    Span4Mux_s3_h I__3883 (
            .O(N__20796),
            .I(N__20784));
    Span4Mux_h I__3882 (
            .O(N__20793),
            .I(N__20781));
    InMux I__3881 (
            .O(N__20790),
            .I(N__20777));
    Span4Mux_v I__3880 (
            .O(N__20787),
            .I(N__20770));
    Span4Mux_v I__3879 (
            .O(N__20784),
            .I(N__20770));
    Span4Mux_v I__3878 (
            .O(N__20781),
            .I(N__20770));
    InMux I__3877 (
            .O(N__20780),
            .I(N__20767));
    LocalMux I__3876 (
            .O(N__20777),
            .I(\c0.data_in_field_96 ));
    Odrv4 I__3875 (
            .O(N__20770),
            .I(\c0.data_in_field_96 ));
    LocalMux I__3874 (
            .O(N__20767),
            .I(\c0.data_in_field_96 ));
    InMux I__3873 (
            .O(N__20760),
            .I(N__20757));
    LocalMux I__3872 (
            .O(N__20757),
            .I(\c0.n5590 ));
    CascadeMux I__3871 (
            .O(N__20754),
            .I(\c0.n40_cascade_ ));
    InMux I__3870 (
            .O(N__20751),
            .I(N__20748));
    LocalMux I__3869 (
            .O(N__20748),
            .I(N__20745));
    Odrv4 I__3868 (
            .O(N__20745),
            .I(\c0.n45_adj_1892 ));
    InMux I__3867 (
            .O(N__20742),
            .I(N__20736));
    InMux I__3866 (
            .O(N__20741),
            .I(N__20733));
    InMux I__3865 (
            .O(N__20740),
            .I(N__20730));
    InMux I__3864 (
            .O(N__20739),
            .I(N__20727));
    LocalMux I__3863 (
            .O(N__20736),
            .I(N__20724));
    LocalMux I__3862 (
            .O(N__20733),
            .I(N__20721));
    LocalMux I__3861 (
            .O(N__20730),
            .I(N__20718));
    LocalMux I__3860 (
            .O(N__20727),
            .I(N__20715));
    Span12Mux_v I__3859 (
            .O(N__20724),
            .I(N__20710));
    Span12Mux_s8_h I__3858 (
            .O(N__20721),
            .I(N__20707));
    Span4Mux_h I__3857 (
            .O(N__20718),
            .I(N__20702));
    Span4Mux_v I__3856 (
            .O(N__20715),
            .I(N__20702));
    InMux I__3855 (
            .O(N__20714),
            .I(N__20697));
    InMux I__3854 (
            .O(N__20713),
            .I(N__20697));
    Odrv12 I__3853 (
            .O(N__20710),
            .I(\c0.data_in_field_132 ));
    Odrv12 I__3852 (
            .O(N__20707),
            .I(\c0.data_in_field_132 ));
    Odrv4 I__3851 (
            .O(N__20702),
            .I(\c0.data_in_field_132 ));
    LocalMux I__3850 (
            .O(N__20697),
            .I(\c0.data_in_field_132 ));
    InMux I__3849 (
            .O(N__20688),
            .I(N__20685));
    LocalMux I__3848 (
            .O(N__20685),
            .I(N__20682));
    Odrv4 I__3847 (
            .O(N__20682),
            .I(\c0.n1969 ));
    InMux I__3846 (
            .O(N__20679),
            .I(N__20676));
    LocalMux I__3845 (
            .O(N__20676),
            .I(N__20672));
    InMux I__3844 (
            .O(N__20675),
            .I(N__20669));
    Span4Mux_h I__3843 (
            .O(N__20672),
            .I(N__20664));
    LocalMux I__3842 (
            .O(N__20669),
            .I(N__20664));
    Odrv4 I__3841 (
            .O(N__20664),
            .I(\c0.n5403 ));
    InMux I__3840 (
            .O(N__20661),
            .I(N__20658));
    LocalMux I__3839 (
            .O(N__20658),
            .I(N__20654));
    InMux I__3838 (
            .O(N__20657),
            .I(N__20650));
    Span4Mux_h I__3837 (
            .O(N__20654),
            .I(N__20647));
    InMux I__3836 (
            .O(N__20653),
            .I(N__20643));
    LocalMux I__3835 (
            .O(N__20650),
            .I(N__20640));
    Span4Mux_v I__3834 (
            .O(N__20647),
            .I(N__20637));
    InMux I__3833 (
            .O(N__20646),
            .I(N__20634));
    LocalMux I__3832 (
            .O(N__20643),
            .I(N__20631));
    Span4Mux_h I__3831 (
            .O(N__20640),
            .I(N__20626));
    Span4Mux_h I__3830 (
            .O(N__20637),
            .I(N__20626));
    LocalMux I__3829 (
            .O(N__20634),
            .I(data_in_19_4));
    Odrv4 I__3828 (
            .O(N__20631),
            .I(data_in_19_4));
    Odrv4 I__3827 (
            .O(N__20626),
            .I(data_in_19_4));
    InMux I__3826 (
            .O(N__20619),
            .I(N__20616));
    LocalMux I__3825 (
            .O(N__20616),
            .I(N__20610));
    InMux I__3824 (
            .O(N__20615),
            .I(N__20607));
    InMux I__3823 (
            .O(N__20614),
            .I(N__20604));
    InMux I__3822 (
            .O(N__20613),
            .I(N__20601));
    Span12Mux_s6_h I__3821 (
            .O(N__20610),
            .I(N__20598));
    LocalMux I__3820 (
            .O(N__20607),
            .I(N__20593));
    LocalMux I__3819 (
            .O(N__20604),
            .I(N__20593));
    LocalMux I__3818 (
            .O(N__20601),
            .I(\c0.data_in_field_115 ));
    Odrv12 I__3817 (
            .O(N__20598),
            .I(\c0.data_in_field_115 ));
    Odrv12 I__3816 (
            .O(N__20593),
            .I(\c0.data_in_field_115 ));
    CascadeMux I__3815 (
            .O(N__20586),
            .I(\c0.n1855_cascade_ ));
    InMux I__3814 (
            .O(N__20583),
            .I(N__20580));
    LocalMux I__3813 (
            .O(N__20580),
            .I(N__20577));
    Span4Mux_v I__3812 (
            .O(N__20577),
            .I(N__20573));
    InMux I__3811 (
            .O(N__20576),
            .I(N__20570));
    Span4Mux_h I__3810 (
            .O(N__20573),
            .I(N__20567));
    LocalMux I__3809 (
            .O(N__20570),
            .I(N__20564));
    Odrv4 I__3808 (
            .O(N__20567),
            .I(\c0.n1917 ));
    Odrv4 I__3807 (
            .O(N__20564),
            .I(\c0.n1917 ));
    InMux I__3806 (
            .O(N__20559),
            .I(N__20556));
    LocalMux I__3805 (
            .O(N__20556),
            .I(N__20552));
    InMux I__3804 (
            .O(N__20555),
            .I(N__20549));
    Span4Mux_h I__3803 (
            .O(N__20552),
            .I(N__20544));
    LocalMux I__3802 (
            .O(N__20549),
            .I(N__20544));
    Span4Mux_h I__3801 (
            .O(N__20544),
            .I(N__20538));
    InMux I__3800 (
            .O(N__20543),
            .I(N__20533));
    InMux I__3799 (
            .O(N__20542),
            .I(N__20533));
    InMux I__3798 (
            .O(N__20541),
            .I(N__20530));
    Odrv4 I__3797 (
            .O(N__20538),
            .I(\c0.data_in_field_34 ));
    LocalMux I__3796 (
            .O(N__20533),
            .I(\c0.data_in_field_34 ));
    LocalMux I__3795 (
            .O(N__20530),
            .I(\c0.data_in_field_34 ));
    InMux I__3794 (
            .O(N__20523),
            .I(N__20520));
    LocalMux I__3793 (
            .O(N__20520),
            .I(N__20517));
    Span4Mux_v I__3792 (
            .O(N__20517),
            .I(N__20513));
    InMux I__3791 (
            .O(N__20516),
            .I(N__20510));
    Span4Mux_h I__3790 (
            .O(N__20513),
            .I(N__20507));
    LocalMux I__3789 (
            .O(N__20510),
            .I(N__20504));
    Odrv4 I__3788 (
            .O(N__20507),
            .I(\c0.n2092 ));
    Odrv4 I__3787 (
            .O(N__20504),
            .I(\c0.n2092 ));
    InMux I__3786 (
            .O(N__20499),
            .I(N__20496));
    LocalMux I__3785 (
            .O(N__20496),
            .I(N__20492));
    InMux I__3784 (
            .O(N__20495),
            .I(N__20489));
    Span4Mux_v I__3783 (
            .O(N__20492),
            .I(N__20484));
    LocalMux I__3782 (
            .O(N__20489),
            .I(N__20484));
    Span4Mux_h I__3781 (
            .O(N__20484),
            .I(N__20481));
    Odrv4 I__3780 (
            .O(N__20481),
            .I(\c0.n5527 ));
    CascadeMux I__3779 (
            .O(N__20478),
            .I(\c0.n5394_cascade_ ));
    InMux I__3778 (
            .O(N__20475),
            .I(N__20472));
    LocalMux I__3777 (
            .O(N__20472),
            .I(N__20468));
    InMux I__3776 (
            .O(N__20471),
            .I(N__20465));
    Span4Mux_v I__3775 (
            .O(N__20468),
            .I(N__20462));
    LocalMux I__3774 (
            .O(N__20465),
            .I(N__20459));
    Span4Mux_h I__3773 (
            .O(N__20462),
            .I(N__20456));
    Span4Mux_h I__3772 (
            .O(N__20459),
            .I(N__20453));
    Odrv4 I__3771 (
            .O(N__20456),
            .I(\c0.n1926 ));
    Odrv4 I__3770 (
            .O(N__20453),
            .I(\c0.n1926 ));
    InMux I__3769 (
            .O(N__20448),
            .I(N__20445));
    LocalMux I__3768 (
            .O(N__20445),
            .I(N__20442));
    Span4Mux_v I__3767 (
            .O(N__20442),
            .I(N__20439));
    Span4Mux_v I__3766 (
            .O(N__20439),
            .I(N__20436));
    Span4Mux_h I__3765 (
            .O(N__20436),
            .I(N__20433));
    Odrv4 I__3764 (
            .O(N__20433),
            .I(\c0.n19_adj_1889 ));
    CascadeMux I__3763 (
            .O(N__20430),
            .I(N__20427));
    InMux I__3762 (
            .O(N__20427),
            .I(N__20424));
    LocalMux I__3761 (
            .O(N__20424),
            .I(N__20421));
    Odrv12 I__3760 (
            .O(N__20421),
            .I(\c0.n22_adj_1886 ));
    InMux I__3759 (
            .O(N__20418),
            .I(N__20413));
    InMux I__3758 (
            .O(N__20417),
            .I(N__20408));
    InMux I__3757 (
            .O(N__20416),
            .I(N__20405));
    LocalMux I__3756 (
            .O(N__20413),
            .I(N__20399));
    InMux I__3755 (
            .O(N__20412),
            .I(N__20396));
    InMux I__3754 (
            .O(N__20411),
            .I(N__20393));
    LocalMux I__3753 (
            .O(N__20408),
            .I(N__20388));
    LocalMux I__3752 (
            .O(N__20405),
            .I(N__20388));
    InMux I__3751 (
            .O(N__20404),
            .I(N__20385));
    InMux I__3750 (
            .O(N__20403),
            .I(N__20382));
    InMux I__3749 (
            .O(N__20402),
            .I(N__20379));
    Odrv4 I__3748 (
            .O(N__20399),
            .I(r_Bit_Index_0));
    LocalMux I__3747 (
            .O(N__20396),
            .I(r_Bit_Index_0));
    LocalMux I__3746 (
            .O(N__20393),
            .I(r_Bit_Index_0));
    Odrv4 I__3745 (
            .O(N__20388),
            .I(r_Bit_Index_0));
    LocalMux I__3744 (
            .O(N__20385),
            .I(r_Bit_Index_0));
    LocalMux I__3743 (
            .O(N__20382),
            .I(r_Bit_Index_0));
    LocalMux I__3742 (
            .O(N__20379),
            .I(r_Bit_Index_0));
    InMux I__3741 (
            .O(N__20364),
            .I(N__20356));
    InMux I__3740 (
            .O(N__20363),
            .I(N__20353));
    InMux I__3739 (
            .O(N__20362),
            .I(N__20350));
    CascadeMux I__3738 (
            .O(N__20361),
            .I(N__20346));
    InMux I__3737 (
            .O(N__20360),
            .I(N__20341));
    CascadeMux I__3736 (
            .O(N__20359),
            .I(N__20338));
    LocalMux I__3735 (
            .O(N__20356),
            .I(N__20335));
    LocalMux I__3734 (
            .O(N__20353),
            .I(N__20330));
    LocalMux I__3733 (
            .O(N__20350),
            .I(N__20330));
    InMux I__3732 (
            .O(N__20349),
            .I(N__20327));
    InMux I__3731 (
            .O(N__20346),
            .I(N__20320));
    InMux I__3730 (
            .O(N__20345),
            .I(N__20320));
    InMux I__3729 (
            .O(N__20344),
            .I(N__20320));
    LocalMux I__3728 (
            .O(N__20341),
            .I(N__20317));
    InMux I__3727 (
            .O(N__20338),
            .I(N__20313));
    Span4Mux_v I__3726 (
            .O(N__20335),
            .I(N__20304));
    Span4Mux_v I__3725 (
            .O(N__20330),
            .I(N__20304));
    LocalMux I__3724 (
            .O(N__20327),
            .I(N__20304));
    LocalMux I__3723 (
            .O(N__20320),
            .I(N__20304));
    Span4Mux_h I__3722 (
            .O(N__20317),
            .I(N__20301));
    CascadeMux I__3721 (
            .O(N__20316),
            .I(N__20296));
    LocalMux I__3720 (
            .O(N__20313),
            .I(N__20293));
    Span4Mux_h I__3719 (
            .O(N__20304),
            .I(N__20290));
    Sp12to4 I__3718 (
            .O(N__20301),
            .I(N__20287));
    InMux I__3717 (
            .O(N__20300),
            .I(N__20284));
    InMux I__3716 (
            .O(N__20299),
            .I(N__20279));
    InMux I__3715 (
            .O(N__20296),
            .I(N__20279));
    Span4Mux_v I__3714 (
            .O(N__20293),
            .I(N__20276));
    Span4Mux_s2_h I__3713 (
            .O(N__20290),
            .I(N__20273));
    Span12Mux_v I__3712 (
            .O(N__20287),
            .I(N__20270));
    LocalMux I__3711 (
            .O(N__20284),
            .I(N__20265));
    LocalMux I__3710 (
            .O(N__20279),
            .I(N__20265));
    Odrv4 I__3709 (
            .O(N__20276),
            .I(r_Rx_Data));
    Odrv4 I__3708 (
            .O(N__20273),
            .I(r_Rx_Data));
    Odrv12 I__3707 (
            .O(N__20270),
            .I(r_Rx_Data));
    Odrv4 I__3706 (
            .O(N__20265),
            .I(r_Rx_Data));
    InMux I__3705 (
            .O(N__20256),
            .I(N__20253));
    LocalMux I__3704 (
            .O(N__20253),
            .I(n1757));
    InMux I__3703 (
            .O(N__20250),
            .I(N__20246));
    InMux I__3702 (
            .O(N__20249),
            .I(N__20243));
    LocalMux I__3701 (
            .O(N__20246),
            .I(N__20240));
    LocalMux I__3700 (
            .O(N__20243),
            .I(N__20237));
    Span4Mux_v I__3699 (
            .O(N__20240),
            .I(N__20230));
    Span4Mux_v I__3698 (
            .O(N__20237),
            .I(N__20230));
    InMux I__3697 (
            .O(N__20236),
            .I(N__20227));
    InMux I__3696 (
            .O(N__20235),
            .I(N__20224));
    Span4Mux_v I__3695 (
            .O(N__20230),
            .I(N__20221));
    LocalMux I__3694 (
            .O(N__20227),
            .I(N__20218));
    LocalMux I__3693 (
            .O(N__20224),
            .I(data_in_3_6));
    Odrv4 I__3692 (
            .O(N__20221),
            .I(data_in_3_6));
    Odrv12 I__3691 (
            .O(N__20218),
            .I(data_in_3_6));
    InMux I__3690 (
            .O(N__20211),
            .I(N__20208));
    LocalMux I__3689 (
            .O(N__20208),
            .I(N__20205));
    Span4Mux_v I__3688 (
            .O(N__20205),
            .I(N__20202));
    Span4Mux_h I__3687 (
            .O(N__20202),
            .I(N__20197));
    InMux I__3686 (
            .O(N__20201),
            .I(N__20194));
    InMux I__3685 (
            .O(N__20200),
            .I(N__20191));
    Odrv4 I__3684 (
            .O(N__20197),
            .I(data_in_0_5));
    LocalMux I__3683 (
            .O(N__20194),
            .I(data_in_0_5));
    LocalMux I__3682 (
            .O(N__20191),
            .I(data_in_0_5));
    InMux I__3681 (
            .O(N__20184),
            .I(N__20181));
    LocalMux I__3680 (
            .O(N__20181),
            .I(N__20178));
    Odrv4 I__3679 (
            .O(N__20178),
            .I(\c0.n22_adj_1924 ));
    InMux I__3678 (
            .O(N__20175),
            .I(N__20172));
    LocalMux I__3677 (
            .O(N__20172),
            .I(N__20168));
    InMux I__3676 (
            .O(N__20171),
            .I(N__20165));
    Span4Mux_v I__3675 (
            .O(N__20168),
            .I(N__20160));
    LocalMux I__3674 (
            .O(N__20165),
            .I(N__20157));
    InMux I__3673 (
            .O(N__20164),
            .I(N__20154));
    InMux I__3672 (
            .O(N__20163),
            .I(N__20151));
    Span4Mux_h I__3671 (
            .O(N__20160),
            .I(N__20147));
    Span4Mux_v I__3670 (
            .O(N__20157),
            .I(N__20142));
    LocalMux I__3669 (
            .O(N__20154),
            .I(N__20142));
    LocalMux I__3668 (
            .O(N__20151),
            .I(N__20139));
    InMux I__3667 (
            .O(N__20150),
            .I(N__20136));
    Span4Mux_v I__3666 (
            .O(N__20147),
            .I(N__20129));
    Span4Mux_h I__3665 (
            .O(N__20142),
            .I(N__20129));
    Span4Mux_v I__3664 (
            .O(N__20139),
            .I(N__20129));
    LocalMux I__3663 (
            .O(N__20136),
            .I(\c0.data_in_field_141 ));
    Odrv4 I__3662 (
            .O(N__20129),
            .I(\c0.data_in_field_141 ));
    CascadeMux I__3661 (
            .O(N__20124),
            .I(N__20119));
    InMux I__3660 (
            .O(N__20123),
            .I(N__20113));
    InMux I__3659 (
            .O(N__20122),
            .I(N__20113));
    InMux I__3658 (
            .O(N__20119),
            .I(N__20110));
    InMux I__3657 (
            .O(N__20118),
            .I(N__20107));
    LocalMux I__3656 (
            .O(N__20113),
            .I(N__20102));
    LocalMux I__3655 (
            .O(N__20110),
            .I(N__20102));
    LocalMux I__3654 (
            .O(N__20107),
            .I(data_in_18_4));
    Odrv4 I__3653 (
            .O(N__20102),
            .I(data_in_18_4));
    CascadeMux I__3652 (
            .O(N__20097),
            .I(\c0.tx.n40_cascade_ ));
    InMux I__3651 (
            .O(N__20094),
            .I(N__20089));
    InMux I__3650 (
            .O(N__20093),
            .I(N__20084));
    InMux I__3649 (
            .O(N__20092),
            .I(N__20084));
    LocalMux I__3648 (
            .O(N__20089),
            .I(N__20081));
    LocalMux I__3647 (
            .O(N__20084),
            .I(N__20078));
    Odrv12 I__3646 (
            .O(N__20081),
            .I(n1760));
    Odrv4 I__3645 (
            .O(N__20078),
            .I(n1760));
    CEMux I__3644 (
            .O(N__20073),
            .I(N__20070));
    LocalMux I__3643 (
            .O(N__20070),
            .I(N__20067));
    Span4Mux_h I__3642 (
            .O(N__20067),
            .I(N__20063));
    InMux I__3641 (
            .O(N__20066),
            .I(N__20060));
    Odrv4 I__3640 (
            .O(N__20063),
            .I(\c0.tx.n2247 ));
    LocalMux I__3639 (
            .O(N__20060),
            .I(\c0.tx.n2247 ));
    SRMux I__3638 (
            .O(N__20055),
            .I(N__20052));
    LocalMux I__3637 (
            .O(N__20052),
            .I(\c0.tx.n2356 ));
    InMux I__3636 (
            .O(N__20049),
            .I(N__20046));
    LocalMux I__3635 (
            .O(N__20046),
            .I(N__20040));
    InMux I__3634 (
            .O(N__20045),
            .I(N__20037));
    InMux I__3633 (
            .O(N__20044),
            .I(N__20034));
    InMux I__3632 (
            .O(N__20043),
            .I(N__20029));
    Span4Mux_h I__3631 (
            .O(N__20040),
            .I(N__20026));
    LocalMux I__3630 (
            .O(N__20037),
            .I(N__20023));
    LocalMux I__3629 (
            .O(N__20034),
            .I(N__20020));
    InMux I__3628 (
            .O(N__20033),
            .I(N__20015));
    InMux I__3627 (
            .O(N__20032),
            .I(N__20015));
    LocalMux I__3626 (
            .O(N__20029),
            .I(\c0.rx.r_Bit_Index_2 ));
    Odrv4 I__3625 (
            .O(N__20026),
            .I(\c0.rx.r_Bit_Index_2 ));
    Odrv4 I__3624 (
            .O(N__20023),
            .I(\c0.rx.r_Bit_Index_2 ));
    Odrv4 I__3623 (
            .O(N__20020),
            .I(\c0.rx.r_Bit_Index_2 ));
    LocalMux I__3622 (
            .O(N__20015),
            .I(\c0.rx.r_Bit_Index_2 ));
    InMux I__3621 (
            .O(N__20004),
            .I(N__20001));
    LocalMux I__3620 (
            .O(N__20001),
            .I(N__19994));
    InMux I__3619 (
            .O(N__20000),
            .I(N__19991));
    InMux I__3618 (
            .O(N__19999),
            .I(N__19986));
    InMux I__3617 (
            .O(N__19998),
            .I(N__19983));
    InMux I__3616 (
            .O(N__19997),
            .I(N__19980));
    Span4Mux_h I__3615 (
            .O(N__19994),
            .I(N__19977));
    LocalMux I__3614 (
            .O(N__19991),
            .I(N__19974));
    InMux I__3613 (
            .O(N__19990),
            .I(N__19969));
    InMux I__3612 (
            .O(N__19989),
            .I(N__19969));
    LocalMux I__3611 (
            .O(N__19986),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__3610 (
            .O(N__19983),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__3609 (
            .O(N__19980),
            .I(\c0.rx.r_Bit_Index_1 ));
    Odrv4 I__3608 (
            .O(N__19977),
            .I(\c0.rx.r_Bit_Index_1 ));
    Odrv4 I__3607 (
            .O(N__19974),
            .I(\c0.rx.r_Bit_Index_1 ));
    LocalMux I__3606 (
            .O(N__19969),
            .I(\c0.rx.r_Bit_Index_1 ));
    InMux I__3605 (
            .O(N__19956),
            .I(N__19953));
    LocalMux I__3604 (
            .O(N__19953),
            .I(N__19948));
    InMux I__3603 (
            .O(N__19952),
            .I(N__19945));
    InMux I__3602 (
            .O(N__19951),
            .I(N__19942));
    Span4Mux_h I__3601 (
            .O(N__19948),
            .I(N__19939));
    LocalMux I__3600 (
            .O(N__19945),
            .I(N__19936));
    LocalMux I__3599 (
            .O(N__19942),
            .I(N__19933));
    Odrv4 I__3598 (
            .O(N__19939),
            .I(\c0.rx.n1706 ));
    Odrv4 I__3597 (
            .O(N__19936),
            .I(\c0.rx.n1706 ));
    Odrv4 I__3596 (
            .O(N__19933),
            .I(\c0.rx.n1706 ));
    CascadeMux I__3595 (
            .O(N__19926),
            .I(n1757_cascade_));
    InMux I__3594 (
            .O(N__19923),
            .I(N__19920));
    LocalMux I__3593 (
            .O(N__19920),
            .I(N__19917));
    Span4Mux_v I__3592 (
            .O(N__19917),
            .I(N__19913));
    InMux I__3591 (
            .O(N__19916),
            .I(N__19910));
    Odrv4 I__3590 (
            .O(N__19913),
            .I(rx_data_0));
    LocalMux I__3589 (
            .O(N__19910),
            .I(rx_data_0));
    CascadeMux I__3588 (
            .O(N__19905),
            .I(N__19902));
    InMux I__3587 (
            .O(N__19902),
            .I(N__19899));
    LocalMux I__3586 (
            .O(N__19899),
            .I(N__19894));
    InMux I__3585 (
            .O(N__19898),
            .I(N__19889));
    InMux I__3584 (
            .O(N__19897),
            .I(N__19889));
    Odrv4 I__3583 (
            .O(N__19894),
            .I(data_in_12_1));
    LocalMux I__3582 (
            .O(N__19889),
            .I(data_in_12_1));
    InMux I__3581 (
            .O(N__19884),
            .I(N__19881));
    LocalMux I__3580 (
            .O(N__19881),
            .I(N__19876));
    InMux I__3579 (
            .O(N__19880),
            .I(N__19873));
    InMux I__3578 (
            .O(N__19879),
            .I(N__19870));
    Span4Mux_v I__3577 (
            .O(N__19876),
            .I(N__19864));
    LocalMux I__3576 (
            .O(N__19873),
            .I(N__19864));
    LocalMux I__3575 (
            .O(N__19870),
            .I(N__19861));
    InMux I__3574 (
            .O(N__19869),
            .I(N__19857));
    Span4Mux_h I__3573 (
            .O(N__19864),
            .I(N__19854));
    Span4Mux_h I__3572 (
            .O(N__19861),
            .I(N__19851));
    InMux I__3571 (
            .O(N__19860),
            .I(N__19848));
    LocalMux I__3570 (
            .O(N__19857),
            .I(\c0.data_in_field_97 ));
    Odrv4 I__3569 (
            .O(N__19854),
            .I(\c0.data_in_field_97 ));
    Odrv4 I__3568 (
            .O(N__19851),
            .I(\c0.data_in_field_97 ));
    LocalMux I__3567 (
            .O(N__19848),
            .I(\c0.data_in_field_97 ));
    InMux I__3566 (
            .O(N__19839),
            .I(N__19836));
    LocalMux I__3565 (
            .O(N__19836),
            .I(N__19833));
    Span4Mux_v I__3564 (
            .O(N__19833),
            .I(N__19829));
    InMux I__3563 (
            .O(N__19832),
            .I(N__19826));
    Span4Mux_h I__3562 (
            .O(N__19829),
            .I(N__19823));
    LocalMux I__3561 (
            .O(N__19826),
            .I(\c0.data_in_frame_19_5 ));
    Odrv4 I__3560 (
            .O(N__19823),
            .I(\c0.data_in_frame_19_5 ));
    InMux I__3559 (
            .O(N__19818),
            .I(N__19815));
    LocalMux I__3558 (
            .O(N__19815),
            .I(N__19811));
    InMux I__3557 (
            .O(N__19814),
            .I(N__19808));
    Span4Mux_h I__3556 (
            .O(N__19811),
            .I(N__19804));
    LocalMux I__3555 (
            .O(N__19808),
            .I(N__19801));
    InMux I__3554 (
            .O(N__19807),
            .I(N__19798));
    Odrv4 I__3553 (
            .O(N__19804),
            .I(data_in_14_6));
    Odrv4 I__3552 (
            .O(N__19801),
            .I(data_in_14_6));
    LocalMux I__3551 (
            .O(N__19798),
            .I(data_in_14_6));
    InMux I__3550 (
            .O(N__19791),
            .I(N__19786));
    CascadeMux I__3549 (
            .O(N__19790),
            .I(N__19783));
    InMux I__3548 (
            .O(N__19789),
            .I(N__19779));
    LocalMux I__3547 (
            .O(N__19786),
            .I(N__19776));
    InMux I__3546 (
            .O(N__19783),
            .I(N__19773));
    InMux I__3545 (
            .O(N__19782),
            .I(N__19770));
    LocalMux I__3544 (
            .O(N__19779),
            .I(N__19767));
    Span4Mux_v I__3543 (
            .O(N__19776),
            .I(N__19764));
    LocalMux I__3542 (
            .O(N__19773),
            .I(N__19761));
    LocalMux I__3541 (
            .O(N__19770),
            .I(data_in_19_7));
    Odrv4 I__3540 (
            .O(N__19767),
            .I(data_in_19_7));
    Odrv4 I__3539 (
            .O(N__19764),
            .I(data_in_19_7));
    Odrv12 I__3538 (
            .O(N__19761),
            .I(data_in_19_7));
    CascadeMux I__3537 (
            .O(N__19752),
            .I(N__19749));
    InMux I__3536 (
            .O(N__19749),
            .I(N__19746));
    LocalMux I__3535 (
            .O(N__19746),
            .I(N__19742));
    InMux I__3534 (
            .O(N__19745),
            .I(N__19739));
    Span4Mux_s3_h I__3533 (
            .O(N__19742),
            .I(N__19736));
    LocalMux I__3532 (
            .O(N__19739),
            .I(\c0.data_in_frame_19_7 ));
    Odrv4 I__3531 (
            .O(N__19736),
            .I(\c0.data_in_frame_19_7 ));
    CascadeMux I__3530 (
            .O(N__19731),
            .I(N__19726));
    InMux I__3529 (
            .O(N__19730),
            .I(N__19721));
    InMux I__3528 (
            .O(N__19729),
            .I(N__19721));
    InMux I__3527 (
            .O(N__19726),
            .I(N__19718));
    LocalMux I__3526 (
            .O(N__19721),
            .I(N__19715));
    LocalMux I__3525 (
            .O(N__19718),
            .I(N__19711));
    Span4Mux_h I__3524 (
            .O(N__19715),
            .I(N__19708));
    InMux I__3523 (
            .O(N__19714),
            .I(N__19705));
    Span4Mux_v I__3522 (
            .O(N__19711),
            .I(N__19702));
    Odrv4 I__3521 (
            .O(N__19708),
            .I(data_in_19_5));
    LocalMux I__3520 (
            .O(N__19705),
            .I(data_in_19_5));
    Odrv4 I__3519 (
            .O(N__19702),
            .I(data_in_19_5));
    CascadeMux I__3518 (
            .O(N__19695),
            .I(N__19692));
    InMux I__3517 (
            .O(N__19692),
            .I(N__19689));
    LocalMux I__3516 (
            .O(N__19689),
            .I(N__19684));
    InMux I__3515 (
            .O(N__19688),
            .I(N__19681));
    InMux I__3514 (
            .O(N__19687),
            .I(N__19678));
    Odrv4 I__3513 (
            .O(N__19684),
            .I(data_in_14_0));
    LocalMux I__3512 (
            .O(N__19681),
            .I(data_in_14_0));
    LocalMux I__3511 (
            .O(N__19678),
            .I(data_in_14_0));
    InMux I__3510 (
            .O(N__19671),
            .I(N__19667));
    InMux I__3509 (
            .O(N__19670),
            .I(N__19664));
    LocalMux I__3508 (
            .O(N__19667),
            .I(N__19661));
    LocalMux I__3507 (
            .O(N__19664),
            .I(N__19658));
    Span12Mux_v I__3506 (
            .O(N__19661),
            .I(N__19654));
    Span4Mux_v I__3505 (
            .O(N__19658),
            .I(N__19651));
    InMux I__3504 (
            .O(N__19657),
            .I(N__19648));
    Odrv12 I__3503 (
            .O(N__19654),
            .I(data_in_13_0));
    Odrv4 I__3502 (
            .O(N__19651),
            .I(data_in_13_0));
    LocalMux I__3501 (
            .O(N__19648),
            .I(data_in_13_0));
    InMux I__3500 (
            .O(N__19641),
            .I(N__19636));
    InMux I__3499 (
            .O(N__19640),
            .I(N__19633));
    InMux I__3498 (
            .O(N__19639),
            .I(N__19630));
    LocalMux I__3497 (
            .O(N__19636),
            .I(N__19627));
    LocalMux I__3496 (
            .O(N__19633),
            .I(N__19624));
    LocalMux I__3495 (
            .O(N__19630),
            .I(N__19621));
    Span4Mux_s2_h I__3494 (
            .O(N__19627),
            .I(N__19618));
    Span12Mux_s6_h I__3493 (
            .O(N__19624),
            .I(N__19613));
    Span4Mux_v I__3492 (
            .O(N__19621),
            .I(N__19610));
    Span4Mux_h I__3491 (
            .O(N__19618),
            .I(N__19607));
    InMux I__3490 (
            .O(N__19617),
            .I(N__19602));
    InMux I__3489 (
            .O(N__19616),
            .I(N__19602));
    Odrv12 I__3488 (
            .O(N__19613),
            .I(\c0.data_in_field_36 ));
    Odrv4 I__3487 (
            .O(N__19610),
            .I(\c0.data_in_field_36 ));
    Odrv4 I__3486 (
            .O(N__19607),
            .I(\c0.data_in_field_36 ));
    LocalMux I__3485 (
            .O(N__19602),
            .I(\c0.data_in_field_36 ));
    InMux I__3484 (
            .O(N__19593),
            .I(N__19590));
    LocalMux I__3483 (
            .O(N__19590),
            .I(N__19586));
    InMux I__3482 (
            .O(N__19589),
            .I(N__19583));
    Span4Mux_s2_h I__3481 (
            .O(N__19586),
            .I(N__19579));
    LocalMux I__3480 (
            .O(N__19583),
            .I(N__19576));
    InMux I__3479 (
            .O(N__19582),
            .I(N__19572));
    Span4Mux_h I__3478 (
            .O(N__19579),
            .I(N__19567));
    Span4Mux_h I__3477 (
            .O(N__19576),
            .I(N__19567));
    InMux I__3476 (
            .O(N__19575),
            .I(N__19564));
    LocalMux I__3475 (
            .O(N__19572),
            .I(\c0.data_in_field_82 ));
    Odrv4 I__3474 (
            .O(N__19567),
            .I(\c0.data_in_field_82 ));
    LocalMux I__3473 (
            .O(N__19564),
            .I(\c0.data_in_field_82 ));
    InMux I__3472 (
            .O(N__19557),
            .I(N__19554));
    LocalMux I__3471 (
            .O(N__19554),
            .I(N__19550));
    InMux I__3470 (
            .O(N__19553),
            .I(N__19546));
    Span4Mux_v I__3469 (
            .O(N__19550),
            .I(N__19543));
    InMux I__3468 (
            .O(N__19549),
            .I(N__19540));
    LocalMux I__3467 (
            .O(N__19546),
            .I(\c0.n1948 ));
    Odrv4 I__3466 (
            .O(N__19543),
            .I(\c0.n1948 ));
    LocalMux I__3465 (
            .O(N__19540),
            .I(\c0.n1948 ));
    InMux I__3464 (
            .O(N__19533),
            .I(N__19530));
    LocalMux I__3463 (
            .O(N__19530),
            .I(N__19526));
    CascadeMux I__3462 (
            .O(N__19529),
            .I(N__19523));
    Span4Mux_v I__3461 (
            .O(N__19526),
            .I(N__19520));
    InMux I__3460 (
            .O(N__19523),
            .I(N__19516));
    Span4Mux_h I__3459 (
            .O(N__19520),
            .I(N__19513));
    InMux I__3458 (
            .O(N__19519),
            .I(N__19510));
    LocalMux I__3457 (
            .O(N__19516),
            .I(data_in_15_1));
    Odrv4 I__3456 (
            .O(N__19513),
            .I(data_in_15_1));
    LocalMux I__3455 (
            .O(N__19510),
            .I(data_in_15_1));
    CascadeMux I__3454 (
            .O(N__19503),
            .I(N__19500));
    InMux I__3453 (
            .O(N__19500),
            .I(N__19496));
    InMux I__3452 (
            .O(N__19499),
            .I(N__19493));
    LocalMux I__3451 (
            .O(N__19496),
            .I(N__19490));
    LocalMux I__3450 (
            .O(N__19493),
            .I(N__19487));
    Span4Mux_h I__3449 (
            .O(N__19490),
            .I(N__19481));
    Span4Mux_v I__3448 (
            .O(N__19487),
            .I(N__19481));
    InMux I__3447 (
            .O(N__19486),
            .I(N__19478));
    Odrv4 I__3446 (
            .O(N__19481),
            .I(data_in_14_1));
    LocalMux I__3445 (
            .O(N__19478),
            .I(data_in_14_1));
    InMux I__3444 (
            .O(N__19473),
            .I(N__19470));
    LocalMux I__3443 (
            .O(N__19470),
            .I(N__19465));
    CascadeMux I__3442 (
            .O(N__19469),
            .I(N__19462));
    InMux I__3441 (
            .O(N__19468),
            .I(N__19458));
    Span4Mux_v I__3440 (
            .O(N__19465),
            .I(N__19455));
    InMux I__3439 (
            .O(N__19462),
            .I(N__19450));
    InMux I__3438 (
            .O(N__19461),
            .I(N__19450));
    LocalMux I__3437 (
            .O(N__19458),
            .I(\c0.data_in_field_127 ));
    Odrv4 I__3436 (
            .O(N__19455),
            .I(\c0.data_in_field_127 ));
    LocalMux I__3435 (
            .O(N__19450),
            .I(\c0.data_in_field_127 ));
    InMux I__3434 (
            .O(N__19443),
            .I(N__19440));
    LocalMux I__3433 (
            .O(N__19440),
            .I(N__19436));
    InMux I__3432 (
            .O(N__19439),
            .I(N__19433));
    Sp12to4 I__3431 (
            .O(N__19436),
            .I(N__19430));
    LocalMux I__3430 (
            .O(N__19433),
            .I(N__19427));
    Span12Mux_v I__3429 (
            .O(N__19430),
            .I(N__19424));
    Span4Mux_v I__3428 (
            .O(N__19427),
            .I(N__19421));
    Odrv12 I__3427 (
            .O(N__19424),
            .I(n4));
    Odrv4 I__3426 (
            .O(N__19421),
            .I(n4));
    CascadeMux I__3425 (
            .O(N__19416),
            .I(N__19413));
    InMux I__3424 (
            .O(N__19413),
            .I(N__19410));
    LocalMux I__3423 (
            .O(N__19410),
            .I(N__19407));
    Span4Mux_h I__3422 (
            .O(N__19407),
            .I(N__19402));
    InMux I__3421 (
            .O(N__19406),
            .I(N__19397));
    InMux I__3420 (
            .O(N__19405),
            .I(N__19397));
    Odrv4 I__3419 (
            .O(N__19402),
            .I(data_in_13_1));
    LocalMux I__3418 (
            .O(N__19397),
            .I(data_in_13_1));
    InMux I__3417 (
            .O(N__19392),
            .I(N__19389));
    LocalMux I__3416 (
            .O(N__19389),
            .I(N__19385));
    InMux I__3415 (
            .O(N__19388),
            .I(N__19382));
    Span4Mux_v I__3414 (
            .O(N__19385),
            .I(N__19377));
    LocalMux I__3413 (
            .O(N__19382),
            .I(N__19377));
    Span4Mux_h I__3412 (
            .O(N__19377),
            .I(N__19373));
    InMux I__3411 (
            .O(N__19376),
            .I(N__19370));
    Span4Mux_v I__3410 (
            .O(N__19373),
            .I(N__19367));
    LocalMux I__3409 (
            .O(N__19370),
            .I(\c0.data_in_field_105 ));
    Odrv4 I__3408 (
            .O(N__19367),
            .I(\c0.data_in_field_105 ));
    InMux I__3407 (
            .O(N__19362),
            .I(N__19359));
    LocalMux I__3406 (
            .O(N__19359),
            .I(\c0.n18_adj_1887 ));
    InMux I__3405 (
            .O(N__19356),
            .I(N__19353));
    LocalMux I__3404 (
            .O(N__19353),
            .I(N__19350));
    Span4Mux_s3_h I__3403 (
            .O(N__19350),
            .I(N__19347));
    Span4Mux_h I__3402 (
            .O(N__19347),
            .I(N__19344));
    Odrv4 I__3401 (
            .O(N__19344),
            .I(\c0.n20_adj_1888 ));
    CascadeMux I__3400 (
            .O(N__19341),
            .I(\c0.tx2_transmit_N_1031_cascade_ ));
    InMux I__3399 (
            .O(N__19338),
            .I(N__19333));
    InMux I__3398 (
            .O(N__19337),
            .I(N__19328));
    InMux I__3397 (
            .O(N__19336),
            .I(N__19328));
    LocalMux I__3396 (
            .O(N__19333),
            .I(\c0.data_in_field_29 ));
    LocalMux I__3395 (
            .O(N__19328),
            .I(\c0.data_in_field_29 ));
    InMux I__3394 (
            .O(N__19323),
            .I(N__19320));
    LocalMux I__3393 (
            .O(N__19320),
            .I(N__19317));
    Odrv12 I__3392 (
            .O(N__19317),
            .I(\c0.n2030 ));
    CascadeMux I__3391 (
            .O(N__19314),
            .I(\c0.n2030_cascade_ ));
    InMux I__3390 (
            .O(N__19311),
            .I(N__19308));
    LocalMux I__3389 (
            .O(N__19308),
            .I(N__19305));
    Span4Mux_v I__3388 (
            .O(N__19305),
            .I(N__19302));
    Span4Mux_h I__3387 (
            .O(N__19302),
            .I(N__19298));
    InMux I__3386 (
            .O(N__19301),
            .I(N__19295));
    Span4Mux_h I__3385 (
            .O(N__19298),
            .I(N__19289));
    LocalMux I__3384 (
            .O(N__19295),
            .I(N__19289));
    InMux I__3383 (
            .O(N__19294),
            .I(N__19286));
    Odrv4 I__3382 (
            .O(N__19289),
            .I(data_in_15_2));
    LocalMux I__3381 (
            .O(N__19286),
            .I(data_in_15_2));
    InMux I__3380 (
            .O(N__19281),
            .I(N__19278));
    LocalMux I__3379 (
            .O(N__19278),
            .I(N__19275));
    Span4Mux_h I__3378 (
            .O(N__19275),
            .I(N__19270));
    InMux I__3377 (
            .O(N__19274),
            .I(N__19265));
    InMux I__3376 (
            .O(N__19273),
            .I(N__19265));
    Odrv4 I__3375 (
            .O(N__19270),
            .I(\c0.data_in_field_22 ));
    LocalMux I__3374 (
            .O(N__19265),
            .I(\c0.data_in_field_22 ));
    InMux I__3373 (
            .O(N__19260),
            .I(N__19257));
    LocalMux I__3372 (
            .O(N__19257),
            .I(N__19254));
    Span4Mux_v I__3371 (
            .O(N__19254),
            .I(N__19251));
    Odrv4 I__3370 (
            .O(N__19251),
            .I(\c0.n5436 ));
    CascadeMux I__3369 (
            .O(N__19248),
            .I(\c0.n5436_cascade_ ));
    InMux I__3368 (
            .O(N__19245),
            .I(N__19242));
    LocalMux I__3367 (
            .O(N__19242),
            .I(\c0.n5509 ));
    InMux I__3366 (
            .O(N__19239),
            .I(N__19236));
    LocalMux I__3365 (
            .O(N__19236),
            .I(N__19229));
    InMux I__3364 (
            .O(N__19235),
            .I(N__19226));
    InMux I__3363 (
            .O(N__19234),
            .I(N__19219));
    InMux I__3362 (
            .O(N__19233),
            .I(N__19219));
    InMux I__3361 (
            .O(N__19232),
            .I(N__19219));
    Odrv4 I__3360 (
            .O(N__19229),
            .I(\c0.data_in_field_78 ));
    LocalMux I__3359 (
            .O(N__19226),
            .I(\c0.data_in_field_78 ));
    LocalMux I__3358 (
            .O(N__19219),
            .I(\c0.data_in_field_78 ));
    CascadeMux I__3357 (
            .O(N__19212),
            .I(\c0.n5509_cascade_ ));
    CascadeMux I__3356 (
            .O(N__19209),
            .I(N__19203));
    InMux I__3355 (
            .O(N__19208),
            .I(N__19200));
    InMux I__3354 (
            .O(N__19207),
            .I(N__19197));
    InMux I__3353 (
            .O(N__19206),
            .I(N__19192));
    InMux I__3352 (
            .O(N__19203),
            .I(N__19192));
    LocalMux I__3351 (
            .O(N__19200),
            .I(N__19185));
    LocalMux I__3350 (
            .O(N__19197),
            .I(N__19185));
    LocalMux I__3349 (
            .O(N__19192),
            .I(N__19182));
    InMux I__3348 (
            .O(N__19191),
            .I(N__19179));
    InMux I__3347 (
            .O(N__19190),
            .I(N__19176));
    Span4Mux_v I__3346 (
            .O(N__19185),
            .I(N__19171));
    Span4Mux_h I__3345 (
            .O(N__19182),
            .I(N__19171));
    LocalMux I__3344 (
            .O(N__19179),
            .I(\c0.data_in_field_92 ));
    LocalMux I__3343 (
            .O(N__19176),
            .I(\c0.data_in_field_92 ));
    Odrv4 I__3342 (
            .O(N__19171),
            .I(\c0.data_in_field_92 ));
    CascadeMux I__3341 (
            .O(N__19164),
            .I(N__19160));
    InMux I__3340 (
            .O(N__19163),
            .I(N__19156));
    InMux I__3339 (
            .O(N__19160),
            .I(N__19153));
    InMux I__3338 (
            .O(N__19159),
            .I(N__19150));
    LocalMux I__3337 (
            .O(N__19156),
            .I(\c0.data_in_field_52 ));
    LocalMux I__3336 (
            .O(N__19153),
            .I(\c0.data_in_field_52 ));
    LocalMux I__3335 (
            .O(N__19150),
            .I(\c0.data_in_field_52 ));
    InMux I__3334 (
            .O(N__19143),
            .I(N__19140));
    LocalMux I__3333 (
            .O(N__19140),
            .I(N__19137));
    Span4Mux_h I__3332 (
            .O(N__19137),
            .I(N__19133));
    InMux I__3331 (
            .O(N__19136),
            .I(N__19129));
    Span4Mux_v I__3330 (
            .O(N__19133),
            .I(N__19126));
    InMux I__3329 (
            .O(N__19132),
            .I(N__19123));
    LocalMux I__3328 (
            .O(N__19129),
            .I(\c0.data_in_field_103 ));
    Odrv4 I__3327 (
            .O(N__19126),
            .I(\c0.data_in_field_103 ));
    LocalMux I__3326 (
            .O(N__19123),
            .I(\c0.data_in_field_103 ));
    InMux I__3325 (
            .O(N__19116),
            .I(N__19113));
    LocalMux I__3324 (
            .O(N__19113),
            .I(\c0.n2152 ));
    InMux I__3323 (
            .O(N__19110),
            .I(N__19107));
    LocalMux I__3322 (
            .O(N__19107),
            .I(N__19102));
    InMux I__3321 (
            .O(N__19106),
            .I(N__19098));
    InMux I__3320 (
            .O(N__19105),
            .I(N__19095));
    Span4Mux_v I__3319 (
            .O(N__19102),
            .I(N__19092));
    InMux I__3318 (
            .O(N__19101),
            .I(N__19089));
    LocalMux I__3317 (
            .O(N__19098),
            .I(N__19084));
    LocalMux I__3316 (
            .O(N__19095),
            .I(N__19084));
    Odrv4 I__3315 (
            .O(N__19092),
            .I(\c0.data_in_field_43 ));
    LocalMux I__3314 (
            .O(N__19089),
            .I(\c0.data_in_field_43 ));
    Odrv4 I__3313 (
            .O(N__19084),
            .I(\c0.data_in_field_43 ));
    CascadeMux I__3312 (
            .O(N__19077),
            .I(\c0.n2152_cascade_ ));
    InMux I__3311 (
            .O(N__19074),
            .I(N__19071));
    LocalMux I__3310 (
            .O(N__19071),
            .I(N__19067));
    InMux I__3309 (
            .O(N__19070),
            .I(N__19064));
    Span4Mux_h I__3308 (
            .O(N__19067),
            .I(N__19061));
    LocalMux I__3307 (
            .O(N__19064),
            .I(N__19058));
    Odrv4 I__3306 (
            .O(N__19061),
            .I(\c0.n5397 ));
    Odrv4 I__3305 (
            .O(N__19058),
            .I(\c0.n5397 ));
    CascadeMux I__3304 (
            .O(N__19053),
            .I(N__19050));
    InMux I__3303 (
            .O(N__19050),
            .I(N__19047));
    LocalMux I__3302 (
            .O(N__19047),
            .I(N__19044));
    Span4Mux_v I__3301 (
            .O(N__19044),
            .I(N__19039));
    InMux I__3300 (
            .O(N__19043),
            .I(N__19036));
    InMux I__3299 (
            .O(N__19042),
            .I(N__19033));
    Odrv4 I__3298 (
            .O(N__19039),
            .I(data_in_11_6));
    LocalMux I__3297 (
            .O(N__19036),
            .I(data_in_11_6));
    LocalMux I__3296 (
            .O(N__19033),
            .I(data_in_11_6));
    InMux I__3295 (
            .O(N__19026),
            .I(N__19023));
    LocalMux I__3294 (
            .O(N__19023),
            .I(N__19017));
    InMux I__3293 (
            .O(N__19022),
            .I(N__19014));
    CascadeMux I__3292 (
            .O(N__19021),
            .I(N__19011));
    InMux I__3291 (
            .O(N__19020),
            .I(N__19008));
    Span4Mux_v I__3290 (
            .O(N__19017),
            .I(N__19005));
    LocalMux I__3289 (
            .O(N__19014),
            .I(N__19002));
    InMux I__3288 (
            .O(N__19011),
            .I(N__18999));
    LocalMux I__3287 (
            .O(N__19008),
            .I(\c0.data_in_field_75 ));
    Odrv4 I__3286 (
            .O(N__19005),
            .I(\c0.data_in_field_75 ));
    Odrv4 I__3285 (
            .O(N__19002),
            .I(\c0.data_in_field_75 ));
    LocalMux I__3284 (
            .O(N__18999),
            .I(\c0.data_in_field_75 ));
    CascadeMux I__3283 (
            .O(N__18990),
            .I(N__18987));
    InMux I__3282 (
            .O(N__18987),
            .I(N__18984));
    LocalMux I__3281 (
            .O(N__18984),
            .I(N__18981));
    Sp12to4 I__3280 (
            .O(N__18981),
            .I(N__18978));
    Span12Mux_v I__3279 (
            .O(N__18978),
            .I(N__18973));
    InMux I__3278 (
            .O(N__18977),
            .I(N__18968));
    InMux I__3277 (
            .O(N__18976),
            .I(N__18968));
    Odrv12 I__3276 (
            .O(N__18973),
            .I(data_in_17_6));
    LocalMux I__3275 (
            .O(N__18968),
            .I(data_in_17_6));
    InMux I__3274 (
            .O(N__18963),
            .I(N__18959));
    CascadeMux I__3273 (
            .O(N__18962),
            .I(N__18955));
    LocalMux I__3272 (
            .O(N__18959),
            .I(N__18952));
    CascadeMux I__3271 (
            .O(N__18958),
            .I(N__18949));
    InMux I__3270 (
            .O(N__18955),
            .I(N__18946));
    Span4Mux_v I__3269 (
            .O(N__18952),
            .I(N__18941));
    InMux I__3268 (
            .O(N__18949),
            .I(N__18938));
    LocalMux I__3267 (
            .O(N__18946),
            .I(N__18935));
    InMux I__3266 (
            .O(N__18945),
            .I(N__18930));
    InMux I__3265 (
            .O(N__18944),
            .I(N__18930));
    Odrv4 I__3264 (
            .O(N__18941),
            .I(\c0.data_in_field_142 ));
    LocalMux I__3263 (
            .O(N__18938),
            .I(\c0.data_in_field_142 ));
    Odrv4 I__3262 (
            .O(N__18935),
            .I(\c0.data_in_field_142 ));
    LocalMux I__3261 (
            .O(N__18930),
            .I(\c0.data_in_field_142 ));
    CascadeMux I__3260 (
            .O(N__18921),
            .I(N__18918));
    InMux I__3259 (
            .O(N__18918),
            .I(N__18915));
    LocalMux I__3258 (
            .O(N__18915),
            .I(N__18911));
    InMux I__3257 (
            .O(N__18914),
            .I(N__18906));
    Span12Mux_s6_h I__3256 (
            .O(N__18911),
            .I(N__18903));
    InMux I__3255 (
            .O(N__18910),
            .I(N__18898));
    InMux I__3254 (
            .O(N__18909),
            .I(N__18898));
    LocalMux I__3253 (
            .O(N__18906),
            .I(N__18895));
    Odrv12 I__3252 (
            .O(N__18903),
            .I(\c0.data_in_field_33 ));
    LocalMux I__3251 (
            .O(N__18898),
            .I(\c0.data_in_field_33 ));
    Odrv4 I__3250 (
            .O(N__18895),
            .I(\c0.data_in_field_33 ));
    InMux I__3249 (
            .O(N__18888),
            .I(N__18885));
    LocalMux I__3248 (
            .O(N__18885),
            .I(N__18882));
    Span4Mux_h I__3247 (
            .O(N__18882),
            .I(N__18878));
    InMux I__3246 (
            .O(N__18881),
            .I(N__18873));
    Span4Mux_v I__3245 (
            .O(N__18878),
            .I(N__18870));
    InMux I__3244 (
            .O(N__18877),
            .I(N__18867));
    InMux I__3243 (
            .O(N__18876),
            .I(N__18864));
    LocalMux I__3242 (
            .O(N__18873),
            .I(\c0.data_in_field_140 ));
    Odrv4 I__3241 (
            .O(N__18870),
            .I(\c0.data_in_field_140 ));
    LocalMux I__3240 (
            .O(N__18867),
            .I(\c0.data_in_field_140 ));
    LocalMux I__3239 (
            .O(N__18864),
            .I(\c0.data_in_field_140 ));
    InMux I__3238 (
            .O(N__18855),
            .I(N__18851));
    InMux I__3237 (
            .O(N__18854),
            .I(N__18848));
    LocalMux I__3236 (
            .O(N__18851),
            .I(N__18845));
    LocalMux I__3235 (
            .O(N__18848),
            .I(N__18842));
    Span4Mux_h I__3234 (
            .O(N__18845),
            .I(N__18836));
    Span4Mux_v I__3233 (
            .O(N__18842),
            .I(N__18836));
    InMux I__3232 (
            .O(N__18841),
            .I(N__18833));
    Odrv4 I__3231 (
            .O(N__18836),
            .I(data_in_12_7));
    LocalMux I__3230 (
            .O(N__18833),
            .I(data_in_12_7));
    InMux I__3229 (
            .O(N__18828),
            .I(N__18825));
    LocalMux I__3228 (
            .O(N__18825),
            .I(N__18820));
    InMux I__3227 (
            .O(N__18824),
            .I(N__18817));
    InMux I__3226 (
            .O(N__18823),
            .I(N__18814));
    Span4Mux_v I__3225 (
            .O(N__18820),
            .I(N__18809));
    LocalMux I__3224 (
            .O(N__18817),
            .I(N__18804));
    LocalMux I__3223 (
            .O(N__18814),
            .I(N__18804));
    InMux I__3222 (
            .O(N__18813),
            .I(N__18799));
    InMux I__3221 (
            .O(N__18812),
            .I(N__18799));
    Odrv4 I__3220 (
            .O(N__18809),
            .I(\c0.data_in_field_126 ));
    Odrv4 I__3219 (
            .O(N__18804),
            .I(\c0.data_in_field_126 ));
    LocalMux I__3218 (
            .O(N__18799),
            .I(\c0.data_in_field_126 ));
    CascadeMux I__3217 (
            .O(N__18792),
            .I(N__18786));
    CascadeMux I__3216 (
            .O(N__18791),
            .I(N__18783));
    InMux I__3215 (
            .O(N__18790),
            .I(N__18780));
    InMux I__3214 (
            .O(N__18789),
            .I(N__18777));
    InMux I__3213 (
            .O(N__18786),
            .I(N__18774));
    InMux I__3212 (
            .O(N__18783),
            .I(N__18771));
    LocalMux I__3211 (
            .O(N__18780),
            .I(N__18768));
    LocalMux I__3210 (
            .O(N__18777),
            .I(N__18763));
    LocalMux I__3209 (
            .O(N__18774),
            .I(N__18763));
    LocalMux I__3208 (
            .O(N__18771),
            .I(N__18758));
    Span4Mux_h I__3207 (
            .O(N__18768),
            .I(N__18758));
    Span4Mux_h I__3206 (
            .O(N__18763),
            .I(N__18755));
    Odrv4 I__3205 (
            .O(N__18758),
            .I(\c0.data_in_field_118 ));
    Odrv4 I__3204 (
            .O(N__18755),
            .I(\c0.data_in_field_118 ));
    CascadeMux I__3203 (
            .O(N__18750),
            .I(N__18747));
    InMux I__3202 (
            .O(N__18747),
            .I(N__18744));
    LocalMux I__3201 (
            .O(N__18744),
            .I(N__18740));
    InMux I__3200 (
            .O(N__18743),
            .I(N__18737));
    Span4Mux_s2_h I__3199 (
            .O(N__18740),
            .I(N__18733));
    LocalMux I__3198 (
            .O(N__18737),
            .I(N__18730));
    InMux I__3197 (
            .O(N__18736),
            .I(N__18727));
    Span4Mux_h I__3196 (
            .O(N__18733),
            .I(N__18719));
    Span4Mux_h I__3195 (
            .O(N__18730),
            .I(N__18719));
    LocalMux I__3194 (
            .O(N__18727),
            .I(N__18719));
    InMux I__3193 (
            .O(N__18726),
            .I(N__18715));
    Span4Mux_v I__3192 (
            .O(N__18719),
            .I(N__18712));
    InMux I__3191 (
            .O(N__18718),
            .I(N__18709));
    LocalMux I__3190 (
            .O(N__18715),
            .I(\c0.data_in_field_51 ));
    Odrv4 I__3189 (
            .O(N__18712),
            .I(\c0.data_in_field_51 ));
    LocalMux I__3188 (
            .O(N__18709),
            .I(\c0.data_in_field_51 ));
    CascadeMux I__3187 (
            .O(N__18702),
            .I(N__18699));
    InMux I__3186 (
            .O(N__18699),
            .I(N__18696));
    LocalMux I__3185 (
            .O(N__18696),
            .I(N__18691));
    InMux I__3184 (
            .O(N__18695),
            .I(N__18686));
    InMux I__3183 (
            .O(N__18694),
            .I(N__18686));
    Odrv4 I__3182 (
            .O(N__18691),
            .I(data_in_16_5));
    LocalMux I__3181 (
            .O(N__18686),
            .I(data_in_16_5));
    CascadeMux I__3180 (
            .O(N__18681),
            .I(N__18678));
    InMux I__3179 (
            .O(N__18678),
            .I(N__18675));
    LocalMux I__3178 (
            .O(N__18675),
            .I(N__18672));
    Span4Mux_v I__3177 (
            .O(N__18672),
            .I(N__18667));
    InMux I__3176 (
            .O(N__18671),
            .I(N__18664));
    InMux I__3175 (
            .O(N__18670),
            .I(N__18661));
    Odrv4 I__3174 (
            .O(N__18667),
            .I(data_in_9_3));
    LocalMux I__3173 (
            .O(N__18664),
            .I(data_in_9_3));
    LocalMux I__3172 (
            .O(N__18661),
            .I(data_in_9_3));
    InMux I__3171 (
            .O(N__18654),
            .I(N__18650));
    InMux I__3170 (
            .O(N__18653),
            .I(N__18647));
    LocalMux I__3169 (
            .O(N__18650),
            .I(N__18641));
    LocalMux I__3168 (
            .O(N__18647),
            .I(N__18641));
    InMux I__3167 (
            .O(N__18646),
            .I(N__18637));
    Span4Mux_h I__3166 (
            .O(N__18641),
            .I(N__18634));
    InMux I__3165 (
            .O(N__18640),
            .I(N__18631));
    LocalMux I__3164 (
            .O(N__18637),
            .I(\c0.data_in_field_3 ));
    Odrv4 I__3163 (
            .O(N__18634),
            .I(\c0.data_in_field_3 ));
    LocalMux I__3162 (
            .O(N__18631),
            .I(\c0.data_in_field_3 ));
    InMux I__3161 (
            .O(N__18624),
            .I(N__18621));
    LocalMux I__3160 (
            .O(N__18621),
            .I(N__18617));
    InMux I__3159 (
            .O(N__18620),
            .I(N__18614));
    Odrv4 I__3158 (
            .O(N__18617),
            .I(\c0.n2125 ));
    LocalMux I__3157 (
            .O(N__18614),
            .I(\c0.n2125 ));
    InMux I__3156 (
            .O(N__18609),
            .I(N__18606));
    LocalMux I__3155 (
            .O(N__18606),
            .I(N__18602));
    InMux I__3154 (
            .O(N__18605),
            .I(N__18598));
    Span4Mux_v I__3153 (
            .O(N__18602),
            .I(N__18595));
    InMux I__3152 (
            .O(N__18601),
            .I(N__18592));
    LocalMux I__3151 (
            .O(N__18598),
            .I(\c0.data_in_field_27 ));
    Odrv4 I__3150 (
            .O(N__18595),
            .I(\c0.data_in_field_27 ));
    LocalMux I__3149 (
            .O(N__18592),
            .I(\c0.data_in_field_27 ));
    InMux I__3148 (
            .O(N__18585),
            .I(N__18582));
    LocalMux I__3147 (
            .O(N__18582),
            .I(\c0.n5469 ));
    CascadeMux I__3146 (
            .O(N__18579),
            .I(N__18574));
    InMux I__3145 (
            .O(N__18578),
            .I(N__18569));
    InMux I__3144 (
            .O(N__18577),
            .I(N__18566));
    InMux I__3143 (
            .O(N__18574),
            .I(N__18563));
    InMux I__3142 (
            .O(N__18573),
            .I(N__18560));
    InMux I__3141 (
            .O(N__18572),
            .I(N__18557));
    LocalMux I__3140 (
            .O(N__18569),
            .I(N__18552));
    LocalMux I__3139 (
            .O(N__18566),
            .I(N__18552));
    LocalMux I__3138 (
            .O(N__18563),
            .I(N__18547));
    LocalMux I__3137 (
            .O(N__18560),
            .I(N__18547));
    LocalMux I__3136 (
            .O(N__18557),
            .I(\c0.data_in_field_83 ));
    Odrv4 I__3135 (
            .O(N__18552),
            .I(\c0.data_in_field_83 ));
    Odrv12 I__3134 (
            .O(N__18547),
            .I(\c0.data_in_field_83 ));
    InMux I__3133 (
            .O(N__18540),
            .I(N__18537));
    LocalMux I__3132 (
            .O(N__18537),
            .I(N__18534));
    Span4Mux_v I__3131 (
            .O(N__18534),
            .I(N__18531));
    Span4Mux_h I__3130 (
            .O(N__18531),
            .I(N__18528));
    Odrv4 I__3129 (
            .O(N__18528),
            .I(\c0.n5454 ));
    CascadeMux I__3128 (
            .O(N__18525),
            .I(\c0.n5469_cascade_ ));
    InMux I__3127 (
            .O(N__18522),
            .I(N__18519));
    LocalMux I__3126 (
            .O(N__18519),
            .I(\c0.n6_adj_1923 ));
    CascadeMux I__3125 (
            .O(N__18516),
            .I(\c0.n5548_cascade_ ));
    InMux I__3124 (
            .O(N__18513),
            .I(N__18510));
    LocalMux I__3123 (
            .O(N__18510),
            .I(N__18505));
    InMux I__3122 (
            .O(N__18509),
            .I(N__18500));
    InMux I__3121 (
            .O(N__18508),
            .I(N__18500));
    Odrv4 I__3120 (
            .O(N__18505),
            .I(data_in_0_4));
    LocalMux I__3119 (
            .O(N__18500),
            .I(data_in_0_4));
    CascadeMux I__3118 (
            .O(N__18495),
            .I(N__18492));
    InMux I__3117 (
            .O(N__18492),
            .I(N__18489));
    LocalMux I__3116 (
            .O(N__18489),
            .I(N__18484));
    InMux I__3115 (
            .O(N__18488),
            .I(N__18479));
    InMux I__3114 (
            .O(N__18487),
            .I(N__18479));
    Odrv12 I__3113 (
            .O(N__18484),
            .I(data_in_7_5));
    LocalMux I__3112 (
            .O(N__18479),
            .I(data_in_7_5));
    CascadeMux I__3111 (
            .O(N__18474),
            .I(\c0.n1729_cascade_ ));
    InMux I__3110 (
            .O(N__18471),
            .I(N__18467));
    InMux I__3109 (
            .O(N__18470),
            .I(N__18461));
    LocalMux I__3108 (
            .O(N__18467),
            .I(N__18458));
    InMux I__3107 (
            .O(N__18466),
            .I(N__18455));
    InMux I__3106 (
            .O(N__18465),
            .I(N__18452));
    InMux I__3105 (
            .O(N__18464),
            .I(N__18449));
    LocalMux I__3104 (
            .O(N__18461),
            .I(N__18446));
    Span12Mux_v I__3103 (
            .O(N__18458),
            .I(N__18441));
    LocalMux I__3102 (
            .O(N__18455),
            .I(N__18441));
    LocalMux I__3101 (
            .O(N__18452),
            .I(\c0.data_in_field_35 ));
    LocalMux I__3100 (
            .O(N__18449),
            .I(\c0.data_in_field_35 ));
    Odrv4 I__3099 (
            .O(N__18446),
            .I(\c0.data_in_field_35 ));
    Odrv12 I__3098 (
            .O(N__18441),
            .I(\c0.data_in_field_35 ));
    InMux I__3097 (
            .O(N__18432),
            .I(N__18427));
    InMux I__3096 (
            .O(N__18431),
            .I(N__18424));
    InMux I__3095 (
            .O(N__18430),
            .I(N__18420));
    LocalMux I__3094 (
            .O(N__18427),
            .I(N__18417));
    LocalMux I__3093 (
            .O(N__18424),
            .I(N__18414));
    CascadeMux I__3092 (
            .O(N__18423),
            .I(N__18411));
    LocalMux I__3091 (
            .O(N__18420),
            .I(N__18408));
    Span4Mux_v I__3090 (
            .O(N__18417),
            .I(N__18403));
    Span4Mux_h I__3089 (
            .O(N__18414),
            .I(N__18403));
    InMux I__3088 (
            .O(N__18411),
            .I(N__18399));
    Span4Mux_h I__3087 (
            .O(N__18408),
            .I(N__18396));
    Span4Mux_v I__3086 (
            .O(N__18403),
            .I(N__18393));
    InMux I__3085 (
            .O(N__18402),
            .I(N__18390));
    LocalMux I__3084 (
            .O(N__18399),
            .I(\c0.data_in_field_9 ));
    Odrv4 I__3083 (
            .O(N__18396),
            .I(\c0.data_in_field_9 ));
    Odrv4 I__3082 (
            .O(N__18393),
            .I(\c0.data_in_field_9 ));
    LocalMux I__3081 (
            .O(N__18390),
            .I(\c0.data_in_field_9 ));
    InMux I__3080 (
            .O(N__18381),
            .I(N__18377));
    InMux I__3079 (
            .O(N__18380),
            .I(N__18374));
    LocalMux I__3078 (
            .O(N__18377),
            .I(N__18371));
    LocalMux I__3077 (
            .O(N__18374),
            .I(N__18368));
    Span4Mux_s3_h I__3076 (
            .O(N__18371),
            .I(N__18365));
    Span4Mux_v I__3075 (
            .O(N__18368),
            .I(N__18362));
    Span4Mux_v I__3074 (
            .O(N__18365),
            .I(N__18359));
    Span4Mux_h I__3073 (
            .O(N__18362),
            .I(N__18354));
    Span4Mux_v I__3072 (
            .O(N__18359),
            .I(N__18351));
    InMux I__3071 (
            .O(N__18358),
            .I(N__18346));
    InMux I__3070 (
            .O(N__18357),
            .I(N__18346));
    Odrv4 I__3069 (
            .O(N__18354),
            .I(\c0.data_in_field_54 ));
    Odrv4 I__3068 (
            .O(N__18351),
            .I(\c0.data_in_field_54 ));
    LocalMux I__3067 (
            .O(N__18346),
            .I(\c0.data_in_field_54 ));
    CascadeMux I__3066 (
            .O(N__18339),
            .I(\c0.n5369_cascade_ ));
    CascadeMux I__3065 (
            .O(N__18336),
            .I(N__18333));
    InMux I__3064 (
            .O(N__18333),
            .I(N__18330));
    LocalMux I__3063 (
            .O(N__18330),
            .I(N__18325));
    InMux I__3062 (
            .O(N__18329),
            .I(N__18322));
    InMux I__3061 (
            .O(N__18328),
            .I(N__18319));
    Odrv4 I__3060 (
            .O(N__18325),
            .I(data_in_0_3));
    LocalMux I__3059 (
            .O(N__18322),
            .I(data_in_0_3));
    LocalMux I__3058 (
            .O(N__18319),
            .I(data_in_0_3));
    InMux I__3057 (
            .O(N__18312),
            .I(N__18309));
    LocalMux I__3056 (
            .O(N__18309),
            .I(\c0.n26 ));
    InMux I__3055 (
            .O(N__18306),
            .I(N__18303));
    LocalMux I__3054 (
            .O(N__18303),
            .I(\c0.n27_adj_1928 ));
    CascadeMux I__3053 (
            .O(N__18300),
            .I(\c0.n28_adj_1926_cascade_ ));
    InMux I__3052 (
            .O(N__18297),
            .I(N__18294));
    LocalMux I__3051 (
            .O(N__18294),
            .I(\c0.n25_adj_1929 ));
    CascadeMux I__3050 (
            .O(N__18291),
            .I(N__18287));
    InMux I__3049 (
            .O(N__18290),
            .I(N__18283));
    InMux I__3048 (
            .O(N__18287),
            .I(N__18280));
    InMux I__3047 (
            .O(N__18286),
            .I(N__18276));
    LocalMux I__3046 (
            .O(N__18283),
            .I(N__18273));
    LocalMux I__3045 (
            .O(N__18280),
            .I(N__18270));
    InMux I__3044 (
            .O(N__18279),
            .I(N__18267));
    LocalMux I__3043 (
            .O(N__18276),
            .I(N__18262));
    Span4Mux_v I__3042 (
            .O(N__18273),
            .I(N__18262));
    Span4Mux_v I__3041 (
            .O(N__18270),
            .I(N__18259));
    LocalMux I__3040 (
            .O(N__18267),
            .I(data_in_2_1));
    Odrv4 I__3039 (
            .O(N__18262),
            .I(data_in_2_1));
    Odrv4 I__3038 (
            .O(N__18259),
            .I(data_in_2_1));
    InMux I__3037 (
            .O(N__18252),
            .I(N__18249));
    LocalMux I__3036 (
            .O(N__18249),
            .I(N__18245));
    InMux I__3035 (
            .O(N__18248),
            .I(N__18242));
    Span4Mux_v I__3034 (
            .O(N__18245),
            .I(N__18237));
    LocalMux I__3033 (
            .O(N__18242),
            .I(N__18237));
    Span4Mux_h I__3032 (
            .O(N__18237),
            .I(N__18232));
    InMux I__3031 (
            .O(N__18236),
            .I(N__18229));
    InMux I__3030 (
            .O(N__18235),
            .I(N__18226));
    Odrv4 I__3029 (
            .O(N__18232),
            .I(data_in_1_0));
    LocalMux I__3028 (
            .O(N__18229),
            .I(data_in_1_0));
    LocalMux I__3027 (
            .O(N__18226),
            .I(data_in_1_0));
    InMux I__3026 (
            .O(N__18219),
            .I(N__18216));
    LocalMux I__3025 (
            .O(N__18216),
            .I(N__18213));
    Span4Mux_v I__3024 (
            .O(N__18213),
            .I(N__18208));
    InMux I__3023 (
            .O(N__18212),
            .I(N__18203));
    InMux I__3022 (
            .O(N__18211),
            .I(N__18203));
    Odrv4 I__3021 (
            .O(N__18208),
            .I(data_in_0_6));
    LocalMux I__3020 (
            .O(N__18203),
            .I(data_in_0_6));
    InMux I__3019 (
            .O(N__18198),
            .I(N__18195));
    LocalMux I__3018 (
            .O(N__18195),
            .I(N__18190));
    InMux I__3017 (
            .O(N__18194),
            .I(N__18187));
    InMux I__3016 (
            .O(N__18193),
            .I(N__18183));
    Span4Mux_v I__3015 (
            .O(N__18190),
            .I(N__18180));
    LocalMux I__3014 (
            .O(N__18187),
            .I(N__18177));
    InMux I__3013 (
            .O(N__18186),
            .I(N__18174));
    LocalMux I__3012 (
            .O(N__18183),
            .I(N__18171));
    Odrv4 I__3011 (
            .O(N__18180),
            .I(data_in_3_7));
    Odrv4 I__3010 (
            .O(N__18177),
            .I(data_in_3_7));
    LocalMux I__3009 (
            .O(N__18174),
            .I(data_in_3_7));
    Odrv4 I__3008 (
            .O(N__18171),
            .I(data_in_3_7));
    CascadeMux I__3007 (
            .O(N__18162),
            .I(N__18159));
    InMux I__3006 (
            .O(N__18159),
            .I(N__18156));
    LocalMux I__3005 (
            .O(N__18156),
            .I(N__18153));
    Span4Mux_v I__3004 (
            .O(N__18153),
            .I(N__18147));
    InMux I__3003 (
            .O(N__18152),
            .I(N__18140));
    InMux I__3002 (
            .O(N__18151),
            .I(N__18140));
    InMux I__3001 (
            .O(N__18150),
            .I(N__18140));
    Odrv4 I__3000 (
            .O(N__18147),
            .I(data_in_1_6));
    LocalMux I__2999 (
            .O(N__18140),
            .I(data_in_1_6));
    InMux I__2998 (
            .O(N__18135),
            .I(N__18128));
    InMux I__2997 (
            .O(N__18134),
            .I(N__18128));
    InMux I__2996 (
            .O(N__18133),
            .I(N__18125));
    LocalMux I__2995 (
            .O(N__18128),
            .I(N__18122));
    LocalMux I__2994 (
            .O(N__18125),
            .I(N__18116));
    Span4Mux_v I__2993 (
            .O(N__18122),
            .I(N__18116));
    InMux I__2992 (
            .O(N__18121),
            .I(N__18113));
    Span4Mux_h I__2991 (
            .O(N__18116),
            .I(N__18110));
    LocalMux I__2990 (
            .O(N__18113),
            .I(data_in_1_7));
    Odrv4 I__2989 (
            .O(N__18110),
            .I(data_in_1_7));
    InMux I__2988 (
            .O(N__18105),
            .I(N__18101));
    CascadeMux I__2987 (
            .O(N__18104),
            .I(N__18097));
    LocalMux I__2986 (
            .O(N__18101),
            .I(N__18094));
    InMux I__2985 (
            .O(N__18100),
            .I(N__18089));
    InMux I__2984 (
            .O(N__18097),
            .I(N__18089));
    Odrv4 I__2983 (
            .O(N__18094),
            .I(data_in_0_7));
    LocalMux I__2982 (
            .O(N__18089),
            .I(data_in_0_7));
    InMux I__2981 (
            .O(N__18084),
            .I(N__18081));
    LocalMux I__2980 (
            .O(N__18081),
            .I(\c0.n30_adj_1941 ));
    InMux I__2979 (
            .O(N__18078),
            .I(N__18075));
    LocalMux I__2978 (
            .O(N__18075),
            .I(\c0.n4795 ));
    CascadeMux I__2977 (
            .O(N__18072),
            .I(N__18069));
    InMux I__2976 (
            .O(N__18069),
            .I(N__18066));
    LocalMux I__2975 (
            .O(N__18066),
            .I(\c0.n26_adj_1940 ));
    InMux I__2974 (
            .O(N__18063),
            .I(N__18060));
    LocalMux I__2973 (
            .O(N__18060),
            .I(\c0.rx.n5633 ));
    InMux I__2972 (
            .O(N__18057),
            .I(N__18053));
    InMux I__2971 (
            .O(N__18056),
            .I(N__18050));
    LocalMux I__2970 (
            .O(N__18053),
            .I(N__18047));
    LocalMux I__2969 (
            .O(N__18050),
            .I(N__18044));
    Odrv4 I__2968 (
            .O(N__18047),
            .I(n3636));
    Odrv4 I__2967 (
            .O(N__18044),
            .I(n3636));
    CascadeMux I__2966 (
            .O(N__18039),
            .I(N__18036));
    InMux I__2965 (
            .O(N__18036),
            .I(N__18032));
    InMux I__2964 (
            .O(N__18035),
            .I(N__18029));
    LocalMux I__2963 (
            .O(N__18032),
            .I(\c0.rx.n3850 ));
    LocalMux I__2962 (
            .O(N__18029),
            .I(\c0.rx.n3850 ));
    CascadeMux I__2961 (
            .O(N__18024),
            .I(N__18019));
    CascadeMux I__2960 (
            .O(N__18023),
            .I(N__18013));
    CascadeMux I__2959 (
            .O(N__18022),
            .I(N__18010));
    InMux I__2958 (
            .O(N__18019),
            .I(N__18007));
    CascadeMux I__2957 (
            .O(N__18018),
            .I(N__18000));
    CascadeMux I__2956 (
            .O(N__18017),
            .I(N__17997));
    CascadeMux I__2955 (
            .O(N__18016),
            .I(N__17993));
    InMux I__2954 (
            .O(N__18013),
            .I(N__17987));
    InMux I__2953 (
            .O(N__18010),
            .I(N__17987));
    LocalMux I__2952 (
            .O(N__18007),
            .I(N__17984));
    CascadeMux I__2951 (
            .O(N__18006),
            .I(N__17980));
    CascadeMux I__2950 (
            .O(N__18005),
            .I(N__17977));
    InMux I__2949 (
            .O(N__18004),
            .I(N__17974));
    InMux I__2948 (
            .O(N__18003),
            .I(N__17967));
    InMux I__2947 (
            .O(N__18000),
            .I(N__17967));
    InMux I__2946 (
            .O(N__17997),
            .I(N__17967));
    InMux I__2945 (
            .O(N__17996),
            .I(N__17962));
    InMux I__2944 (
            .O(N__17993),
            .I(N__17962));
    InMux I__2943 (
            .O(N__17992),
            .I(N__17959));
    LocalMux I__2942 (
            .O(N__17987),
            .I(N__17956));
    Span4Mux_h I__2941 (
            .O(N__17984),
            .I(N__17953));
    InMux I__2940 (
            .O(N__17983),
            .I(N__17946));
    InMux I__2939 (
            .O(N__17980),
            .I(N__17946));
    InMux I__2938 (
            .O(N__17977),
            .I(N__17946));
    LocalMux I__2937 (
            .O(N__17974),
            .I(r_SM_Main_1_adj_1990));
    LocalMux I__2936 (
            .O(N__17967),
            .I(r_SM_Main_1_adj_1990));
    LocalMux I__2935 (
            .O(N__17962),
            .I(r_SM_Main_1_adj_1990));
    LocalMux I__2934 (
            .O(N__17959),
            .I(r_SM_Main_1_adj_1990));
    Odrv12 I__2933 (
            .O(N__17956),
            .I(r_SM_Main_1_adj_1990));
    Odrv4 I__2932 (
            .O(N__17953),
            .I(r_SM_Main_1_adj_1990));
    LocalMux I__2931 (
            .O(N__17946),
            .I(r_SM_Main_1_adj_1990));
    CascadeMux I__2930 (
            .O(N__17931),
            .I(\c0.rx.n3850_cascade_ ));
    CEMux I__2929 (
            .O(N__17928),
            .I(N__17924));
    CEMux I__2928 (
            .O(N__17927),
            .I(N__17921));
    LocalMux I__2927 (
            .O(N__17924),
            .I(N__17918));
    LocalMux I__2926 (
            .O(N__17921),
            .I(N__17915));
    Span4Mux_h I__2925 (
            .O(N__17918),
            .I(N__17911));
    Span4Mux_v I__2924 (
            .O(N__17915),
            .I(N__17908));
    InMux I__2923 (
            .O(N__17914),
            .I(N__17905));
    Odrv4 I__2922 (
            .O(N__17911),
            .I(\c0.rx.n2259 ));
    Odrv4 I__2921 (
            .O(N__17908),
            .I(\c0.rx.n2259 ));
    LocalMux I__2920 (
            .O(N__17905),
            .I(\c0.rx.n2259 ));
    SRMux I__2919 (
            .O(N__17898),
            .I(N__17894));
    SRMux I__2918 (
            .O(N__17897),
            .I(N__17891));
    LocalMux I__2917 (
            .O(N__17894),
            .I(N__17888));
    LocalMux I__2916 (
            .O(N__17891),
            .I(N__17885));
    Span4Mux_h I__2915 (
            .O(N__17888),
            .I(N__17880));
    Span4Mux_h I__2914 (
            .O(N__17885),
            .I(N__17880));
    Odrv4 I__2913 (
            .O(N__17880),
            .I(\c0.rx.n2367 ));
    CascadeMux I__2912 (
            .O(N__17877),
            .I(N__17874));
    InMux I__2911 (
            .O(N__17874),
            .I(N__17871));
    LocalMux I__2910 (
            .O(N__17871),
            .I(N__17866));
    CascadeMux I__2909 (
            .O(N__17870),
            .I(N__17862));
    InMux I__2908 (
            .O(N__17869),
            .I(N__17859));
    Span4Mux_h I__2907 (
            .O(N__17866),
            .I(N__17856));
    InMux I__2906 (
            .O(N__17865),
            .I(N__17851));
    InMux I__2905 (
            .O(N__17862),
            .I(N__17851));
    LocalMux I__2904 (
            .O(N__17859),
            .I(data_in_2_5));
    Odrv4 I__2903 (
            .O(N__17856),
            .I(data_in_2_5));
    LocalMux I__2902 (
            .O(N__17851),
            .I(data_in_2_5));
    InMux I__2901 (
            .O(N__17844),
            .I(N__17841));
    LocalMux I__2900 (
            .O(N__17841),
            .I(N__17838));
    Span4Mux_v I__2899 (
            .O(N__17838),
            .I(N__17833));
    InMux I__2898 (
            .O(N__17837),
            .I(N__17828));
    InMux I__2897 (
            .O(N__17836),
            .I(N__17828));
    Span4Mux_h I__2896 (
            .O(N__17833),
            .I(N__17825));
    LocalMux I__2895 (
            .O(N__17828),
            .I(data_in_10_1));
    Odrv4 I__2894 (
            .O(N__17825),
            .I(data_in_10_1));
    InMux I__2893 (
            .O(N__17820),
            .I(N__17816));
    InMux I__2892 (
            .O(N__17819),
            .I(N__17813));
    LocalMux I__2891 (
            .O(N__17816),
            .I(N__17810));
    LocalMux I__2890 (
            .O(N__17813),
            .I(N__17805));
    Span4Mux_v I__2889 (
            .O(N__17810),
            .I(N__17805));
    Span4Mux_v I__2888 (
            .O(N__17805),
            .I(N__17801));
    InMux I__2887 (
            .O(N__17804),
            .I(N__17798));
    Odrv4 I__2886 (
            .O(N__17801),
            .I(data_in_9_1));
    LocalMux I__2885 (
            .O(N__17798),
            .I(data_in_9_1));
    CascadeMux I__2884 (
            .O(N__17793),
            .I(N__17790));
    InMux I__2883 (
            .O(N__17790),
            .I(N__17787));
    LocalMux I__2882 (
            .O(N__17787),
            .I(N__17784));
    Span4Mux_h I__2881 (
            .O(N__17784),
            .I(N__17779));
    InMux I__2880 (
            .O(N__17783),
            .I(N__17774));
    InMux I__2879 (
            .O(N__17782),
            .I(N__17774));
    Odrv4 I__2878 (
            .O(N__17779),
            .I(data_in_12_6));
    LocalMux I__2877 (
            .O(N__17774),
            .I(data_in_12_6));
    InMux I__2876 (
            .O(N__17769),
            .I(N__17766));
    LocalMux I__2875 (
            .O(N__17766),
            .I(N__17763));
    Span4Mux_v I__2874 (
            .O(N__17763),
            .I(N__17760));
    Span4Mux_v I__2873 (
            .O(N__17760),
            .I(N__17756));
    InMux I__2872 (
            .O(N__17759),
            .I(N__17753));
    Odrv4 I__2871 (
            .O(N__17756),
            .I(n1764));
    LocalMux I__2870 (
            .O(N__17753),
            .I(n1764));
    InMux I__2869 (
            .O(N__17748),
            .I(N__17744));
    CascadeMux I__2868 (
            .O(N__17747),
            .I(N__17741));
    LocalMux I__2867 (
            .O(N__17744),
            .I(N__17738));
    InMux I__2866 (
            .O(N__17741),
            .I(N__17735));
    Odrv4 I__2865 (
            .O(N__17738),
            .I(rx_data_7));
    LocalMux I__2864 (
            .O(N__17735),
            .I(rx_data_7));
    InMux I__2863 (
            .O(N__17730),
            .I(N__17727));
    LocalMux I__2862 (
            .O(N__17727),
            .I(N__17723));
    InMux I__2861 (
            .O(N__17726),
            .I(N__17720));
    Span4Mux_h I__2860 (
            .O(N__17723),
            .I(N__17717));
    LocalMux I__2859 (
            .O(N__17720),
            .I(N__17714));
    Span4Mux_v I__2858 (
            .O(N__17717),
            .I(N__17709));
    Span4Mux_h I__2857 (
            .O(N__17714),
            .I(N__17709));
    Span4Mux_h I__2856 (
            .O(N__17709),
            .I(N__17705));
    InMux I__2855 (
            .O(N__17708),
            .I(N__17702));
    Odrv4 I__2854 (
            .O(N__17705),
            .I(data_in_15_6));
    LocalMux I__2853 (
            .O(N__17702),
            .I(data_in_15_6));
    CascadeMux I__2852 (
            .O(N__17697),
            .I(N__17692));
    CascadeMux I__2851 (
            .O(N__17696),
            .I(N__17685));
    InMux I__2850 (
            .O(N__17695),
            .I(N__17680));
    InMux I__2849 (
            .O(N__17692),
            .I(N__17675));
    InMux I__2848 (
            .O(N__17691),
            .I(N__17675));
    InMux I__2847 (
            .O(N__17690),
            .I(N__17670));
    InMux I__2846 (
            .O(N__17689),
            .I(N__17670));
    InMux I__2845 (
            .O(N__17688),
            .I(N__17667));
    InMux I__2844 (
            .O(N__17685),
            .I(N__17660));
    InMux I__2843 (
            .O(N__17684),
            .I(N__17660));
    InMux I__2842 (
            .O(N__17683),
            .I(N__17660));
    LocalMux I__2841 (
            .O(N__17680),
            .I(N__17655));
    LocalMux I__2840 (
            .O(N__17675),
            .I(N__17655));
    LocalMux I__2839 (
            .O(N__17670),
            .I(r_SM_Main_0_adj_1991));
    LocalMux I__2838 (
            .O(N__17667),
            .I(r_SM_Main_0_adj_1991));
    LocalMux I__2837 (
            .O(N__17660),
            .I(r_SM_Main_0_adj_1991));
    Odrv4 I__2836 (
            .O(N__17655),
            .I(r_SM_Main_0_adj_1991));
    InMux I__2835 (
            .O(N__17646),
            .I(N__17642));
    InMux I__2834 (
            .O(N__17645),
            .I(N__17639));
    LocalMux I__2833 (
            .O(N__17642),
            .I(N__17631));
    LocalMux I__2832 (
            .O(N__17639),
            .I(N__17627));
    InMux I__2831 (
            .O(N__17638),
            .I(N__17622));
    InMux I__2830 (
            .O(N__17637),
            .I(N__17622));
    InMux I__2829 (
            .O(N__17636),
            .I(N__17615));
    InMux I__2828 (
            .O(N__17635),
            .I(N__17615));
    InMux I__2827 (
            .O(N__17634),
            .I(N__17615));
    Span4Mux_h I__2826 (
            .O(N__17631),
            .I(N__17612));
    InMux I__2825 (
            .O(N__17630),
            .I(N__17609));
    Odrv4 I__2824 (
            .O(N__17627),
            .I(r_SM_Main_2_N_1824_2));
    LocalMux I__2823 (
            .O(N__17622),
            .I(r_SM_Main_2_N_1824_2));
    LocalMux I__2822 (
            .O(N__17615),
            .I(r_SM_Main_2_N_1824_2));
    Odrv4 I__2821 (
            .O(N__17612),
            .I(r_SM_Main_2_N_1824_2));
    LocalMux I__2820 (
            .O(N__17609),
            .I(r_SM_Main_2_N_1824_2));
    InMux I__2819 (
            .O(N__17598),
            .I(N__17595));
    LocalMux I__2818 (
            .O(N__17595),
            .I(\c0.rx.n6291 ));
    InMux I__2817 (
            .O(N__17592),
            .I(N__17589));
    LocalMux I__2816 (
            .O(N__17589),
            .I(N__17585));
    InMux I__2815 (
            .O(N__17588),
            .I(N__17582));
    Odrv4 I__2814 (
            .O(N__17585),
            .I(\c0.n1889 ));
    LocalMux I__2813 (
            .O(N__17582),
            .I(\c0.n1889 ));
    InMux I__2812 (
            .O(N__17577),
            .I(N__17573));
    CascadeMux I__2811 (
            .O(N__17576),
            .I(N__17570));
    LocalMux I__2810 (
            .O(N__17573),
            .I(N__17567));
    InMux I__2809 (
            .O(N__17570),
            .I(N__17561));
    Span4Mux_v I__2808 (
            .O(N__17567),
            .I(N__17558));
    InMux I__2807 (
            .O(N__17566),
            .I(N__17551));
    InMux I__2806 (
            .O(N__17565),
            .I(N__17551));
    InMux I__2805 (
            .O(N__17564),
            .I(N__17551));
    LocalMux I__2804 (
            .O(N__17561),
            .I(\c0.data_in_field_76 ));
    Odrv4 I__2803 (
            .O(N__17558),
            .I(\c0.data_in_field_76 ));
    LocalMux I__2802 (
            .O(N__17551),
            .I(\c0.data_in_field_76 ));
    InMux I__2801 (
            .O(N__17544),
            .I(N__17540));
    InMux I__2800 (
            .O(N__17543),
            .I(N__17537));
    LocalMux I__2799 (
            .O(N__17540),
            .I(N__17534));
    LocalMux I__2798 (
            .O(N__17537),
            .I(\c0.data_in_frame_18_4 ));
    Odrv4 I__2797 (
            .O(N__17534),
            .I(\c0.data_in_frame_18_4 ));
    CascadeMux I__2796 (
            .O(N__17529),
            .I(\c0.n6243_cascade_ ));
    CascadeMux I__2795 (
            .O(N__17526),
            .I(\c0.n5698_cascade_ ));
    InMux I__2794 (
            .O(N__17523),
            .I(N__17520));
    LocalMux I__2793 (
            .O(N__17520),
            .I(N__17517));
    Odrv4 I__2792 (
            .O(N__17517),
            .I(\c0.n6231 ));
    InMux I__2791 (
            .O(N__17514),
            .I(N__17511));
    LocalMux I__2790 (
            .O(N__17511),
            .I(\c0.n6237 ));
    CascadeMux I__2789 (
            .O(N__17508),
            .I(N__17505));
    InMux I__2788 (
            .O(N__17505),
            .I(N__17501));
    InMux I__2787 (
            .O(N__17504),
            .I(N__17496));
    LocalMux I__2786 (
            .O(N__17501),
            .I(N__17493));
    InMux I__2785 (
            .O(N__17500),
            .I(N__17488));
    InMux I__2784 (
            .O(N__17499),
            .I(N__17488));
    LocalMux I__2783 (
            .O(N__17496),
            .I(\c0.data_in_field_102 ));
    Odrv4 I__2782 (
            .O(N__17493),
            .I(\c0.data_in_field_102 ));
    LocalMux I__2781 (
            .O(N__17488),
            .I(\c0.data_in_field_102 ));
    InMux I__2780 (
            .O(N__17481),
            .I(N__17478));
    LocalMux I__2779 (
            .O(N__17478),
            .I(\c0.n5701 ));
    InMux I__2778 (
            .O(N__17475),
            .I(N__17471));
    InMux I__2777 (
            .O(N__17474),
            .I(N__17468));
    LocalMux I__2776 (
            .O(N__17471),
            .I(N__17465));
    LocalMux I__2775 (
            .O(N__17468),
            .I(N__17462));
    Span4Mux_v I__2774 (
            .O(N__17465),
            .I(N__17458));
    Span12Mux_v I__2773 (
            .O(N__17462),
            .I(N__17455));
    InMux I__2772 (
            .O(N__17461),
            .I(N__17452));
    Odrv4 I__2771 (
            .O(N__17458),
            .I(data_in_10_6));
    Odrv12 I__2770 (
            .O(N__17455),
            .I(data_in_10_6));
    LocalMux I__2769 (
            .O(N__17452),
            .I(data_in_10_6));
    InMux I__2768 (
            .O(N__17445),
            .I(N__17442));
    LocalMux I__2767 (
            .O(N__17442),
            .I(N__17436));
    InMux I__2766 (
            .O(N__17441),
            .I(N__17432));
    InMux I__2765 (
            .O(N__17440),
            .I(N__17427));
    InMux I__2764 (
            .O(N__17439),
            .I(N__17427));
    Span4Mux_v I__2763 (
            .O(N__17436),
            .I(N__17424));
    InMux I__2762 (
            .O(N__17435),
            .I(N__17421));
    LocalMux I__2761 (
            .O(N__17432),
            .I(N__17418));
    LocalMux I__2760 (
            .O(N__17427),
            .I(\c0.data_in_field_86 ));
    Odrv4 I__2759 (
            .O(N__17424),
            .I(\c0.data_in_field_86 ));
    LocalMux I__2758 (
            .O(N__17421),
            .I(\c0.data_in_field_86 ));
    Odrv4 I__2757 (
            .O(N__17418),
            .I(\c0.data_in_field_86 ));
    CascadeMux I__2756 (
            .O(N__17409),
            .I(N__17406));
    InMux I__2755 (
            .O(N__17406),
            .I(N__17403));
    LocalMux I__2754 (
            .O(N__17403),
            .I(\c0.n5388 ));
    InMux I__2753 (
            .O(N__17400),
            .I(N__17397));
    LocalMux I__2752 (
            .O(N__17397),
            .I(\c0.n5418 ));
    InMux I__2751 (
            .O(N__17394),
            .I(N__17391));
    LocalMux I__2750 (
            .O(N__17391),
            .I(N__17387));
    InMux I__2749 (
            .O(N__17390),
            .I(N__17384));
    Odrv4 I__2748 (
            .O(N__17387),
            .I(\c0.n5491 ));
    LocalMux I__2747 (
            .O(N__17384),
            .I(\c0.n5491 ));
    InMux I__2746 (
            .O(N__17379),
            .I(N__17376));
    LocalMux I__2745 (
            .O(N__17376),
            .I(\c0.n44_adj_1894 ));
    InMux I__2744 (
            .O(N__17373),
            .I(N__17368));
    InMux I__2743 (
            .O(N__17372),
            .I(N__17365));
    InMux I__2742 (
            .O(N__17371),
            .I(N__17362));
    LocalMux I__2741 (
            .O(N__17368),
            .I(\c0.data_in_field_112 ));
    LocalMux I__2740 (
            .O(N__17365),
            .I(\c0.data_in_field_112 ));
    LocalMux I__2739 (
            .O(N__17362),
            .I(\c0.data_in_field_112 ));
    CascadeMux I__2738 (
            .O(N__17355),
            .I(N__17350));
    InMux I__2737 (
            .O(N__17354),
            .I(N__17347));
    CascadeMux I__2736 (
            .O(N__17353),
            .I(N__17343));
    InMux I__2735 (
            .O(N__17350),
            .I(N__17340));
    LocalMux I__2734 (
            .O(N__17347),
            .I(N__17337));
    InMux I__2733 (
            .O(N__17346),
            .I(N__17334));
    InMux I__2732 (
            .O(N__17343),
            .I(N__17331));
    LocalMux I__2731 (
            .O(N__17340),
            .I(\c0.data_in_field_30 ));
    Odrv4 I__2730 (
            .O(N__17337),
            .I(\c0.data_in_field_30 ));
    LocalMux I__2729 (
            .O(N__17334),
            .I(\c0.data_in_field_30 ));
    LocalMux I__2728 (
            .O(N__17331),
            .I(\c0.data_in_field_30 ));
    InMux I__2727 (
            .O(N__17322),
            .I(N__17319));
    LocalMux I__2726 (
            .O(N__17319),
            .I(N__17315));
    InMux I__2725 (
            .O(N__17318),
            .I(N__17312));
    Span4Mux_v I__2724 (
            .O(N__17315),
            .I(N__17304));
    LocalMux I__2723 (
            .O(N__17312),
            .I(N__17304));
    InMux I__2722 (
            .O(N__17311),
            .I(N__17301));
    InMux I__2721 (
            .O(N__17310),
            .I(N__17296));
    InMux I__2720 (
            .O(N__17309),
            .I(N__17296));
    Odrv4 I__2719 (
            .O(N__17304),
            .I(\c0.data_in_field_125 ));
    LocalMux I__2718 (
            .O(N__17301),
            .I(\c0.data_in_field_125 ));
    LocalMux I__2717 (
            .O(N__17296),
            .I(\c0.data_in_field_125 ));
    InMux I__2716 (
            .O(N__17289),
            .I(N__17286));
    LocalMux I__2715 (
            .O(N__17286),
            .I(N__17280));
    InMux I__2714 (
            .O(N__17285),
            .I(N__17277));
    InMux I__2713 (
            .O(N__17284),
            .I(N__17274));
    CascadeMux I__2712 (
            .O(N__17283),
            .I(N__17270));
    Span4Mux_s2_h I__2711 (
            .O(N__17280),
            .I(N__17265));
    LocalMux I__2710 (
            .O(N__17277),
            .I(N__17265));
    LocalMux I__2709 (
            .O(N__17274),
            .I(N__17262));
    InMux I__2708 (
            .O(N__17273),
            .I(N__17259));
    InMux I__2707 (
            .O(N__17270),
            .I(N__17256));
    Span4Mux_h I__2706 (
            .O(N__17265),
            .I(N__17253));
    Span4Mux_h I__2705 (
            .O(N__17262),
            .I(N__17248));
    LocalMux I__2704 (
            .O(N__17259),
            .I(N__17248));
    LocalMux I__2703 (
            .O(N__17256),
            .I(\c0.data_in_field_135 ));
    Odrv4 I__2702 (
            .O(N__17253),
            .I(\c0.data_in_field_135 ));
    Odrv4 I__2701 (
            .O(N__17248),
            .I(\c0.data_in_field_135 ));
    InMux I__2700 (
            .O(N__17241),
            .I(N__17238));
    LocalMux I__2699 (
            .O(N__17238),
            .I(N__17234));
    InMux I__2698 (
            .O(N__17237),
            .I(N__17231));
    Span4Mux_h I__2697 (
            .O(N__17234),
            .I(N__17228));
    LocalMux I__2696 (
            .O(N__17231),
            .I(\c0.n1908 ));
    Odrv4 I__2695 (
            .O(N__17228),
            .I(\c0.n1908 ));
    InMux I__2694 (
            .O(N__17223),
            .I(N__17220));
    LocalMux I__2693 (
            .O(N__17220),
            .I(N__17216));
    InMux I__2692 (
            .O(N__17219),
            .I(N__17213));
    Span4Mux_v I__2691 (
            .O(N__17216),
            .I(N__17204));
    LocalMux I__2690 (
            .O(N__17213),
            .I(N__17204));
    InMux I__2689 (
            .O(N__17212),
            .I(N__17201));
    InMux I__2688 (
            .O(N__17211),
            .I(N__17198));
    InMux I__2687 (
            .O(N__17210),
            .I(N__17195));
    CascadeMux I__2686 (
            .O(N__17209),
            .I(N__17192));
    Span4Mux_v I__2685 (
            .O(N__17204),
            .I(N__17187));
    LocalMux I__2684 (
            .O(N__17201),
            .I(N__17187));
    LocalMux I__2683 (
            .O(N__17198),
            .I(N__17182));
    LocalMux I__2682 (
            .O(N__17195),
            .I(N__17182));
    InMux I__2681 (
            .O(N__17192),
            .I(N__17179));
    Span4Mux_h I__2680 (
            .O(N__17187),
            .I(N__17176));
    Span4Mux_v I__2679 (
            .O(N__17182),
            .I(N__17173));
    LocalMux I__2678 (
            .O(N__17179),
            .I(\c0.data_in_field_99 ));
    Odrv4 I__2677 (
            .O(N__17176),
            .I(\c0.data_in_field_99 ));
    Odrv4 I__2676 (
            .O(N__17173),
            .I(\c0.data_in_field_99 ));
    InMux I__2675 (
            .O(N__17166),
            .I(N__17163));
    LocalMux I__2674 (
            .O(N__17163),
            .I(N__17159));
    InMux I__2673 (
            .O(N__17162),
            .I(N__17156));
    Span4Mux_v I__2672 (
            .O(N__17159),
            .I(N__17150));
    LocalMux I__2671 (
            .O(N__17156),
            .I(N__17147));
    InMux I__2670 (
            .O(N__17155),
            .I(N__17140));
    InMux I__2669 (
            .O(N__17154),
            .I(N__17140));
    InMux I__2668 (
            .O(N__17153),
            .I(N__17140));
    Odrv4 I__2667 (
            .O(N__17150),
            .I(\c0.data_in_field_65 ));
    Odrv12 I__2666 (
            .O(N__17147),
            .I(\c0.data_in_field_65 ));
    LocalMux I__2665 (
            .O(N__17140),
            .I(\c0.data_in_field_65 ));
    InMux I__2664 (
            .O(N__17133),
            .I(N__17130));
    LocalMux I__2663 (
            .O(N__17130),
            .I(N__17127));
    Span4Mux_v I__2662 (
            .O(N__17127),
            .I(N__17121));
    InMux I__2661 (
            .O(N__17126),
            .I(N__17118));
    InMux I__2660 (
            .O(N__17125),
            .I(N__17113));
    InMux I__2659 (
            .O(N__17124),
            .I(N__17113));
    Odrv4 I__2658 (
            .O(N__17121),
            .I(\c0.data_in_field_129 ));
    LocalMux I__2657 (
            .O(N__17118),
            .I(\c0.data_in_field_129 ));
    LocalMux I__2656 (
            .O(N__17113),
            .I(\c0.data_in_field_129 ));
    InMux I__2655 (
            .O(N__17106),
            .I(N__17103));
    LocalMux I__2654 (
            .O(N__17103),
            .I(N__17100));
    Span4Mux_h I__2653 (
            .O(N__17100),
            .I(N__17097));
    Odrv4 I__2652 (
            .O(N__17097),
            .I(\c0.n5569 ));
    CascadeMux I__2651 (
            .O(N__17094),
            .I(\c0.n5569_cascade_ ));
    InMux I__2650 (
            .O(N__17091),
            .I(N__17088));
    LocalMux I__2649 (
            .O(N__17088),
            .I(N__17082));
    CascadeMux I__2648 (
            .O(N__17087),
            .I(N__17079));
    InMux I__2647 (
            .O(N__17086),
            .I(N__17076));
    InMux I__2646 (
            .O(N__17085),
            .I(N__17073));
    Span4Mux_h I__2645 (
            .O(N__17082),
            .I(N__17070));
    InMux I__2644 (
            .O(N__17079),
            .I(N__17067));
    LocalMux I__2643 (
            .O(N__17076),
            .I(\c0.data_in_field_114 ));
    LocalMux I__2642 (
            .O(N__17073),
            .I(\c0.data_in_field_114 ));
    Odrv4 I__2641 (
            .O(N__17070),
            .I(\c0.data_in_field_114 ));
    LocalMux I__2640 (
            .O(N__17067),
            .I(\c0.data_in_field_114 ));
    InMux I__2639 (
            .O(N__17058),
            .I(N__17055));
    LocalMux I__2638 (
            .O(N__17055),
            .I(N__17052));
    Span4Mux_v I__2637 (
            .O(N__17052),
            .I(N__17049));
    Odrv4 I__2636 (
            .O(N__17049),
            .I(\c0.n20_adj_1882 ));
    CascadeMux I__2635 (
            .O(N__17046),
            .I(\c0.n2062_cascade_ ));
    InMux I__2634 (
            .O(N__17043),
            .I(N__17040));
    LocalMux I__2633 (
            .O(N__17040),
            .I(N__17037));
    Span4Mux_h I__2632 (
            .O(N__17037),
            .I(N__17034));
    Odrv4 I__2631 (
            .O(N__17034),
            .I(\c0.n44 ));
    InMux I__2630 (
            .O(N__17031),
            .I(N__17028));
    LocalMux I__2629 (
            .O(N__17028),
            .I(N__17023));
    InMux I__2628 (
            .O(N__17027),
            .I(N__17020));
    InMux I__2627 (
            .O(N__17026),
            .I(N__17017));
    Span4Mux_v I__2626 (
            .O(N__17023),
            .I(N__17014));
    LocalMux I__2625 (
            .O(N__17020),
            .I(N__17011));
    LocalMux I__2624 (
            .O(N__17017),
            .I(N__17007));
    Span4Mux_s2_h I__2623 (
            .O(N__17014),
            .I(N__17002));
    Span4Mux_h I__2622 (
            .O(N__17011),
            .I(N__17002));
    InMux I__2621 (
            .O(N__17010),
            .I(N__16999));
    Odrv4 I__2620 (
            .O(N__17007),
            .I(\c0.data_in_field_134 ));
    Odrv4 I__2619 (
            .O(N__17002),
            .I(\c0.data_in_field_134 ));
    LocalMux I__2618 (
            .O(N__16999),
            .I(\c0.data_in_field_134 ));
    InMux I__2617 (
            .O(N__16992),
            .I(N__16989));
    LocalMux I__2616 (
            .O(N__16989),
            .I(N__16986));
    Span4Mux_s3_h I__2615 (
            .O(N__16986),
            .I(N__16983));
    Span4Mux_v I__2614 (
            .O(N__16983),
            .I(N__16979));
    InMux I__2613 (
            .O(N__16982),
            .I(N__16976));
    Odrv4 I__2612 (
            .O(N__16979),
            .I(\c0.n5503 ));
    LocalMux I__2611 (
            .O(N__16976),
            .I(\c0.n5503 ));
    InMux I__2610 (
            .O(N__16971),
            .I(N__16968));
    LocalMux I__2609 (
            .O(N__16968),
            .I(N__16964));
    InMux I__2608 (
            .O(N__16967),
            .I(N__16961));
    Span4Mux_v I__2607 (
            .O(N__16964),
            .I(N__16958));
    LocalMux I__2606 (
            .O(N__16961),
            .I(N__16955));
    Odrv4 I__2605 (
            .O(N__16958),
            .I(\c0.n2095 ));
    Odrv12 I__2604 (
            .O(N__16955),
            .I(\c0.n2095 ));
    InMux I__2603 (
            .O(N__16950),
            .I(N__16947));
    LocalMux I__2602 (
            .O(N__16947),
            .I(\c0.n16_adj_1871 ));
    InMux I__2601 (
            .O(N__16944),
            .I(N__16940));
    InMux I__2600 (
            .O(N__16943),
            .I(N__16937));
    LocalMux I__2599 (
            .O(N__16940),
            .I(N__16934));
    LocalMux I__2598 (
            .O(N__16937),
            .I(N__16930));
    Span4Mux_v I__2597 (
            .O(N__16934),
            .I(N__16927));
    InMux I__2596 (
            .O(N__16933),
            .I(N__16924));
    Span4Mux_v I__2595 (
            .O(N__16930),
            .I(N__16921));
    Span4Mux_s2_h I__2594 (
            .O(N__16927),
            .I(N__16918));
    LocalMux I__2593 (
            .O(N__16924),
            .I(data_in_11_3));
    Odrv4 I__2592 (
            .O(N__16921),
            .I(data_in_11_3));
    Odrv4 I__2591 (
            .O(N__16918),
            .I(data_in_11_3));
    InMux I__2590 (
            .O(N__16911),
            .I(N__16908));
    LocalMux I__2589 (
            .O(N__16908),
            .I(\c0.n2021 ));
    InMux I__2588 (
            .O(N__16905),
            .I(N__16901));
    InMux I__2587 (
            .O(N__16904),
            .I(N__16898));
    LocalMux I__2586 (
            .O(N__16901),
            .I(N__16894));
    LocalMux I__2585 (
            .O(N__16898),
            .I(N__16891));
    InMux I__2584 (
            .O(N__16897),
            .I(N__16887));
    Span4Mux_h I__2583 (
            .O(N__16894),
            .I(N__16882));
    Span4Mux_h I__2582 (
            .O(N__16891),
            .I(N__16882));
    InMux I__2581 (
            .O(N__16890),
            .I(N__16879));
    LocalMux I__2580 (
            .O(N__16887),
            .I(\c0.data_in_field_10 ));
    Odrv4 I__2579 (
            .O(N__16882),
            .I(\c0.data_in_field_10 ));
    LocalMux I__2578 (
            .O(N__16879),
            .I(\c0.data_in_field_10 ));
    CascadeMux I__2577 (
            .O(N__16872),
            .I(\c0.n2021_cascade_ ));
    InMux I__2576 (
            .O(N__16869),
            .I(N__16864));
    CascadeMux I__2575 (
            .O(N__16868),
            .I(N__16861));
    InMux I__2574 (
            .O(N__16867),
            .I(N__16857));
    LocalMux I__2573 (
            .O(N__16864),
            .I(N__16854));
    InMux I__2572 (
            .O(N__16861),
            .I(N__16851));
    InMux I__2571 (
            .O(N__16860),
            .I(N__16848));
    LocalMux I__2570 (
            .O(N__16857),
            .I(\c0.data_in_field_41 ));
    Odrv12 I__2569 (
            .O(N__16854),
            .I(\c0.data_in_field_41 ));
    LocalMux I__2568 (
            .O(N__16851),
            .I(\c0.data_in_field_41 ));
    LocalMux I__2567 (
            .O(N__16848),
            .I(\c0.data_in_field_41 ));
    CascadeMux I__2566 (
            .O(N__16839),
            .I(\c0.n2074_cascade_ ));
    InMux I__2565 (
            .O(N__16836),
            .I(N__16830));
    InMux I__2564 (
            .O(N__16835),
            .I(N__16830));
    LocalMux I__2563 (
            .O(N__16830),
            .I(\c0.n2000 ));
    InMux I__2562 (
            .O(N__16827),
            .I(N__16823));
    InMux I__2561 (
            .O(N__16826),
            .I(N__16820));
    LocalMux I__2560 (
            .O(N__16823),
            .I(N__16817));
    LocalMux I__2559 (
            .O(N__16820),
            .I(N__16814));
    Span4Mux_h I__2558 (
            .O(N__16817),
            .I(N__16809));
    Span4Mux_h I__2557 (
            .O(N__16814),
            .I(N__16806));
    InMux I__2556 (
            .O(N__16813),
            .I(N__16801));
    InMux I__2555 (
            .O(N__16812),
            .I(N__16801));
    Odrv4 I__2554 (
            .O(N__16809),
            .I(\c0.data_in_field_26 ));
    Odrv4 I__2553 (
            .O(N__16806),
            .I(\c0.data_in_field_26 ));
    LocalMux I__2552 (
            .O(N__16801),
            .I(\c0.data_in_field_26 ));
    InMux I__2551 (
            .O(N__16794),
            .I(N__16791));
    LocalMux I__2550 (
            .O(N__16791),
            .I(N__16785));
    InMux I__2549 (
            .O(N__16790),
            .I(N__16782));
    InMux I__2548 (
            .O(N__16789),
            .I(N__16779));
    InMux I__2547 (
            .O(N__16788),
            .I(N__16776));
    Span4Mux_v I__2546 (
            .O(N__16785),
            .I(N__16771));
    LocalMux I__2545 (
            .O(N__16782),
            .I(N__16771));
    LocalMux I__2544 (
            .O(N__16779),
            .I(N__16768));
    LocalMux I__2543 (
            .O(N__16776),
            .I(N__16763));
    Span4Mux_h I__2542 (
            .O(N__16771),
            .I(N__16760));
    Span4Mux_h I__2541 (
            .O(N__16768),
            .I(N__16757));
    InMux I__2540 (
            .O(N__16767),
            .I(N__16752));
    InMux I__2539 (
            .O(N__16766),
            .I(N__16752));
    Odrv12 I__2538 (
            .O(N__16763),
            .I(\c0.data_in_field_64 ));
    Odrv4 I__2537 (
            .O(N__16760),
            .I(\c0.data_in_field_64 ));
    Odrv4 I__2536 (
            .O(N__16757),
            .I(\c0.data_in_field_64 ));
    LocalMux I__2535 (
            .O(N__16752),
            .I(\c0.data_in_field_64 ));
    CascadeMux I__2534 (
            .O(N__16743),
            .I(N__16740));
    InMux I__2533 (
            .O(N__16740),
            .I(N__16737));
    LocalMux I__2532 (
            .O(N__16737),
            .I(N__16733));
    InMux I__2531 (
            .O(N__16736),
            .I(N__16730));
    Span4Mux_v I__2530 (
            .O(N__16733),
            .I(N__16726));
    LocalMux I__2529 (
            .O(N__16730),
            .I(N__16723));
    InMux I__2528 (
            .O(N__16729),
            .I(N__16720));
    Odrv4 I__2527 (
            .O(N__16726),
            .I(data_in_8_2));
    Odrv4 I__2526 (
            .O(N__16723),
            .I(data_in_8_2));
    LocalMux I__2525 (
            .O(N__16720),
            .I(data_in_8_2));
    InMux I__2524 (
            .O(N__16713),
            .I(N__16709));
    CascadeMux I__2523 (
            .O(N__16712),
            .I(N__16706));
    LocalMux I__2522 (
            .O(N__16709),
            .I(N__16703));
    InMux I__2521 (
            .O(N__16706),
            .I(N__16700));
    Span4Mux_v I__2520 (
            .O(N__16703),
            .I(N__16695));
    LocalMux I__2519 (
            .O(N__16700),
            .I(N__16695));
    Span4Mux_v I__2518 (
            .O(N__16695),
            .I(N__16691));
    InMux I__2517 (
            .O(N__16694),
            .I(N__16688));
    Sp12to4 I__2516 (
            .O(N__16691),
            .I(N__16685));
    LocalMux I__2515 (
            .O(N__16688),
            .I(data_in_5_3));
    Odrv12 I__2514 (
            .O(N__16685),
            .I(data_in_5_3));
    CascadeMux I__2513 (
            .O(N__16680),
            .I(N__16677));
    InMux I__2512 (
            .O(N__16677),
            .I(N__16674));
    LocalMux I__2511 (
            .O(N__16674),
            .I(N__16671));
    Span4Mux_v I__2510 (
            .O(N__16671),
            .I(N__16668));
    Odrv4 I__2509 (
            .O(N__16668),
            .I(\c0.n6183 ));
    InMux I__2508 (
            .O(N__16665),
            .I(N__16662));
    LocalMux I__2507 (
            .O(N__16662),
            .I(\c0.n20_adj_1958 ));
    CascadeMux I__2506 (
            .O(N__16659),
            .I(\c0.n31_adj_1896_cascade_ ));
    InMux I__2505 (
            .O(N__16656),
            .I(N__16653));
    LocalMux I__2504 (
            .O(N__16653),
            .I(\c0.n41 ));
    InMux I__2503 (
            .O(N__16650),
            .I(N__16647));
    LocalMux I__2502 (
            .O(N__16647),
            .I(N__16642));
    InMux I__2501 (
            .O(N__16646),
            .I(N__16638));
    InMux I__2500 (
            .O(N__16645),
            .I(N__16635));
    Span4Mux_v I__2499 (
            .O(N__16642),
            .I(N__16632));
    InMux I__2498 (
            .O(N__16641),
            .I(N__16629));
    LocalMux I__2497 (
            .O(N__16638),
            .I(N__16626));
    LocalMux I__2496 (
            .O(N__16635),
            .I(\c0.data_in_field_6 ));
    Odrv4 I__2495 (
            .O(N__16632),
            .I(\c0.data_in_field_6 ));
    LocalMux I__2494 (
            .O(N__16629),
            .I(\c0.data_in_field_6 ));
    Odrv4 I__2493 (
            .O(N__16626),
            .I(\c0.data_in_field_6 ));
    InMux I__2492 (
            .O(N__16617),
            .I(N__16614));
    LocalMux I__2491 (
            .O(N__16614),
            .I(\c0.n10_adj_1915 ));
    InMux I__2490 (
            .O(N__16611),
            .I(N__16608));
    LocalMux I__2489 (
            .O(N__16608),
            .I(N__16605));
    Odrv4 I__2488 (
            .O(N__16605),
            .I(\c0.n1913 ));
    CascadeMux I__2487 (
            .O(N__16602),
            .I(N__16599));
    InMux I__2486 (
            .O(N__16599),
            .I(N__16595));
    InMux I__2485 (
            .O(N__16598),
            .I(N__16591));
    LocalMux I__2484 (
            .O(N__16595),
            .I(N__16588));
    InMux I__2483 (
            .O(N__16594),
            .I(N__16584));
    LocalMux I__2482 (
            .O(N__16591),
            .I(N__16581));
    Span4Mux_h I__2481 (
            .O(N__16588),
            .I(N__16578));
    InMux I__2480 (
            .O(N__16587),
            .I(N__16575));
    LocalMux I__2479 (
            .O(N__16584),
            .I(\c0.data_in_field_7 ));
    Odrv4 I__2478 (
            .O(N__16581),
            .I(\c0.data_in_field_7 ));
    Odrv4 I__2477 (
            .O(N__16578),
            .I(\c0.data_in_field_7 ));
    LocalMux I__2476 (
            .O(N__16575),
            .I(\c0.data_in_field_7 ));
    CascadeMux I__2475 (
            .O(N__16566),
            .I(N__16562));
    InMux I__2474 (
            .O(N__16565),
            .I(N__16558));
    InMux I__2473 (
            .O(N__16562),
            .I(N__16555));
    InMux I__2472 (
            .O(N__16561),
            .I(N__16552));
    LocalMux I__2471 (
            .O(N__16558),
            .I(data_in_0_1));
    LocalMux I__2470 (
            .O(N__16555),
            .I(data_in_0_1));
    LocalMux I__2469 (
            .O(N__16552),
            .I(data_in_0_1));
    InMux I__2468 (
            .O(N__16545),
            .I(N__16542));
    LocalMux I__2467 (
            .O(N__16542),
            .I(N__16539));
    Sp12to4 I__2466 (
            .O(N__16539),
            .I(N__16536));
    Odrv12 I__2465 (
            .O(N__16536),
            .I(\c0.n2104 ));
    InMux I__2464 (
            .O(N__16533),
            .I(N__16530));
    LocalMux I__2463 (
            .O(N__16530),
            .I(\c0.n1835 ));
    CascadeMux I__2462 (
            .O(N__16527),
            .I(\c0.n2104_cascade_ ));
    CascadeMux I__2461 (
            .O(N__16524),
            .I(N__16521));
    InMux I__2460 (
            .O(N__16521),
            .I(N__16518));
    LocalMux I__2459 (
            .O(N__16518),
            .I(N__16515));
    Span4Mux_h I__2458 (
            .O(N__16515),
            .I(N__16512));
    Span4Mux_s2_h I__2457 (
            .O(N__16512),
            .I(N__16507));
    InMux I__2456 (
            .O(N__16511),
            .I(N__16502));
    InMux I__2455 (
            .O(N__16510),
            .I(N__16502));
    Odrv4 I__2454 (
            .O(N__16507),
            .I(data_in_8_1));
    LocalMux I__2453 (
            .O(N__16502),
            .I(data_in_8_1));
    InMux I__2452 (
            .O(N__16497),
            .I(N__16494));
    LocalMux I__2451 (
            .O(N__16494),
            .I(N__16491));
    Span4Mux_h I__2450 (
            .O(N__16491),
            .I(N__16485));
    InMux I__2449 (
            .O(N__16490),
            .I(N__16478));
    InMux I__2448 (
            .O(N__16489),
            .I(N__16478));
    InMux I__2447 (
            .O(N__16488),
            .I(N__16478));
    Odrv4 I__2446 (
            .O(N__16485),
            .I(data_in_1_3));
    LocalMux I__2445 (
            .O(N__16478),
            .I(data_in_1_3));
    CascadeMux I__2444 (
            .O(N__16473),
            .I(N__16470));
    InMux I__2443 (
            .O(N__16470),
            .I(N__16466));
    InMux I__2442 (
            .O(N__16469),
            .I(N__16463));
    LocalMux I__2441 (
            .O(N__16466),
            .I(N__16459));
    LocalMux I__2440 (
            .O(N__16463),
            .I(N__16456));
    InMux I__2439 (
            .O(N__16462),
            .I(N__16453));
    Odrv12 I__2438 (
            .O(N__16459),
            .I(data_in_6_3));
    Odrv4 I__2437 (
            .O(N__16456),
            .I(data_in_6_3));
    LocalMux I__2436 (
            .O(N__16453),
            .I(data_in_6_3));
    InMux I__2435 (
            .O(N__16446),
            .I(N__16439));
    InMux I__2434 (
            .O(N__16445),
            .I(N__16439));
    InMux I__2433 (
            .O(N__16444),
            .I(N__16436));
    LocalMux I__2432 (
            .O(N__16439),
            .I(data_in_12_3));
    LocalMux I__2431 (
            .O(N__16436),
            .I(data_in_12_3));
    CascadeMux I__2430 (
            .O(N__16431),
            .I(N__16427));
    InMux I__2429 (
            .O(N__16430),
            .I(N__16423));
    InMux I__2428 (
            .O(N__16427),
            .I(N__16420));
    CascadeMux I__2427 (
            .O(N__16426),
            .I(N__16417));
    LocalMux I__2426 (
            .O(N__16423),
            .I(N__16413));
    LocalMux I__2425 (
            .O(N__16420),
            .I(N__16410));
    InMux I__2424 (
            .O(N__16417),
            .I(N__16407));
    InMux I__2423 (
            .O(N__16416),
            .I(N__16404));
    Span4Mux_s1_h I__2422 (
            .O(N__16413),
            .I(N__16399));
    Span4Mux_v I__2421 (
            .O(N__16410),
            .I(N__16399));
    LocalMux I__2420 (
            .O(N__16407),
            .I(data_in_2_7));
    LocalMux I__2419 (
            .O(N__16404),
            .I(data_in_2_7));
    Odrv4 I__2418 (
            .O(N__16399),
            .I(data_in_2_7));
    InMux I__2417 (
            .O(N__16392),
            .I(N__16388));
    InMux I__2416 (
            .O(N__16391),
            .I(N__16385));
    LocalMux I__2415 (
            .O(N__16388),
            .I(N__16382));
    LocalMux I__2414 (
            .O(N__16385),
            .I(N__16378));
    Span4Mux_h I__2413 (
            .O(N__16382),
            .I(N__16375));
    InMux I__2412 (
            .O(N__16381),
            .I(N__16372));
    Span4Mux_h I__2411 (
            .O(N__16378),
            .I(N__16368));
    Span4Mux_v I__2410 (
            .O(N__16375),
            .I(N__16363));
    LocalMux I__2409 (
            .O(N__16372),
            .I(N__16363));
    InMux I__2408 (
            .O(N__16371),
            .I(N__16358));
    Span4Mux_v I__2407 (
            .O(N__16368),
            .I(N__16355));
    Span4Mux_h I__2406 (
            .O(N__16363),
            .I(N__16352));
    InMux I__2405 (
            .O(N__16362),
            .I(N__16349));
    InMux I__2404 (
            .O(N__16361),
            .I(N__16346));
    LocalMux I__2403 (
            .O(N__16358),
            .I(\c0.data_in_field_131 ));
    Odrv4 I__2402 (
            .O(N__16355),
            .I(\c0.data_in_field_131 ));
    Odrv4 I__2401 (
            .O(N__16352),
            .I(\c0.data_in_field_131 ));
    LocalMux I__2400 (
            .O(N__16349),
            .I(\c0.data_in_field_131 ));
    LocalMux I__2399 (
            .O(N__16346),
            .I(\c0.data_in_field_131 ));
    InMux I__2398 (
            .O(N__16335),
            .I(N__16332));
    LocalMux I__2397 (
            .O(N__16332),
            .I(N__16326));
    InMux I__2396 (
            .O(N__16331),
            .I(N__16323));
    InMux I__2395 (
            .O(N__16330),
            .I(N__16318));
    InMux I__2394 (
            .O(N__16329),
            .I(N__16318));
    Odrv4 I__2393 (
            .O(N__16326),
            .I(data_in_1_1));
    LocalMux I__2392 (
            .O(N__16323),
            .I(data_in_1_1));
    LocalMux I__2391 (
            .O(N__16318),
            .I(data_in_1_1));
    CascadeMux I__2390 (
            .O(N__16311),
            .I(\c0.rx.n6294_cascade_ ));
    InMux I__2389 (
            .O(N__16308),
            .I(N__16298));
    InMux I__2388 (
            .O(N__16307),
            .I(N__16298));
    InMux I__2387 (
            .O(N__16306),
            .I(N__16298));
    InMux I__2386 (
            .O(N__16305),
            .I(N__16290));
    LocalMux I__2385 (
            .O(N__16298),
            .I(N__16287));
    InMux I__2384 (
            .O(N__16297),
            .I(N__16277));
    InMux I__2383 (
            .O(N__16296),
            .I(N__16277));
    InMux I__2382 (
            .O(N__16295),
            .I(N__16277));
    InMux I__2381 (
            .O(N__16294),
            .I(N__16277));
    InMux I__2380 (
            .O(N__16293),
            .I(N__16274));
    LocalMux I__2379 (
            .O(N__16290),
            .I(N__16269));
    Span4Mux_v I__2378 (
            .O(N__16287),
            .I(N__16269));
    InMux I__2377 (
            .O(N__16286),
            .I(N__16266));
    LocalMux I__2376 (
            .O(N__16277),
            .I(N__16263));
    LocalMux I__2375 (
            .O(N__16274),
            .I(N__16260));
    Odrv4 I__2374 (
            .O(N__16269),
            .I(r_SM_Main_2_adj_1989));
    LocalMux I__2373 (
            .O(N__16266),
            .I(r_SM_Main_2_adj_1989));
    Odrv12 I__2372 (
            .O(N__16263),
            .I(r_SM_Main_2_adj_1989));
    Odrv4 I__2371 (
            .O(N__16260),
            .I(r_SM_Main_2_adj_1989));
    CascadeMux I__2370 (
            .O(N__16251),
            .I(\c0.rx.n75_cascade_ ));
    InMux I__2369 (
            .O(N__16248),
            .I(N__16245));
    LocalMux I__2368 (
            .O(N__16245),
            .I(N__16242));
    Odrv12 I__2367 (
            .O(N__16242),
            .I(\c0.rx.n5815 ));
    CascadeMux I__2366 (
            .O(N__16239),
            .I(n4_adj_1980_cascade_));
    InMux I__2365 (
            .O(N__16236),
            .I(N__16230));
    InMux I__2364 (
            .O(N__16235),
            .I(N__16230));
    LocalMux I__2363 (
            .O(N__16230),
            .I(rx_data_4));
    CascadeMux I__2362 (
            .O(N__16227),
            .I(n2198_cascade_));
    InMux I__2361 (
            .O(N__16224),
            .I(N__16219));
    InMux I__2360 (
            .O(N__16223),
            .I(N__16216));
    CascadeMux I__2359 (
            .O(N__16222),
            .I(N__16213));
    LocalMux I__2358 (
            .O(N__16219),
            .I(N__16203));
    LocalMux I__2357 (
            .O(N__16216),
            .I(N__16203));
    InMux I__2356 (
            .O(N__16213),
            .I(N__16194));
    InMux I__2355 (
            .O(N__16212),
            .I(N__16194));
    InMux I__2354 (
            .O(N__16211),
            .I(N__16194));
    InMux I__2353 (
            .O(N__16210),
            .I(N__16194));
    InMux I__2352 (
            .O(N__16209),
            .I(N__16189));
    InMux I__2351 (
            .O(N__16208),
            .I(N__16189));
    Span4Mux_v I__2350 (
            .O(N__16203),
            .I(N__16184));
    LocalMux I__2349 (
            .O(N__16194),
            .I(N__16184));
    LocalMux I__2348 (
            .O(N__16189),
            .I(\c0.rx.n359 ));
    Odrv4 I__2347 (
            .O(N__16184),
            .I(\c0.rx.n359 ));
    InMux I__2346 (
            .O(N__16179),
            .I(N__16176));
    LocalMux I__2345 (
            .O(N__16176),
            .I(\c0.rx.n5859 ));
    InMux I__2344 (
            .O(N__16173),
            .I(N__16168));
    InMux I__2343 (
            .O(N__16172),
            .I(N__16165));
    InMux I__2342 (
            .O(N__16171),
            .I(N__16162));
    LocalMux I__2341 (
            .O(N__16168),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__2340 (
            .O(N__16165),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__2339 (
            .O(N__16162),
            .I(\c0.rx.r_Clock_Count_7 ));
    InMux I__2338 (
            .O(N__16155),
            .I(N__16152));
    LocalMux I__2337 (
            .O(N__16152),
            .I(N__16149));
    Odrv4 I__2336 (
            .O(N__16149),
            .I(\c0.rx.n5823 ));
    CascadeMux I__2335 (
            .O(N__16146),
            .I(N__16142));
    InMux I__2334 (
            .O(N__16145),
            .I(N__16139));
    InMux I__2333 (
            .O(N__16142),
            .I(N__16135));
    LocalMux I__2332 (
            .O(N__16139),
            .I(N__16132));
    InMux I__2331 (
            .O(N__16138),
            .I(N__16128));
    LocalMux I__2330 (
            .O(N__16135),
            .I(N__16125));
    Span4Mux_v I__2329 (
            .O(N__16132),
            .I(N__16122));
    InMux I__2328 (
            .O(N__16131),
            .I(N__16119));
    LocalMux I__2327 (
            .O(N__16128),
            .I(data_in_18_6));
    Odrv4 I__2326 (
            .O(N__16125),
            .I(data_in_18_6));
    Odrv4 I__2325 (
            .O(N__16122),
            .I(data_in_18_6));
    LocalMux I__2324 (
            .O(N__16119),
            .I(data_in_18_6));
    InMux I__2323 (
            .O(N__16110),
            .I(N__16106));
    InMux I__2322 (
            .O(N__16109),
            .I(N__16103));
    LocalMux I__2321 (
            .O(N__16106),
            .I(N__16100));
    LocalMux I__2320 (
            .O(N__16103),
            .I(\c0.data_in_frame_18_6 ));
    Odrv4 I__2319 (
            .O(N__16100),
            .I(\c0.data_in_frame_18_6 ));
    InMux I__2318 (
            .O(N__16095),
            .I(N__16091));
    InMux I__2317 (
            .O(N__16094),
            .I(N__16088));
    LocalMux I__2316 (
            .O(N__16091),
            .I(N__16085));
    LocalMux I__2315 (
            .O(N__16088),
            .I(\c0.data_in_frame_18_7 ));
    Odrv4 I__2314 (
            .O(N__16085),
            .I(\c0.data_in_frame_18_7 ));
    CascadeMux I__2313 (
            .O(N__16080),
            .I(N__16076));
    InMux I__2312 (
            .O(N__16079),
            .I(N__16073));
    InMux I__2311 (
            .O(N__16076),
            .I(N__16070));
    LocalMux I__2310 (
            .O(N__16073),
            .I(N__16067));
    LocalMux I__2309 (
            .O(N__16070),
            .I(N__16063));
    Span12Mux_v I__2308 (
            .O(N__16067),
            .I(N__16060));
    InMux I__2307 (
            .O(N__16066),
            .I(N__16057));
    Odrv4 I__2306 (
            .O(N__16063),
            .I(data_in_7_1));
    Odrv12 I__2305 (
            .O(N__16060),
            .I(data_in_7_1));
    LocalMux I__2304 (
            .O(N__16057),
            .I(data_in_7_1));
    CascadeMux I__2303 (
            .O(N__16050),
            .I(n1764_cascade_));
    InMux I__2302 (
            .O(N__16047),
            .I(N__16044));
    LocalMux I__2301 (
            .O(N__16044),
            .I(N__16040));
    InMux I__2300 (
            .O(N__16043),
            .I(N__16037));
    Odrv4 I__2299 (
            .O(N__16040),
            .I(rx_data_5));
    LocalMux I__2298 (
            .O(N__16037),
            .I(rx_data_5));
    InMux I__2297 (
            .O(N__16032),
            .I(N__16029));
    LocalMux I__2296 (
            .O(N__16029),
            .I(N__16025));
    InMux I__2295 (
            .O(N__16028),
            .I(N__16022));
    Odrv12 I__2294 (
            .O(N__16025),
            .I(rx_data_6));
    LocalMux I__2293 (
            .O(N__16022),
            .I(rx_data_6));
    InMux I__2292 (
            .O(N__16017),
            .I(N__16014));
    LocalMux I__2291 (
            .O(N__16014),
            .I(\c0.rx.n5822 ));
    InMux I__2290 (
            .O(N__16011),
            .I(N__16006));
    InMux I__2289 (
            .O(N__16010),
            .I(N__16003));
    InMux I__2288 (
            .O(N__16009),
            .I(N__16000));
    LocalMux I__2287 (
            .O(N__16006),
            .I(N__15997));
    LocalMux I__2286 (
            .O(N__16003),
            .I(\c0.rx.r_Clock_Count_2 ));
    LocalMux I__2285 (
            .O(N__16000),
            .I(\c0.rx.r_Clock_Count_2 ));
    Odrv4 I__2284 (
            .O(N__15997),
            .I(\c0.rx.r_Clock_Count_2 ));
    InMux I__2283 (
            .O(N__15990),
            .I(N__15987));
    LocalMux I__2282 (
            .O(N__15987),
            .I(n4_adj_1980));
    CascadeMux I__2281 (
            .O(N__15984),
            .I(N__15978));
    InMux I__2280 (
            .O(N__15983),
            .I(N__15975));
    InMux I__2279 (
            .O(N__15982),
            .I(N__15968));
    InMux I__2278 (
            .O(N__15981),
            .I(N__15968));
    InMux I__2277 (
            .O(N__15978),
            .I(N__15968));
    LocalMux I__2276 (
            .O(N__15975),
            .I(data_in_19_6));
    LocalMux I__2275 (
            .O(N__15968),
            .I(data_in_19_6));
    CascadeMux I__2274 (
            .O(N__15963),
            .I(N__15959));
    InMux I__2273 (
            .O(N__15962),
            .I(N__15956));
    InMux I__2272 (
            .O(N__15959),
            .I(N__15953));
    LocalMux I__2271 (
            .O(N__15956),
            .I(N__15950));
    LocalMux I__2270 (
            .O(N__15953),
            .I(\c0.data_in_frame_19_0 ));
    Odrv12 I__2269 (
            .O(N__15950),
            .I(\c0.data_in_frame_19_0 ));
    InMux I__2268 (
            .O(N__15945),
            .I(N__15940));
    InMux I__2267 (
            .O(N__15944),
            .I(N__15935));
    InMux I__2266 (
            .O(N__15943),
            .I(N__15935));
    LocalMux I__2265 (
            .O(N__15940),
            .I(\c0.data_in_field_17 ));
    LocalMux I__2264 (
            .O(N__15935),
            .I(\c0.data_in_field_17 ));
    CascadeMux I__2263 (
            .O(N__15930),
            .I(\c0.n6093_cascade_ ));
    InMux I__2262 (
            .O(N__15927),
            .I(N__15924));
    LocalMux I__2261 (
            .O(N__15924),
            .I(N__15921));
    Span4Mux_h I__2260 (
            .O(N__15921),
            .I(N__15918));
    Odrv4 I__2259 (
            .O(N__15918),
            .I(\c0.n5767 ));
    InMux I__2258 (
            .O(N__15915),
            .I(N__15911));
    InMux I__2257 (
            .O(N__15914),
            .I(N__15908));
    LocalMux I__2256 (
            .O(N__15911),
            .I(N__15902));
    LocalMux I__2255 (
            .O(N__15908),
            .I(N__15902));
    InMux I__2254 (
            .O(N__15907),
            .I(N__15899));
    Odrv12 I__2253 (
            .O(N__15902),
            .I(data_in_16_2));
    LocalMux I__2252 (
            .O(N__15899),
            .I(data_in_16_2));
    InMux I__2251 (
            .O(N__15894),
            .I(N__15891));
    LocalMux I__2250 (
            .O(N__15891),
            .I(N__15888));
    Odrv4 I__2249 (
            .O(N__15888),
            .I(\c0.n5512 ));
    CascadeMux I__2248 (
            .O(N__15885),
            .I(\c0.n5512_cascade_ ));
    InMux I__2247 (
            .O(N__15882),
            .I(N__15879));
    LocalMux I__2246 (
            .O(N__15879),
            .I(\c0.n22 ));
    InMux I__2245 (
            .O(N__15876),
            .I(N__15873));
    LocalMux I__2244 (
            .O(N__15873),
            .I(N__15869));
    InMux I__2243 (
            .O(N__15872),
            .I(N__15866));
    Odrv12 I__2242 (
            .O(N__15869),
            .I(\c0.n2155 ));
    LocalMux I__2241 (
            .O(N__15866),
            .I(\c0.n2155 ));
    CascadeMux I__2240 (
            .O(N__15861),
            .I(\c0.n2155_cascade_ ));
    CascadeMux I__2239 (
            .O(N__15858),
            .I(N__15855));
    InMux I__2238 (
            .O(N__15855),
            .I(N__15852));
    LocalMux I__2237 (
            .O(N__15852),
            .I(N__15849));
    Span4Mux_v I__2236 (
            .O(N__15849),
            .I(N__15846));
    Span4Mux_h I__2235 (
            .O(N__15846),
            .I(N__15843));
    Odrv4 I__2234 (
            .O(N__15843),
            .I(\c0.n43 ));
    InMux I__2233 (
            .O(N__15840),
            .I(N__15837));
    LocalMux I__2232 (
            .O(N__15837),
            .I(N__15834));
    Span4Mux_v I__2231 (
            .O(N__15834),
            .I(N__15830));
    InMux I__2230 (
            .O(N__15833),
            .I(N__15827));
    Odrv4 I__2229 (
            .O(N__15830),
            .I(\c0.n2026 ));
    LocalMux I__2228 (
            .O(N__15827),
            .I(\c0.n2026 ));
    CascadeMux I__2227 (
            .O(N__15822),
            .I(N__15819));
    InMux I__2226 (
            .O(N__15819),
            .I(N__15816));
    LocalMux I__2225 (
            .O(N__15816),
            .I(N__15812));
    InMux I__2224 (
            .O(N__15815),
            .I(N__15809));
    Span4Mux_v I__2223 (
            .O(N__15812),
            .I(N__15805));
    LocalMux I__2222 (
            .O(N__15809),
            .I(N__15802));
    InMux I__2221 (
            .O(N__15808),
            .I(N__15799));
    Odrv4 I__2220 (
            .O(N__15805),
            .I(data_in_16_1));
    Odrv12 I__2219 (
            .O(N__15802),
            .I(data_in_16_1));
    LocalMux I__2218 (
            .O(N__15799),
            .I(data_in_16_1));
    InMux I__2217 (
            .O(N__15792),
            .I(N__15786));
    InMux I__2216 (
            .O(N__15791),
            .I(N__15786));
    LocalMux I__2215 (
            .O(N__15786),
            .I(N__15783));
    Span4Mux_v I__2214 (
            .O(N__15783),
            .I(N__15780));
    Odrv4 I__2213 (
            .O(N__15780),
            .I(\c0.n2080 ));
    InMux I__2212 (
            .O(N__15777),
            .I(N__15774));
    LocalMux I__2211 (
            .O(N__15774),
            .I(N__15770));
    InMux I__2210 (
            .O(N__15773),
            .I(N__15767));
    Odrv4 I__2209 (
            .O(N__15770),
            .I(\c0.n2012 ));
    LocalMux I__2208 (
            .O(N__15767),
            .I(\c0.n2012 ));
    CascadeMux I__2207 (
            .O(N__15762),
            .I(N__15759));
    InMux I__2206 (
            .O(N__15759),
            .I(N__15755));
    InMux I__2205 (
            .O(N__15758),
            .I(N__15752));
    LocalMux I__2204 (
            .O(N__15755),
            .I(\c0.n1973 ));
    LocalMux I__2203 (
            .O(N__15752),
            .I(\c0.n1973 ));
    InMux I__2202 (
            .O(N__15747),
            .I(N__15743));
    InMux I__2201 (
            .O(N__15746),
            .I(N__15740));
    LocalMux I__2200 (
            .O(N__15743),
            .I(N__15737));
    LocalMux I__2199 (
            .O(N__15740),
            .I(N__15730));
    Span4Mux_h I__2198 (
            .O(N__15737),
            .I(N__15730));
    InMux I__2197 (
            .O(N__15736),
            .I(N__15727));
    InMux I__2196 (
            .O(N__15735),
            .I(N__15724));
    Sp12to4 I__2195 (
            .O(N__15730),
            .I(N__15719));
    LocalMux I__2194 (
            .O(N__15727),
            .I(N__15719));
    LocalMux I__2193 (
            .O(N__15724),
            .I(data_in_19_3));
    Odrv12 I__2192 (
            .O(N__15719),
            .I(data_in_19_3));
    CascadeMux I__2191 (
            .O(N__15714),
            .I(\c0.n18_adj_1959_cascade_ ));
    InMux I__2190 (
            .O(N__15711),
            .I(N__15708));
    LocalMux I__2189 (
            .O(N__15708),
            .I(N__15705));
    Odrv4 I__2188 (
            .O(N__15705),
            .I(\c0.n16 ));
    CascadeMux I__2187 (
            .O(N__15702),
            .I(\c0.n20_adj_1870_cascade_ ));
    InMux I__2186 (
            .O(N__15699),
            .I(N__15696));
    LocalMux I__2185 (
            .O(N__15696),
            .I(\c0.n5577 ));
    CascadeMux I__2184 (
            .O(N__15693),
            .I(\c0.n2101_cascade_ ));
    CascadeMux I__2183 (
            .O(N__15690),
            .I(\c0.n6_adj_1917_cascade_ ));
    InMux I__2182 (
            .O(N__15687),
            .I(N__15684));
    LocalMux I__2181 (
            .O(N__15684),
            .I(N__15680));
    InMux I__2180 (
            .O(N__15683),
            .I(N__15677));
    Span4Mux_v I__2179 (
            .O(N__15680),
            .I(N__15672));
    LocalMux I__2178 (
            .O(N__15677),
            .I(N__15669));
    InMux I__2177 (
            .O(N__15676),
            .I(N__15664));
    InMux I__2176 (
            .O(N__15675),
            .I(N__15664));
    Odrv4 I__2175 (
            .O(N__15672),
            .I(\c0.data_in_field_68 ));
    Odrv12 I__2174 (
            .O(N__15669),
            .I(\c0.data_in_field_68 ));
    LocalMux I__2173 (
            .O(N__15664),
            .I(\c0.data_in_field_68 ));
    InMux I__2172 (
            .O(N__15657),
            .I(N__15654));
    LocalMux I__2171 (
            .O(N__15654),
            .I(N__15650));
    InMux I__2170 (
            .O(N__15653),
            .I(N__15647));
    Span4Mux_h I__2169 (
            .O(N__15650),
            .I(N__15644));
    LocalMux I__2168 (
            .O(N__15647),
            .I(\c0.n5557 ));
    Odrv4 I__2167 (
            .O(N__15644),
            .I(\c0.n5557 ));
    CascadeMux I__2166 (
            .O(N__15639),
            .I(\c0.n17_cascade_ ));
    InMux I__2165 (
            .O(N__15636),
            .I(N__15633));
    LocalMux I__2164 (
            .O(N__15633),
            .I(\c0.n5574 ));
    InMux I__2163 (
            .O(N__15630),
            .I(N__15627));
    LocalMux I__2162 (
            .O(N__15627),
            .I(N__15624));
    Span4Mux_v I__2161 (
            .O(N__15624),
            .I(N__15620));
    InMux I__2160 (
            .O(N__15623),
            .I(N__15617));
    Odrv4 I__2159 (
            .O(N__15620),
            .I(\c0.n5572 ));
    LocalMux I__2158 (
            .O(N__15617),
            .I(\c0.n5572 ));
    InMux I__2157 (
            .O(N__15612),
            .I(N__15608));
    InMux I__2156 (
            .O(N__15611),
            .I(N__15605));
    LocalMux I__2155 (
            .O(N__15608),
            .I(N__15602));
    LocalMux I__2154 (
            .O(N__15605),
            .I(N__15599));
    Span4Mux_h I__2153 (
            .O(N__15602),
            .I(N__15595));
    Span4Mux_v I__2152 (
            .O(N__15599),
            .I(N__15592));
    InMux I__2151 (
            .O(N__15598),
            .I(N__15589));
    Odrv4 I__2150 (
            .O(N__15595),
            .I(data_in_8_7));
    Odrv4 I__2149 (
            .O(N__15592),
            .I(data_in_8_7));
    LocalMux I__2148 (
            .O(N__15589),
            .I(data_in_8_7));
    CascadeMux I__2147 (
            .O(N__15582),
            .I(N__15579));
    InMux I__2146 (
            .O(N__15579),
            .I(N__15576));
    LocalMux I__2145 (
            .O(N__15576),
            .I(N__15572));
    InMux I__2144 (
            .O(N__15575),
            .I(N__15569));
    Span4Mux_v I__2143 (
            .O(N__15572),
            .I(N__15565));
    LocalMux I__2142 (
            .O(N__15569),
            .I(N__15562));
    InMux I__2141 (
            .O(N__15568),
            .I(N__15559));
    Odrv4 I__2140 (
            .O(N__15565),
            .I(data_in_17_1));
    Odrv4 I__2139 (
            .O(N__15562),
            .I(data_in_17_1));
    LocalMux I__2138 (
            .O(N__15559),
            .I(data_in_17_1));
    InMux I__2137 (
            .O(N__15552),
            .I(N__15548));
    CascadeMux I__2136 (
            .O(N__15551),
            .I(N__15545));
    LocalMux I__2135 (
            .O(N__15548),
            .I(N__15541));
    InMux I__2134 (
            .O(N__15545),
            .I(N__15536));
    InMux I__2133 (
            .O(N__15544),
            .I(N__15533));
    Span12Mux_v I__2132 (
            .O(N__15541),
            .I(N__15530));
    InMux I__2131 (
            .O(N__15540),
            .I(N__15525));
    InMux I__2130 (
            .O(N__15539),
            .I(N__15525));
    LocalMux I__2129 (
            .O(N__15536),
            .I(\c0.data_in_field_138 ));
    LocalMux I__2128 (
            .O(N__15533),
            .I(\c0.data_in_field_138 ));
    Odrv12 I__2127 (
            .O(N__15530),
            .I(\c0.data_in_field_138 ));
    LocalMux I__2126 (
            .O(N__15525),
            .I(\c0.data_in_field_138 ));
    CascadeMux I__2125 (
            .O(N__15516),
            .I(N__15513));
    InMux I__2124 (
            .O(N__15513),
            .I(N__15509));
    InMux I__2123 (
            .O(N__15512),
            .I(N__15505));
    LocalMux I__2122 (
            .O(N__15509),
            .I(N__15502));
    CascadeMux I__2121 (
            .O(N__15508),
            .I(N__15499));
    LocalMux I__2120 (
            .O(N__15505),
            .I(N__15494));
    Span4Mux_h I__2119 (
            .O(N__15502),
            .I(N__15494));
    InMux I__2118 (
            .O(N__15499),
            .I(N__15489));
    Span4Mux_v I__2117 (
            .O(N__15494),
            .I(N__15486));
    InMux I__2116 (
            .O(N__15493),
            .I(N__15481));
    InMux I__2115 (
            .O(N__15492),
            .I(N__15481));
    LocalMux I__2114 (
            .O(N__15489),
            .I(\c0.data_in_field_130 ));
    Odrv4 I__2113 (
            .O(N__15486),
            .I(\c0.data_in_field_130 ));
    LocalMux I__2112 (
            .O(N__15481),
            .I(\c0.data_in_field_130 ));
    CascadeMux I__2111 (
            .O(N__15474),
            .I(N__15471));
    InMux I__2110 (
            .O(N__15471),
            .I(N__15468));
    LocalMux I__2109 (
            .O(N__15468),
            .I(N__15465));
    Span4Mux_v I__2108 (
            .O(N__15465),
            .I(N__15462));
    Odrv4 I__2107 (
            .O(N__15462),
            .I(\c0.n6213 ));
    InMux I__2106 (
            .O(N__15459),
            .I(N__15454));
    InMux I__2105 (
            .O(N__15458),
            .I(N__15451));
    CascadeMux I__2104 (
            .O(N__15457),
            .I(N__15448));
    LocalMux I__2103 (
            .O(N__15454),
            .I(N__15445));
    LocalMux I__2102 (
            .O(N__15451),
            .I(N__15442));
    InMux I__2101 (
            .O(N__15448),
            .I(N__15437));
    Span4Mux_s3_h I__2100 (
            .O(N__15445),
            .I(N__15434));
    Span4Mux_h I__2099 (
            .O(N__15442),
            .I(N__15431));
    InMux I__2098 (
            .O(N__15441),
            .I(N__15426));
    InMux I__2097 (
            .O(N__15440),
            .I(N__15426));
    LocalMux I__2096 (
            .O(N__15437),
            .I(\c0.data_in_field_73 ));
    Odrv4 I__2095 (
            .O(N__15434),
            .I(\c0.data_in_field_73 ));
    Odrv4 I__2094 (
            .O(N__15431),
            .I(\c0.data_in_field_73 ));
    LocalMux I__2093 (
            .O(N__15426),
            .I(\c0.data_in_field_73 ));
    CascadeMux I__2092 (
            .O(N__15417),
            .I(\c0.n14_adj_1957_cascade_ ));
    InMux I__2091 (
            .O(N__15414),
            .I(N__15406));
    InMux I__2090 (
            .O(N__15413),
            .I(N__15406));
    InMux I__2089 (
            .O(N__15412),
            .I(N__15401));
    InMux I__2088 (
            .O(N__15411),
            .I(N__15401));
    LocalMux I__2087 (
            .O(N__15406),
            .I(\c0.data_in_field_53 ));
    LocalMux I__2086 (
            .O(N__15401),
            .I(\c0.data_in_field_53 ));
    CascadeMux I__2085 (
            .O(N__15396),
            .I(\c0.n22_adj_1903_cascade_ ));
    InMux I__2084 (
            .O(N__15393),
            .I(N__15390));
    LocalMux I__2083 (
            .O(N__15390),
            .I(\c0.n18_adj_1904 ));
    InMux I__2082 (
            .O(N__15387),
            .I(N__15384));
    LocalMux I__2081 (
            .O(N__15384),
            .I(\c0.n20_adj_1905 ));
    CascadeMux I__2080 (
            .O(N__15381),
            .I(\c0.n5589_cascade_ ));
    CascadeMux I__2079 (
            .O(N__15378),
            .I(N__15375));
    InMux I__2078 (
            .O(N__15375),
            .I(N__15372));
    LocalMux I__2077 (
            .O(N__15372),
            .I(N__15369));
    Span4Mux_h I__2076 (
            .O(N__15369),
            .I(N__15366));
    Span4Mux_v I__2075 (
            .O(N__15366),
            .I(N__15363));
    Odrv4 I__2074 (
            .O(N__15363),
            .I(\c0.n29 ));
    InMux I__2073 (
            .O(N__15360),
            .I(N__15354));
    InMux I__2072 (
            .O(N__15359),
            .I(N__15354));
    LocalMux I__2071 (
            .O(N__15354),
            .I(\c0.n5458 ));
    CascadeMux I__2070 (
            .O(N__15351),
            .I(N__15348));
    InMux I__2069 (
            .O(N__15348),
            .I(N__15345));
    LocalMux I__2068 (
            .O(N__15345),
            .I(N__15342));
    Span4Mux_h I__2067 (
            .O(N__15342),
            .I(N__15338));
    InMux I__2066 (
            .O(N__15341),
            .I(N__15335));
    Odrv4 I__2065 (
            .O(N__15338),
            .I(\c0.n1994 ));
    LocalMux I__2064 (
            .O(N__15335),
            .I(\c0.n1994 ));
    CascadeMux I__2063 (
            .O(N__15330),
            .I(\c0.n6009_cascade_ ));
    InMux I__2062 (
            .O(N__15327),
            .I(N__15324));
    LocalMux I__2061 (
            .O(N__15324),
            .I(N__15321));
    Span4Mux_v I__2060 (
            .O(N__15321),
            .I(N__15318));
    Odrv4 I__2059 (
            .O(N__15318),
            .I(\c0.n6012 ));
    InMux I__2058 (
            .O(N__15315),
            .I(N__15310));
    InMux I__2057 (
            .O(N__15314),
            .I(N__15305));
    InMux I__2056 (
            .O(N__15313),
            .I(N__15305));
    LocalMux I__2055 (
            .O(N__15310),
            .I(\c0.data_in_field_15 ));
    LocalMux I__2054 (
            .O(N__15305),
            .I(\c0.data_in_field_15 ));
    InMux I__2053 (
            .O(N__15300),
            .I(N__15297));
    LocalMux I__2052 (
            .O(N__15297),
            .I(N__15294));
    Span4Mux_s2_h I__2051 (
            .O(N__15294),
            .I(N__15291));
    Span4Mux_v I__2050 (
            .O(N__15291),
            .I(N__15286));
    InMux I__2049 (
            .O(N__15290),
            .I(N__15281));
    InMux I__2048 (
            .O(N__15289),
            .I(N__15281));
    Odrv4 I__2047 (
            .O(N__15286),
            .I(\c0.data_in_field_8 ));
    LocalMux I__2046 (
            .O(N__15281),
            .I(\c0.data_in_field_8 ));
    InMux I__2045 (
            .O(N__15276),
            .I(N__15273));
    LocalMux I__2044 (
            .O(N__15273),
            .I(\c0.n2039 ));
    CascadeMux I__2043 (
            .O(N__15270),
            .I(\c0.n2039_cascade_ ));
    InMux I__2042 (
            .O(N__15267),
            .I(N__15262));
    InMux I__2041 (
            .O(N__15266),
            .I(N__15258));
    InMux I__2040 (
            .O(N__15265),
            .I(N__15255));
    LocalMux I__2039 (
            .O(N__15262),
            .I(N__15252));
    InMux I__2038 (
            .O(N__15261),
            .I(N__15249));
    LocalMux I__2037 (
            .O(N__15258),
            .I(\c0.data_in_field_23 ));
    LocalMux I__2036 (
            .O(N__15255),
            .I(\c0.data_in_field_23 ));
    Odrv4 I__2035 (
            .O(N__15252),
            .I(\c0.data_in_field_23 ));
    LocalMux I__2034 (
            .O(N__15249),
            .I(\c0.data_in_field_23 ));
    InMux I__2033 (
            .O(N__15240),
            .I(N__15237));
    LocalMux I__2032 (
            .O(N__15237),
            .I(\c0.rx.n5857 ));
    CascadeMux I__2031 (
            .O(N__15234),
            .I(N__15230));
    InMux I__2030 (
            .O(N__15233),
            .I(N__15226));
    InMux I__2029 (
            .O(N__15230),
            .I(N__15223));
    InMux I__2028 (
            .O(N__15229),
            .I(N__15220));
    LocalMux I__2027 (
            .O(N__15226),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__2026 (
            .O(N__15223),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__2025 (
            .O(N__15220),
            .I(\c0.rx.r_Clock_Count_4 ));
    IoInMux I__2024 (
            .O(N__15213),
            .I(N__15210));
    LocalMux I__2023 (
            .O(N__15210),
            .I(tx_enable));
    CascadeMux I__2022 (
            .O(N__15207),
            .I(N__15204));
    InMux I__2021 (
            .O(N__15204),
            .I(N__15201));
    LocalMux I__2020 (
            .O(N__15201),
            .I(N__15197));
    InMux I__2019 (
            .O(N__15200),
            .I(N__15194));
    Span4Mux_v I__2018 (
            .O(N__15197),
            .I(N__15190));
    LocalMux I__2017 (
            .O(N__15194),
            .I(N__15187));
    InMux I__2016 (
            .O(N__15193),
            .I(N__15184));
    Odrv4 I__2015 (
            .O(N__15190),
            .I(data_in_16_3));
    Odrv4 I__2014 (
            .O(N__15187),
            .I(data_in_16_3));
    LocalMux I__2013 (
            .O(N__15184),
            .I(data_in_16_3));
    CascadeMux I__2012 (
            .O(N__15177),
            .I(N__15174));
    InMux I__2011 (
            .O(N__15174),
            .I(N__15168));
    InMux I__2010 (
            .O(N__15173),
            .I(N__15168));
    LocalMux I__2009 (
            .O(N__15168),
            .I(rx_data_3));
    CascadeMux I__2008 (
            .O(N__15165),
            .I(N__15162));
    InMux I__2007 (
            .O(N__15162),
            .I(N__15158));
    InMux I__2006 (
            .O(N__15161),
            .I(N__15155));
    LocalMux I__2005 (
            .O(N__15158),
            .I(N__15152));
    LocalMux I__2004 (
            .O(N__15155),
            .I(N__15149));
    Span4Mux_v I__2003 (
            .O(N__15152),
            .I(N__15144));
    Span4Mux_v I__2002 (
            .O(N__15149),
            .I(N__15141));
    InMux I__2001 (
            .O(N__15148),
            .I(N__15138));
    InMux I__2000 (
            .O(N__15147),
            .I(N__15135));
    Span4Mux_v I__1999 (
            .O(N__15144),
            .I(N__15132));
    Odrv4 I__1998 (
            .O(N__15141),
            .I(data_in_18_1));
    LocalMux I__1997 (
            .O(N__15138),
            .I(data_in_18_1));
    LocalMux I__1996 (
            .O(N__15135),
            .I(data_in_18_1));
    Odrv4 I__1995 (
            .O(N__15132),
            .I(data_in_18_1));
    InMux I__1994 (
            .O(N__15123),
            .I(N__15111));
    InMux I__1993 (
            .O(N__15122),
            .I(N__15111));
    InMux I__1992 (
            .O(N__15121),
            .I(N__15111));
    InMux I__1991 (
            .O(N__15120),
            .I(N__15111));
    LocalMux I__1990 (
            .O(N__15111),
            .I(N__15104));
    InMux I__1989 (
            .O(N__15110),
            .I(N__15095));
    InMux I__1988 (
            .O(N__15109),
            .I(N__15095));
    InMux I__1987 (
            .O(N__15108),
            .I(N__15095));
    InMux I__1986 (
            .O(N__15107),
            .I(N__15095));
    Odrv4 I__1985 (
            .O(N__15104),
            .I(\c0.rx.n36 ));
    LocalMux I__1984 (
            .O(N__15095),
            .I(\c0.rx.n36 ));
    InMux I__1983 (
            .O(N__15090),
            .I(\c0.rx.n4778 ));
    InMux I__1982 (
            .O(N__15087),
            .I(N__15084));
    LocalMux I__1981 (
            .O(N__15084),
            .I(\c0.rx.n5361 ));
    InMux I__1980 (
            .O(N__15081),
            .I(N__15078));
    LocalMux I__1979 (
            .O(N__15078),
            .I(\c0.rx.n5858 ));
    InMux I__1978 (
            .O(N__15075),
            .I(N__15072));
    LocalMux I__1977 (
            .O(N__15072),
            .I(\c0.rx.n5854 ));
    InMux I__1976 (
            .O(N__15069),
            .I(N__15064));
    InMux I__1975 (
            .O(N__15068),
            .I(N__15061));
    InMux I__1974 (
            .O(N__15067),
            .I(N__15058));
    LocalMux I__1973 (
            .O(N__15064),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__1972 (
            .O(N__15061),
            .I(\c0.rx.r_Clock_Count_3 ));
    LocalMux I__1971 (
            .O(N__15058),
            .I(\c0.rx.r_Clock_Count_3 ));
    InMux I__1970 (
            .O(N__15051),
            .I(N__15046));
    InMux I__1969 (
            .O(N__15050),
            .I(N__15041));
    InMux I__1968 (
            .O(N__15049),
            .I(N__15041));
    LocalMux I__1967 (
            .O(N__15046),
            .I(\c0.rx.r_Clock_Count_6 ));
    LocalMux I__1966 (
            .O(N__15041),
            .I(\c0.rx.r_Clock_Count_6 ));
    InMux I__1965 (
            .O(N__15036),
            .I(N__15031));
    InMux I__1964 (
            .O(N__15035),
            .I(N__15028));
    InMux I__1963 (
            .O(N__15034),
            .I(N__15025));
    LocalMux I__1962 (
            .O(N__15031),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__1961 (
            .O(N__15028),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__1960 (
            .O(N__15025),
            .I(\c0.rx.r_Clock_Count_5 ));
    CascadeMux I__1959 (
            .O(N__15018),
            .I(\c0.rx.n8_cascade_ ));
    InMux I__1958 (
            .O(N__15015),
            .I(N__15003));
    InMux I__1957 (
            .O(N__15014),
            .I(N__15003));
    InMux I__1956 (
            .O(N__15013),
            .I(N__15003));
    InMux I__1955 (
            .O(N__15012),
            .I(N__15003));
    LocalMux I__1954 (
            .O(N__15003),
            .I(\c0.rx.n1724 ));
    CascadeMux I__1953 (
            .O(N__15000),
            .I(\c0.rx.n1724_cascade_ ));
    InMux I__1952 (
            .O(N__14997),
            .I(N__14988));
    InMux I__1951 (
            .O(N__14996),
            .I(N__14985));
    InMux I__1950 (
            .O(N__14995),
            .I(N__14982));
    InMux I__1949 (
            .O(N__14994),
            .I(N__14975));
    InMux I__1948 (
            .O(N__14993),
            .I(N__14975));
    InMux I__1947 (
            .O(N__14992),
            .I(N__14975));
    InMux I__1946 (
            .O(N__14991),
            .I(N__14972));
    LocalMux I__1945 (
            .O(N__14988),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__1944 (
            .O(N__14985),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__1943 (
            .O(N__14982),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__1942 (
            .O(N__14975),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__1941 (
            .O(N__14972),
            .I(\c0.rx.r_Clock_Count_1 ));
    InMux I__1940 (
            .O(N__14961),
            .I(N__14958));
    LocalMux I__1939 (
            .O(N__14958),
            .I(\c0.rx.n5855 ));
    InMux I__1938 (
            .O(N__14955),
            .I(N__14946));
    InMux I__1937 (
            .O(N__14954),
            .I(N__14943));
    InMux I__1936 (
            .O(N__14953),
            .I(N__14938));
    InMux I__1935 (
            .O(N__14952),
            .I(N__14938));
    InMux I__1934 (
            .O(N__14951),
            .I(N__14931));
    InMux I__1933 (
            .O(N__14950),
            .I(N__14931));
    InMux I__1932 (
            .O(N__14949),
            .I(N__14931));
    LocalMux I__1931 (
            .O(N__14946),
            .I(\c0.rx.r_Clock_Count_0 ));
    LocalMux I__1930 (
            .O(N__14943),
            .I(\c0.rx.r_Clock_Count_0 ));
    LocalMux I__1929 (
            .O(N__14938),
            .I(\c0.rx.r_Clock_Count_0 ));
    LocalMux I__1928 (
            .O(N__14931),
            .I(\c0.rx.r_Clock_Count_0 ));
    CascadeMux I__1927 (
            .O(N__14922),
            .I(N__14918));
    InMux I__1926 (
            .O(N__14921),
            .I(N__14915));
    InMux I__1925 (
            .O(N__14918),
            .I(N__14911));
    LocalMux I__1924 (
            .O(N__14915),
            .I(N__14908));
    InMux I__1923 (
            .O(N__14914),
            .I(N__14905));
    LocalMux I__1922 (
            .O(N__14911),
            .I(\c0.data_in_field_104 ));
    Odrv12 I__1921 (
            .O(N__14908),
            .I(\c0.data_in_field_104 ));
    LocalMux I__1920 (
            .O(N__14905),
            .I(\c0.data_in_field_104 ));
    CascadeMux I__1919 (
            .O(N__14898),
            .I(\c0.n6021_cascade_ ));
    InMux I__1918 (
            .O(N__14895),
            .I(N__14892));
    LocalMux I__1917 (
            .O(N__14892),
            .I(N__14889));
    Span4Mux_s3_h I__1916 (
            .O(N__14889),
            .I(N__14886));
    Odrv4 I__1915 (
            .O(N__14886),
            .I(\c0.n5797 ));
    InMux I__1914 (
            .O(N__14883),
            .I(bfn_4_27_0_));
    InMux I__1913 (
            .O(N__14880),
            .I(N__14877));
    LocalMux I__1912 (
            .O(N__14877),
            .I(\c0.rx.n5860 ));
    InMux I__1911 (
            .O(N__14874),
            .I(\c0.rx.n4772 ));
    InMux I__1910 (
            .O(N__14871),
            .I(\c0.rx.n4773 ));
    InMux I__1909 (
            .O(N__14868),
            .I(N__14865));
    LocalMux I__1908 (
            .O(N__14865),
            .I(\c0.rx.n5856 ));
    InMux I__1907 (
            .O(N__14862),
            .I(\c0.rx.n4774 ));
    InMux I__1906 (
            .O(N__14859),
            .I(\c0.rx.n4775 ));
    InMux I__1905 (
            .O(N__14856),
            .I(\c0.rx.n4776 ));
    InMux I__1904 (
            .O(N__14853),
            .I(\c0.rx.n4777 ));
    CascadeMux I__1903 (
            .O(N__14850),
            .I(\c0.n6147_cascade_ ));
    InMux I__1902 (
            .O(N__14847),
            .I(N__14844));
    LocalMux I__1901 (
            .O(N__14844),
            .I(N__14841));
    Span4Mux_v I__1900 (
            .O(N__14841),
            .I(N__14838));
    IoSpan4Mux I__1899 (
            .O(N__14838),
            .I(N__14835));
    Span4Mux_s1_h I__1898 (
            .O(N__14835),
            .I(N__14832));
    Odrv4 I__1897 (
            .O(N__14832),
            .I(\c0.n6150 ));
    InMux I__1896 (
            .O(N__14829),
            .I(N__14825));
    InMux I__1895 (
            .O(N__14828),
            .I(N__14822));
    LocalMux I__1894 (
            .O(N__14825),
            .I(N__14819));
    LocalMux I__1893 (
            .O(N__14822),
            .I(\c0.data_in_frame_19_4 ));
    Odrv4 I__1892 (
            .O(N__14819),
            .I(\c0.data_in_frame_19_4 ));
    InMux I__1891 (
            .O(N__14814),
            .I(N__14811));
    LocalMux I__1890 (
            .O(N__14811),
            .I(N__14808));
    Span4Mux_v I__1889 (
            .O(N__14808),
            .I(N__14803));
    InMux I__1888 (
            .O(N__14807),
            .I(N__14798));
    InMux I__1887 (
            .O(N__14806),
            .I(N__14798));
    Odrv4 I__1886 (
            .O(N__14803),
            .I(\c0.data_in_field_14 ));
    LocalMux I__1885 (
            .O(N__14798),
            .I(\c0.data_in_field_14 ));
    CascadeMux I__1884 (
            .O(N__14793),
            .I(\c0.n6255_cascade_ ));
    CascadeMux I__1883 (
            .O(N__14790),
            .I(N__14787));
    InMux I__1882 (
            .O(N__14787),
            .I(N__14784));
    LocalMux I__1881 (
            .O(N__14784),
            .I(\c0.n5692 ));
    InMux I__1880 (
            .O(N__14781),
            .I(N__14778));
    LocalMux I__1879 (
            .O(N__14778),
            .I(N__14775));
    Span4Mux_v I__1878 (
            .O(N__14775),
            .I(N__14770));
    InMux I__1877 (
            .O(N__14774),
            .I(N__14765));
    InMux I__1876 (
            .O(N__14773),
            .I(N__14765));
    Odrv4 I__1875 (
            .O(N__14770),
            .I(\c0.data_in_field_119 ));
    LocalMux I__1874 (
            .O(N__14765),
            .I(\c0.data_in_field_119 ));
    CascadeMux I__1873 (
            .O(N__14760),
            .I(\c0.n6273_cascade_ ));
    InMux I__1872 (
            .O(N__14757),
            .I(N__14754));
    LocalMux I__1871 (
            .O(N__14754),
            .I(N__14750));
    InMux I__1870 (
            .O(N__14753),
            .I(N__14746));
    Span4Mux_v I__1869 (
            .O(N__14750),
            .I(N__14743));
    InMux I__1868 (
            .O(N__14749),
            .I(N__14740));
    LocalMux I__1867 (
            .O(N__14746),
            .I(\c0.data_in_field_111 ));
    Odrv4 I__1866 (
            .O(N__14743),
            .I(\c0.data_in_field_111 ));
    LocalMux I__1865 (
            .O(N__14740),
            .I(\c0.data_in_field_111 ));
    InMux I__1864 (
            .O(N__14733),
            .I(N__14730));
    LocalMux I__1863 (
            .O(N__14730),
            .I(\c0.n5994 ));
    CascadeMux I__1862 (
            .O(N__14727),
            .I(\c0.n5686_cascade_ ));
    CascadeMux I__1861 (
            .O(N__14724),
            .I(\c0.n6261_cascade_ ));
    InMux I__1860 (
            .O(N__14721),
            .I(N__14718));
    LocalMux I__1859 (
            .O(N__14718),
            .I(\c0.n6264 ));
    InMux I__1858 (
            .O(N__14715),
            .I(N__14710));
    InMux I__1857 (
            .O(N__14714),
            .I(N__14707));
    CascadeMux I__1856 (
            .O(N__14713),
            .I(N__14704));
    LocalMux I__1855 (
            .O(N__14710),
            .I(N__14701));
    LocalMux I__1854 (
            .O(N__14707),
            .I(N__14698));
    InMux I__1853 (
            .O(N__14704),
            .I(N__14695));
    Span4Mux_s3_h I__1852 (
            .O(N__14701),
            .I(N__14691));
    Span4Mux_h I__1851 (
            .O(N__14698),
            .I(N__14688));
    LocalMux I__1850 (
            .O(N__14695),
            .I(N__14685));
    InMux I__1849 (
            .O(N__14694),
            .I(N__14682));
    Sp12to4 I__1848 (
            .O(N__14691),
            .I(N__14679));
    Span4Mux_v I__1847 (
            .O(N__14688),
            .I(N__14674));
    Span4Mux_h I__1846 (
            .O(N__14685),
            .I(N__14674));
    LocalMux I__1845 (
            .O(N__14682),
            .I(data_in_18_3));
    Odrv12 I__1844 (
            .O(N__14679),
            .I(data_in_18_3));
    Odrv4 I__1843 (
            .O(N__14674),
            .I(data_in_18_3));
    InMux I__1842 (
            .O(N__14667),
            .I(N__14664));
    LocalMux I__1841 (
            .O(N__14664),
            .I(N__14661));
    Odrv12 I__1840 (
            .O(N__14661),
            .I(\c0.n5725 ));
    InMux I__1839 (
            .O(N__14658),
            .I(N__14655));
    LocalMux I__1838 (
            .O(N__14655),
            .I(N__14652));
    Odrv4 I__1837 (
            .O(N__14652),
            .I(\c0.n6165 ));
    InMux I__1836 (
            .O(N__14649),
            .I(N__14646));
    LocalMux I__1835 (
            .O(N__14646),
            .I(N__14643));
    Span4Mux_v I__1834 (
            .O(N__14643),
            .I(N__14640));
    Odrv4 I__1833 (
            .O(N__14640),
            .I(\c0.n6168 ));
    CascadeMux I__1832 (
            .O(N__14637),
            .I(N__14634));
    InMux I__1831 (
            .O(N__14634),
            .I(N__14631));
    LocalMux I__1830 (
            .O(N__14631),
            .I(\c0.n20_adj_1878 ));
    CascadeMux I__1829 (
            .O(N__14628),
            .I(N__14625));
    InMux I__1828 (
            .O(N__14625),
            .I(N__14622));
    LocalMux I__1827 (
            .O(N__14622),
            .I(N__14618));
    InMux I__1826 (
            .O(N__14621),
            .I(N__14615));
    Span12Mux_s11_v I__1825 (
            .O(N__14618),
            .I(N__14611));
    LocalMux I__1824 (
            .O(N__14615),
            .I(N__14608));
    InMux I__1823 (
            .O(N__14614),
            .I(N__14605));
    Odrv12 I__1822 (
            .O(N__14611),
            .I(data_in_7_2));
    Odrv4 I__1821 (
            .O(N__14608),
            .I(data_in_7_2));
    LocalMux I__1820 (
            .O(N__14605),
            .I(data_in_7_2));
    InMux I__1819 (
            .O(N__14598),
            .I(N__14595));
    LocalMux I__1818 (
            .O(N__14595),
            .I(N__14591));
    CascadeMux I__1817 (
            .O(N__14594),
            .I(N__14587));
    Span4Mux_v I__1816 (
            .O(N__14591),
            .I(N__14583));
    InMux I__1815 (
            .O(N__14590),
            .I(N__14576));
    InMux I__1814 (
            .O(N__14587),
            .I(N__14576));
    InMux I__1813 (
            .O(N__14586),
            .I(N__14576));
    Odrv4 I__1812 (
            .O(N__14583),
            .I(\c0.data_in_field_58 ));
    LocalMux I__1811 (
            .O(N__14576),
            .I(\c0.data_in_field_58 ));
    CascadeMux I__1810 (
            .O(N__14571),
            .I(N__14567));
    InMux I__1809 (
            .O(N__14570),
            .I(N__14564));
    InMux I__1808 (
            .O(N__14567),
            .I(N__14561));
    LocalMux I__1807 (
            .O(N__14564),
            .I(\c0.data_in_frame_19_6 ));
    LocalMux I__1806 (
            .O(N__14561),
            .I(\c0.data_in_frame_19_6 ));
    InMux I__1805 (
            .O(N__14556),
            .I(N__14553));
    LocalMux I__1804 (
            .O(N__14553),
            .I(N__14550));
    Odrv4 I__1803 (
            .O(N__14550),
            .I(\c0.n5578 ));
    CascadeMux I__1802 (
            .O(N__14547),
            .I(\c0.n6177_cascade_ ));
    CascadeMux I__1801 (
            .O(N__14544),
            .I(\c0.n5728_cascade_ ));
    CascadeMux I__1800 (
            .O(N__14541),
            .I(\c0.n16_adj_1873_cascade_ ));
    InMux I__1799 (
            .O(N__14538),
            .I(N__14535));
    LocalMux I__1798 (
            .O(N__14535),
            .I(\c0.n24 ));
    InMux I__1797 (
            .O(N__14532),
            .I(N__14526));
    InMux I__1796 (
            .O(N__14531),
            .I(N__14521));
    InMux I__1795 (
            .O(N__14530),
            .I(N__14521));
    InMux I__1794 (
            .O(N__14529),
            .I(N__14518));
    LocalMux I__1793 (
            .O(N__14526),
            .I(\c0.data_in_field_81 ));
    LocalMux I__1792 (
            .O(N__14521),
            .I(\c0.data_in_field_81 ));
    LocalMux I__1791 (
            .O(N__14518),
            .I(\c0.data_in_field_81 ));
    CascadeMux I__1790 (
            .O(N__14511),
            .I(N__14508));
    InMux I__1789 (
            .O(N__14508),
            .I(N__14505));
    LocalMux I__1788 (
            .O(N__14505),
            .I(N__14502));
    Span4Mux_v I__1787 (
            .O(N__14502),
            .I(N__14499));
    Odrv4 I__1786 (
            .O(N__14499),
            .I(\c0.n5551 ));
    CascadeMux I__1785 (
            .O(N__14496),
            .I(\c0.n5551_cascade_ ));
    InMux I__1784 (
            .O(N__14493),
            .I(N__14490));
    LocalMux I__1783 (
            .O(N__14490),
            .I(N__14487));
    Span4Mux_h I__1782 (
            .O(N__14487),
            .I(N__14483));
    InMux I__1781 (
            .O(N__14486),
            .I(N__14480));
    Odrv4 I__1780 (
            .O(N__14483),
            .I(\c0.n1892 ));
    LocalMux I__1779 (
            .O(N__14480),
            .I(\c0.n1892 ));
    InMux I__1778 (
            .O(N__14475),
            .I(N__14472));
    LocalMux I__1777 (
            .O(N__14472),
            .I(\c0.n20 ));
    CascadeMux I__1776 (
            .O(N__14469),
            .I(\c0.n19_cascade_ ));
    InMux I__1775 (
            .O(N__14466),
            .I(N__14461));
    InMux I__1774 (
            .O(N__14465),
            .I(N__14458));
    InMux I__1773 (
            .O(N__14464),
            .I(N__14455));
    LocalMux I__1772 (
            .O(N__14461),
            .I(data_in_10_3));
    LocalMux I__1771 (
            .O(N__14458),
            .I(data_in_10_3));
    LocalMux I__1770 (
            .O(N__14455),
            .I(data_in_10_3));
    CascadeMux I__1769 (
            .O(N__14448),
            .I(\c0.n5412_cascade_ ));
    InMux I__1768 (
            .O(N__14445),
            .I(N__14442));
    LocalMux I__1767 (
            .O(N__14442),
            .I(N__14439));
    Odrv4 I__1766 (
            .O(N__14439),
            .I(\c0.n16_adj_1880 ));
    CascadeMux I__1765 (
            .O(N__14436),
            .I(\c0.n22_adj_1881_cascade_ ));
    InMux I__1764 (
            .O(N__14433),
            .I(N__14430));
    LocalMux I__1763 (
            .O(N__14430),
            .I(N__14427));
    Span4Mux_s3_h I__1762 (
            .O(N__14427),
            .I(N__14424));
    Sp12to4 I__1761 (
            .O(N__14424),
            .I(N__14421));
    Odrv12 I__1760 (
            .O(N__14421),
            .I(\c0.n24_adj_1884 ));
    InMux I__1759 (
            .O(N__14418),
            .I(N__14415));
    LocalMux I__1758 (
            .O(N__14415),
            .I(N__14411));
    InMux I__1757 (
            .O(N__14414),
            .I(N__14406));
    Span4Mux_v I__1756 (
            .O(N__14411),
            .I(N__14403));
    InMux I__1755 (
            .O(N__14410),
            .I(N__14398));
    InMux I__1754 (
            .O(N__14409),
            .I(N__14398));
    LocalMux I__1753 (
            .O(N__14406),
            .I(\c0.data_in_field_11 ));
    Odrv4 I__1752 (
            .O(N__14403),
            .I(\c0.data_in_field_11 ));
    LocalMux I__1751 (
            .O(N__14398),
            .I(\c0.data_in_field_11 ));
    CascadeMux I__1750 (
            .O(N__14391),
            .I(N__14387));
    InMux I__1749 (
            .O(N__14390),
            .I(N__14384));
    InMux I__1748 (
            .O(N__14387),
            .I(N__14380));
    LocalMux I__1747 (
            .O(N__14384),
            .I(N__14377));
    InMux I__1746 (
            .O(N__14383),
            .I(N__14374));
    LocalMux I__1745 (
            .O(N__14380),
            .I(data_in_8_3));
    Odrv4 I__1744 (
            .O(N__14377),
            .I(data_in_8_3));
    LocalMux I__1743 (
            .O(N__14374),
            .I(data_in_8_3));
    CascadeMux I__1742 (
            .O(N__14367),
            .I(N__14361));
    InMux I__1741 (
            .O(N__14366),
            .I(N__14358));
    InMux I__1740 (
            .O(N__14365),
            .I(N__14355));
    InMux I__1739 (
            .O(N__14364),
            .I(N__14352));
    InMux I__1738 (
            .O(N__14361),
            .I(N__14349));
    LocalMux I__1737 (
            .O(N__14358),
            .I(\c0.data_in_field_67 ));
    LocalMux I__1736 (
            .O(N__14355),
            .I(\c0.data_in_field_67 ));
    LocalMux I__1735 (
            .O(N__14352),
            .I(\c0.data_in_field_67 ));
    LocalMux I__1734 (
            .O(N__14349),
            .I(\c0.data_in_field_67 ));
    CascadeMux I__1733 (
            .O(N__14340),
            .I(\c0.rx.n3589_cascade_ ));
    CascadeMux I__1732 (
            .O(N__14337),
            .I(\c0.rx.n17_cascade_ ));
    InMux I__1731 (
            .O(N__14334),
            .I(N__14331));
    LocalMux I__1730 (
            .O(N__14331),
            .I(\c0.rx.n5817 ));
    CascadeMux I__1729 (
            .O(N__14328),
            .I(N__14325));
    InMux I__1728 (
            .O(N__14325),
            .I(N__14322));
    LocalMux I__1727 (
            .O(N__14322),
            .I(N__14317));
    InMux I__1726 (
            .O(N__14321),
            .I(N__14314));
    InMux I__1725 (
            .O(N__14320),
            .I(N__14311));
    Span4Mux_h I__1724 (
            .O(N__14317),
            .I(N__14308));
    LocalMux I__1723 (
            .O(N__14314),
            .I(data_in_15_3));
    LocalMux I__1722 (
            .O(N__14311),
            .I(data_in_15_3));
    Odrv4 I__1721 (
            .O(N__14308),
            .I(data_in_15_3));
    InMux I__1720 (
            .O(N__14301),
            .I(N__14298));
    LocalMux I__1719 (
            .O(N__14298),
            .I(N__14294));
    InMux I__1718 (
            .O(N__14297),
            .I(N__14290));
    Span4Mux_v I__1717 (
            .O(N__14294),
            .I(N__14287));
    InMux I__1716 (
            .O(N__14293),
            .I(N__14284));
    LocalMux I__1715 (
            .O(N__14290),
            .I(\c0.data_in_field_59 ));
    Odrv4 I__1714 (
            .O(N__14287),
            .I(\c0.data_in_field_59 ));
    LocalMux I__1713 (
            .O(N__14284),
            .I(\c0.data_in_field_59 ));
    InMux I__1712 (
            .O(N__14277),
            .I(N__14274));
    LocalMux I__1711 (
            .O(N__14274),
            .I(N__14268));
    InMux I__1710 (
            .O(N__14273),
            .I(N__14263));
    InMux I__1709 (
            .O(N__14272),
            .I(N__14263));
    InMux I__1708 (
            .O(N__14271),
            .I(N__14260));
    Span4Mux_s3_h I__1707 (
            .O(N__14268),
            .I(N__14257));
    LocalMux I__1706 (
            .O(N__14263),
            .I(N__14254));
    LocalMux I__1705 (
            .O(N__14260),
            .I(\c0.data_in_field_123 ));
    Odrv4 I__1704 (
            .O(N__14257),
            .I(\c0.data_in_field_123 ));
    Odrv4 I__1703 (
            .O(N__14254),
            .I(\c0.data_in_field_123 ));
    CascadeMux I__1702 (
            .O(N__14247),
            .I(N__14243));
    InMux I__1701 (
            .O(N__14246),
            .I(N__14239));
    InMux I__1700 (
            .O(N__14243),
            .I(N__14234));
    InMux I__1699 (
            .O(N__14242),
            .I(N__14234));
    LocalMux I__1698 (
            .O(N__14239),
            .I(data_in_7_3));
    LocalMux I__1697 (
            .O(N__14234),
            .I(data_in_7_3));
    InMux I__1696 (
            .O(N__14229),
            .I(\c0.n4738 ));
    InMux I__1695 (
            .O(N__14226),
            .I(N__14222));
    InMux I__1694 (
            .O(N__14225),
            .I(N__14214));
    LocalMux I__1693 (
            .O(N__14222),
            .I(N__14211));
    CascadeMux I__1692 (
            .O(N__14221),
            .I(N__14208));
    InMux I__1691 (
            .O(N__14220),
            .I(N__14200));
    InMux I__1690 (
            .O(N__14219),
            .I(N__14200));
    InMux I__1689 (
            .O(N__14218),
            .I(N__14195));
    InMux I__1688 (
            .O(N__14217),
            .I(N__14195));
    LocalMux I__1687 (
            .O(N__14214),
            .I(N__14190));
    Span4Mux_v I__1686 (
            .O(N__14211),
            .I(N__14190));
    InMux I__1685 (
            .O(N__14208),
            .I(N__14187));
    InMux I__1684 (
            .O(N__14207),
            .I(N__14182));
    InMux I__1683 (
            .O(N__14206),
            .I(N__14182));
    InMux I__1682 (
            .O(N__14205),
            .I(N__14179));
    LocalMux I__1681 (
            .O(N__14200),
            .I(N__14174));
    LocalMux I__1680 (
            .O(N__14195),
            .I(N__14174));
    Span4Mux_v I__1679 (
            .O(N__14190),
            .I(N__14171));
    LocalMux I__1678 (
            .O(N__14187),
            .I(N__14168));
    LocalMux I__1677 (
            .O(N__14182),
            .I(\c0.byte_transmit_counter2_4 ));
    LocalMux I__1676 (
            .O(N__14179),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__1675 (
            .O(N__14174),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__1674 (
            .O(N__14171),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__1673 (
            .O(N__14168),
            .I(\c0.byte_transmit_counter2_4 ));
    CEMux I__1672 (
            .O(N__14157),
            .I(N__14154));
    LocalMux I__1671 (
            .O(N__14154),
            .I(N__14151));
    Odrv12 I__1670 (
            .O(N__14151),
            .I(\c0.n195 ));
    SRMux I__1669 (
            .O(N__14148),
            .I(N__14145));
    LocalMux I__1668 (
            .O(N__14145),
            .I(N__14142));
    Span4Mux_h I__1667 (
            .O(N__14142),
            .I(N__14139));
    Odrv4 I__1666 (
            .O(N__14139),
            .I(\c0.n2325 ));
    CascadeMux I__1665 (
            .O(N__14136),
            .I(N__14133));
    InMux I__1664 (
            .O(N__14133),
            .I(N__14129));
    CascadeMux I__1663 (
            .O(N__14132),
            .I(N__14120));
    LocalMux I__1662 (
            .O(N__14129),
            .I(N__14116));
    CascadeMux I__1661 (
            .O(N__14128),
            .I(N__14108));
    CascadeMux I__1660 (
            .O(N__14127),
            .I(N__14105));
    InMux I__1659 (
            .O(N__14126),
            .I(N__14101));
    InMux I__1658 (
            .O(N__14125),
            .I(N__14092));
    InMux I__1657 (
            .O(N__14124),
            .I(N__14092));
    InMux I__1656 (
            .O(N__14123),
            .I(N__14092));
    InMux I__1655 (
            .O(N__14120),
            .I(N__14089));
    InMux I__1654 (
            .O(N__14119),
            .I(N__14086));
    Span4Mux_v I__1653 (
            .O(N__14116),
            .I(N__14083));
    InMux I__1652 (
            .O(N__14115),
            .I(N__14078));
    InMux I__1651 (
            .O(N__14114),
            .I(N__14078));
    InMux I__1650 (
            .O(N__14113),
            .I(N__14071));
    InMux I__1649 (
            .O(N__14112),
            .I(N__14071));
    InMux I__1648 (
            .O(N__14111),
            .I(N__14071));
    InMux I__1647 (
            .O(N__14108),
            .I(N__14064));
    InMux I__1646 (
            .O(N__14105),
            .I(N__14064));
    InMux I__1645 (
            .O(N__14104),
            .I(N__14064));
    LocalMux I__1644 (
            .O(N__14101),
            .I(N__14061));
    InMux I__1643 (
            .O(N__14100),
            .I(N__14056));
    InMux I__1642 (
            .O(N__14099),
            .I(N__14056));
    LocalMux I__1641 (
            .O(N__14092),
            .I(N__14049));
    LocalMux I__1640 (
            .O(N__14089),
            .I(N__14049));
    LocalMux I__1639 (
            .O(N__14086),
            .I(N__14049));
    Span4Mux_v I__1638 (
            .O(N__14083),
            .I(N__14044));
    LocalMux I__1637 (
            .O(N__14078),
            .I(N__14044));
    LocalMux I__1636 (
            .O(N__14071),
            .I(r_SM_Main_2_adj_1992));
    LocalMux I__1635 (
            .O(N__14064),
            .I(r_SM_Main_2_adj_1992));
    Odrv4 I__1634 (
            .O(N__14061),
            .I(r_SM_Main_2_adj_1992));
    LocalMux I__1633 (
            .O(N__14056),
            .I(r_SM_Main_2_adj_1992));
    Odrv4 I__1632 (
            .O(N__14049),
            .I(r_SM_Main_2_adj_1992));
    Odrv4 I__1631 (
            .O(N__14044),
            .I(r_SM_Main_2_adj_1992));
    InMux I__1630 (
            .O(N__14031),
            .I(N__14028));
    LocalMux I__1629 (
            .O(N__14028),
            .I(\c0.tx2.n14 ));
    InMux I__1628 (
            .O(N__14025),
            .I(N__14021));
    InMux I__1627 (
            .O(N__14024),
            .I(N__14018));
    LocalMux I__1626 (
            .O(N__14021),
            .I(N__14013));
    LocalMux I__1625 (
            .O(N__14018),
            .I(N__14008));
    CascadeMux I__1624 (
            .O(N__14017),
            .I(N__14003));
    InMux I__1623 (
            .O(N__14016),
            .I(N__14000));
    Span4Mux_s2_h I__1622 (
            .O(N__14013),
            .I(N__13997));
    InMux I__1621 (
            .O(N__14012),
            .I(N__13992));
    InMux I__1620 (
            .O(N__14011),
            .I(N__13992));
    Span4Mux_s2_h I__1619 (
            .O(N__14008),
            .I(N__13989));
    InMux I__1618 (
            .O(N__14007),
            .I(N__13982));
    InMux I__1617 (
            .O(N__14006),
            .I(N__13982));
    InMux I__1616 (
            .O(N__14003),
            .I(N__13982));
    LocalMux I__1615 (
            .O(N__14000),
            .I(\c0.tx2.r_SM_Main_0 ));
    Odrv4 I__1614 (
            .O(N__13997),
            .I(\c0.tx2.r_SM_Main_0 ));
    LocalMux I__1613 (
            .O(N__13992),
            .I(\c0.tx2.r_SM_Main_0 ));
    Odrv4 I__1612 (
            .O(N__13989),
            .I(\c0.tx2.r_SM_Main_0 ));
    LocalMux I__1611 (
            .O(N__13982),
            .I(\c0.tx2.r_SM_Main_0 ));
    CEMux I__1610 (
            .O(N__13971),
            .I(N__13968));
    LocalMux I__1609 (
            .O(N__13968),
            .I(N__13965));
    Span4Mux_s2_h I__1608 (
            .O(N__13965),
            .I(N__13960));
    InMux I__1607 (
            .O(N__13964),
            .I(N__13957));
    InMux I__1606 (
            .O(N__13963),
            .I(N__13954));
    Odrv4 I__1605 (
            .O(N__13960),
            .I(n2208));
    LocalMux I__1604 (
            .O(N__13957),
            .I(n2208));
    LocalMux I__1603 (
            .O(N__13954),
            .I(n2208));
    SRMux I__1602 (
            .O(N__13947),
            .I(N__13944));
    LocalMux I__1601 (
            .O(N__13944),
            .I(N__13941));
    Span4Mux_v I__1600 (
            .O(N__13941),
            .I(N__13937));
    InMux I__1599 (
            .O(N__13940),
            .I(N__13934));
    Odrv4 I__1598 (
            .O(N__13937),
            .I(n2339));
    LocalMux I__1597 (
            .O(N__13934),
            .I(n2339));
    InMux I__1596 (
            .O(N__13929),
            .I(N__13922));
    InMux I__1595 (
            .O(N__13928),
            .I(N__13922));
    InMux I__1594 (
            .O(N__13927),
            .I(N__13919));
    LocalMux I__1593 (
            .O(N__13922),
            .I(N__13915));
    LocalMux I__1592 (
            .O(N__13919),
            .I(N__13909));
    InMux I__1591 (
            .O(N__13918),
            .I(N__13906));
    Span4Mux_v I__1590 (
            .O(N__13915),
            .I(N__13903));
    InMux I__1589 (
            .O(N__13914),
            .I(N__13900));
    InMux I__1588 (
            .O(N__13913),
            .I(N__13895));
    InMux I__1587 (
            .O(N__13912),
            .I(N__13895));
    Span4Mux_v I__1586 (
            .O(N__13909),
            .I(N__13890));
    LocalMux I__1585 (
            .O(N__13906),
            .I(N__13890));
    Odrv4 I__1584 (
            .O(N__13903),
            .I(r_Bit_Index_0_adj_1995));
    LocalMux I__1583 (
            .O(N__13900),
            .I(r_Bit_Index_0_adj_1995));
    LocalMux I__1582 (
            .O(N__13895),
            .I(r_Bit_Index_0_adj_1995));
    Odrv4 I__1581 (
            .O(N__13890),
            .I(r_Bit_Index_0_adj_1995));
    InMux I__1580 (
            .O(N__13881),
            .I(N__13874));
    InMux I__1579 (
            .O(N__13880),
            .I(N__13871));
    InMux I__1578 (
            .O(N__13879),
            .I(N__13868));
    InMux I__1577 (
            .O(N__13878),
            .I(N__13863));
    InMux I__1576 (
            .O(N__13877),
            .I(N__13863));
    LocalMux I__1575 (
            .O(N__13874),
            .I(\c0.tx2.r_SM_Main_2_N_1767_1 ));
    LocalMux I__1574 (
            .O(N__13871),
            .I(\c0.tx2.r_SM_Main_2_N_1767_1 ));
    LocalMux I__1573 (
            .O(N__13868),
            .I(\c0.tx2.r_SM_Main_2_N_1767_1 ));
    LocalMux I__1572 (
            .O(N__13863),
            .I(\c0.tx2.r_SM_Main_2_N_1767_1 ));
    InMux I__1571 (
            .O(N__13854),
            .I(N__13851));
    LocalMux I__1570 (
            .O(N__13851),
            .I(\c0.tx2.n5847 ));
    InMux I__1569 (
            .O(N__13848),
            .I(N__13845));
    LocalMux I__1568 (
            .O(N__13845),
            .I(\c0.rx.n3589 ));
    CascadeMux I__1567 (
            .O(N__13842),
            .I(N__13839));
    InMux I__1566 (
            .O(N__13839),
            .I(N__13836));
    LocalMux I__1565 (
            .O(N__13836),
            .I(N__13833));
    Span4Mux_s2_h I__1564 (
            .O(N__13833),
            .I(N__13830));
    Odrv4 I__1563 (
            .O(N__13830),
            .I(\c0.n6081 ));
    InMux I__1562 (
            .O(N__13827),
            .I(N__13824));
    LocalMux I__1561 (
            .O(N__13824),
            .I(N__13821));
    Span4Mux_h I__1560 (
            .O(N__13821),
            .I(N__13818));
    Span4Mux_v I__1559 (
            .O(N__13818),
            .I(N__13815));
    Odrv4 I__1558 (
            .O(N__13815),
            .I(\c0.n6084 ));
    InMux I__1557 (
            .O(N__13812),
            .I(N__13809));
    LocalMux I__1556 (
            .O(N__13809),
            .I(\c0.n5695 ));
    CascadeMux I__1555 (
            .O(N__13806),
            .I(\c0.n6234_cascade_ ));
    CascadeMux I__1554 (
            .O(N__13803),
            .I(N__13799));
    InMux I__1553 (
            .O(N__13802),
            .I(N__13793));
    InMux I__1552 (
            .O(N__13799),
            .I(N__13790));
    InMux I__1551 (
            .O(N__13798),
            .I(N__13784));
    InMux I__1550 (
            .O(N__13797),
            .I(N__13779));
    InMux I__1549 (
            .O(N__13796),
            .I(N__13779));
    LocalMux I__1548 (
            .O(N__13793),
            .I(N__13774));
    LocalMux I__1547 (
            .O(N__13790),
            .I(N__13774));
    InMux I__1546 (
            .O(N__13789),
            .I(N__13767));
    InMux I__1545 (
            .O(N__13788),
            .I(N__13767));
    InMux I__1544 (
            .O(N__13787),
            .I(N__13767));
    LocalMux I__1543 (
            .O(N__13784),
            .I(N__13761));
    LocalMux I__1542 (
            .O(N__13779),
            .I(N__13761));
    Span4Mux_h I__1541 (
            .O(N__13774),
            .I(N__13758));
    LocalMux I__1540 (
            .O(N__13767),
            .I(N__13755));
    InMux I__1539 (
            .O(N__13766),
            .I(N__13752));
    Span4Mux_v I__1538 (
            .O(N__13761),
            .I(N__13749));
    Sp12to4 I__1537 (
            .O(N__13758),
            .I(N__13744));
    Span12Mux_h I__1536 (
            .O(N__13755),
            .I(N__13744));
    LocalMux I__1535 (
            .O(N__13752),
            .I(\c0.n1081 ));
    Odrv4 I__1534 (
            .O(N__13749),
            .I(\c0.n1081 ));
    Odrv12 I__1533 (
            .O(N__13744),
            .I(\c0.n1081 ));
    CEMux I__1532 (
            .O(N__13737),
            .I(N__13733));
    CEMux I__1531 (
            .O(N__13736),
            .I(N__13729));
    LocalMux I__1530 (
            .O(N__13733),
            .I(N__13724));
    CEMux I__1529 (
            .O(N__13732),
            .I(N__13721));
    LocalMux I__1528 (
            .O(N__13729),
            .I(N__13718));
    CEMux I__1527 (
            .O(N__13728),
            .I(N__13715));
    CEMux I__1526 (
            .O(N__13727),
            .I(N__13712));
    Span4Mux_h I__1525 (
            .O(N__13724),
            .I(N__13707));
    LocalMux I__1524 (
            .O(N__13721),
            .I(N__13707));
    Span4Mux_s1_h I__1523 (
            .O(N__13718),
            .I(N__13702));
    LocalMux I__1522 (
            .O(N__13715),
            .I(N__13702));
    LocalMux I__1521 (
            .O(N__13712),
            .I(N__13699));
    Span4Mux_v I__1520 (
            .O(N__13707),
            .I(N__13696));
    Span4Mux_v I__1519 (
            .O(N__13702),
            .I(N__13693));
    Sp12to4 I__1518 (
            .O(N__13699),
            .I(N__13690));
    Span4Mux_v I__1517 (
            .O(N__13696),
            .I(N__13687));
    Odrv4 I__1516 (
            .O(N__13693),
            .I(\c0.tx2.n1624 ));
    Odrv12 I__1515 (
            .O(N__13690),
            .I(\c0.tx2.n1624 ));
    Odrv4 I__1514 (
            .O(N__13687),
            .I(\c0.tx2.n1624 ));
    InMux I__1513 (
            .O(N__13680),
            .I(N__13677));
    LocalMux I__1512 (
            .O(N__13677),
            .I(\c0.tx2.r_Tx_Data_7 ));
    InMux I__1511 (
            .O(N__13674),
            .I(N__13671));
    LocalMux I__1510 (
            .O(N__13671),
            .I(\c0.tx2.r_Tx_Data_6 ));
    CascadeMux I__1509 (
            .O(N__13668),
            .I(N__13665));
    InMux I__1508 (
            .O(N__13665),
            .I(N__13660));
    CascadeMux I__1507 (
            .O(N__13664),
            .I(N__13656));
    InMux I__1506 (
            .O(N__13663),
            .I(N__13653));
    LocalMux I__1505 (
            .O(N__13660),
            .I(N__13650));
    CascadeMux I__1504 (
            .O(N__13659),
            .I(N__13647));
    InMux I__1503 (
            .O(N__13656),
            .I(N__13641));
    LocalMux I__1502 (
            .O(N__13653),
            .I(N__13638));
    Span4Mux_v I__1501 (
            .O(N__13650),
            .I(N__13635));
    InMux I__1500 (
            .O(N__13647),
            .I(N__13630));
    InMux I__1499 (
            .O(N__13646),
            .I(N__13630));
    InMux I__1498 (
            .O(N__13645),
            .I(N__13627));
    InMux I__1497 (
            .O(N__13644),
            .I(N__13624));
    LocalMux I__1496 (
            .O(N__13641),
            .I(N__13619));
    Span4Mux_v I__1495 (
            .O(N__13638),
            .I(N__13619));
    Span4Mux_h I__1494 (
            .O(N__13635),
            .I(N__13616));
    LocalMux I__1493 (
            .O(N__13630),
            .I(\c0.tx2.r_Bit_Index_1 ));
    LocalMux I__1492 (
            .O(N__13627),
            .I(\c0.tx2.r_Bit_Index_1 ));
    LocalMux I__1491 (
            .O(N__13624),
            .I(\c0.tx2.r_Bit_Index_1 ));
    Odrv4 I__1490 (
            .O(N__13619),
            .I(\c0.tx2.r_Bit_Index_1 ));
    Odrv4 I__1489 (
            .O(N__13616),
            .I(\c0.tx2.r_Bit_Index_1 ));
    InMux I__1488 (
            .O(N__13605),
            .I(N__13602));
    LocalMux I__1487 (
            .O(N__13602),
            .I(N__13599));
    Span4Mux_v I__1486 (
            .O(N__13599),
            .I(N__13596));
    Odrv4 I__1485 (
            .O(N__13596),
            .I(\c0.tx2.n6003 ));
    CascadeMux I__1484 (
            .O(N__13593),
            .I(N__13588));
    InMux I__1483 (
            .O(N__13592),
            .I(N__13583));
    InMux I__1482 (
            .O(N__13591),
            .I(N__13583));
    InMux I__1481 (
            .O(N__13588),
            .I(N__13580));
    LocalMux I__1480 (
            .O(N__13583),
            .I(N__13577));
    LocalMux I__1479 (
            .O(N__13580),
            .I(N__13574));
    Odrv4 I__1478 (
            .O(N__13577),
            .I(\c0.FRAME_MATCHER_wait_for_transmission_N_909 ));
    Odrv4 I__1477 (
            .O(N__13574),
            .I(\c0.FRAME_MATCHER_wait_for_transmission_N_909 ));
    InMux I__1476 (
            .O(N__13569),
            .I(\c0.n4735 ));
    InMux I__1475 (
            .O(N__13566),
            .I(\c0.n4736 ));
    InMux I__1474 (
            .O(N__13563),
            .I(\c0.n4737 ));
    InMux I__1473 (
            .O(N__13560),
            .I(N__13556));
    InMux I__1472 (
            .O(N__13559),
            .I(N__13553));
    LocalMux I__1471 (
            .O(N__13556),
            .I(\c0.data_in_frame_18_5 ));
    LocalMux I__1470 (
            .O(N__13553),
            .I(\c0.data_in_frame_18_5 ));
    CascadeMux I__1469 (
            .O(N__13548),
            .I(\c0.n6225_cascade_ ));
    CascadeMux I__1468 (
            .O(N__13545),
            .I(\c0.n6228_cascade_ ));
    InMux I__1467 (
            .O(N__13542),
            .I(N__13539));
    LocalMux I__1466 (
            .O(N__13539),
            .I(N__13536));
    Span4Mux_v I__1465 (
            .O(N__13536),
            .I(N__13533));
    Odrv4 I__1464 (
            .O(N__13533),
            .I(\c0.tx2.r_Tx_Data_5 ));
    CascadeMux I__1463 (
            .O(N__13530),
            .I(\c0.n6267_cascade_ ));
    CascadeMux I__1462 (
            .O(N__13527),
            .I(\c0.n6270_cascade_ ));
    CascadeMux I__1461 (
            .O(N__13524),
            .I(N__13521));
    InMux I__1460 (
            .O(N__13521),
            .I(N__13518));
    LocalMux I__1459 (
            .O(N__13518),
            .I(N__13515));
    Span4Mux_v I__1458 (
            .O(N__13515),
            .I(N__13512));
    Odrv4 I__1457 (
            .O(N__13512),
            .I(\c0.tx2.r_Tx_Data_4 ));
    CascadeMux I__1456 (
            .O(N__13509),
            .I(N__13506));
    InMux I__1455 (
            .O(N__13506),
            .I(N__13502));
    InMux I__1454 (
            .O(N__13505),
            .I(N__13499));
    LocalMux I__1453 (
            .O(N__13502),
            .I(\c0.data_in_frame_19_3 ));
    LocalMux I__1452 (
            .O(N__13499),
            .I(\c0.data_in_frame_19_3 ));
    InMux I__1451 (
            .O(N__13494),
            .I(N__13491));
    LocalMux I__1450 (
            .O(N__13491),
            .I(N__13488));
    Odrv4 I__1449 (
            .O(N__13488),
            .I(\c0.n22_adj_1876 ));
    InMux I__1448 (
            .O(N__13485),
            .I(N__13482));
    LocalMux I__1447 (
            .O(N__13482),
            .I(N__13478));
    InMux I__1446 (
            .O(N__13481),
            .I(N__13474));
    Span4Mux_s2_h I__1445 (
            .O(N__13478),
            .I(N__13471));
    InMux I__1444 (
            .O(N__13477),
            .I(N__13468));
    LocalMux I__1443 (
            .O(N__13474),
            .I(\c0.data_in_field_49 ));
    Odrv4 I__1442 (
            .O(N__13471),
            .I(\c0.data_in_field_49 ));
    LocalMux I__1441 (
            .O(N__13468),
            .I(\c0.data_in_field_49 ));
    CascadeMux I__1440 (
            .O(N__13461),
            .I(\c0.n5991_cascade_ ));
    InMux I__1439 (
            .O(N__13458),
            .I(N__13455));
    LocalMux I__1438 (
            .O(N__13455),
            .I(N__13452));
    Span4Mux_s2_h I__1437 (
            .O(N__13452),
            .I(N__13449));
    Odrv4 I__1436 (
            .O(N__13449),
            .I(\c0.n6105 ));
    CascadeMux I__1435 (
            .O(N__13446),
            .I(\c0.n5488_cascade_ ));
    CascadeMux I__1434 (
            .O(N__13443),
            .I(\c0.n36_cascade_ ));
    InMux I__1433 (
            .O(N__13440),
            .I(N__13437));
    LocalMux I__1432 (
            .O(N__13437),
            .I(\c0.n45 ));
    InMux I__1431 (
            .O(N__13434),
            .I(N__13431));
    LocalMux I__1430 (
            .O(N__13431),
            .I(\c0.n12 ));
    InMux I__1429 (
            .O(N__13428),
            .I(N__13425));
    LocalMux I__1428 (
            .O(N__13425),
            .I(\c0.n5488 ));
    InMux I__1427 (
            .O(N__13422),
            .I(N__13419));
    LocalMux I__1426 (
            .O(N__13419),
            .I(\c0.n5489 ));
    InMux I__1425 (
            .O(N__13416),
            .I(N__13413));
    LocalMux I__1424 (
            .O(N__13413),
            .I(\c0.n1886 ));
    InMux I__1423 (
            .O(N__13410),
            .I(N__13407));
    LocalMux I__1422 (
            .O(N__13407),
            .I(\c0.n1942 ));
    InMux I__1421 (
            .O(N__13404),
            .I(N__13401));
    LocalMux I__1420 (
            .O(N__13401),
            .I(\c0.n12_adj_1951 ));
    CascadeMux I__1419 (
            .O(N__13398),
            .I(N__13395));
    InMux I__1418 (
            .O(N__13395),
            .I(N__13392));
    LocalMux I__1417 (
            .O(N__13392),
            .I(N__13389));
    Span4Mux_v I__1416 (
            .O(N__13389),
            .I(N__13384));
    InMux I__1415 (
            .O(N__13388),
            .I(N__13381));
    InMux I__1414 (
            .O(N__13387),
            .I(N__13378));
    Odrv4 I__1413 (
            .O(N__13384),
            .I(data_in_14_2));
    LocalMux I__1412 (
            .O(N__13381),
            .I(data_in_14_2));
    LocalMux I__1411 (
            .O(N__13378),
            .I(data_in_14_2));
    InMux I__1410 (
            .O(N__13371),
            .I(N__13368));
    LocalMux I__1409 (
            .O(N__13368),
            .I(N__13365));
    Span4Mux_h I__1408 (
            .O(N__13365),
            .I(N__13362));
    Odrv4 I__1407 (
            .O(N__13362),
            .I(\c0.n5536 ));
    InMux I__1406 (
            .O(N__13359),
            .I(N__13356));
    LocalMux I__1405 (
            .O(N__13356),
            .I(\c0.n5586 ));
    CascadeMux I__1404 (
            .O(N__13353),
            .I(\c0.n5381_cascade_ ));
    CascadeMux I__1403 (
            .O(N__13350),
            .I(N__13347));
    InMux I__1402 (
            .O(N__13347),
            .I(N__13343));
    InMux I__1401 (
            .O(N__13346),
            .I(N__13340));
    LocalMux I__1400 (
            .O(N__13343),
            .I(N__13336));
    LocalMux I__1399 (
            .O(N__13340),
            .I(N__13333));
    InMux I__1398 (
            .O(N__13339),
            .I(N__13330));
    Odrv4 I__1397 (
            .O(N__13336),
            .I(data_in_13_7));
    Odrv4 I__1396 (
            .O(N__13333),
            .I(data_in_13_7));
    LocalMux I__1395 (
            .O(N__13330),
            .I(data_in_13_7));
    InMux I__1394 (
            .O(N__13323),
            .I(N__13320));
    LocalMux I__1393 (
            .O(N__13320),
            .I(\c0.n2009 ));
    InMux I__1392 (
            .O(N__13317),
            .I(N__13314));
    LocalMux I__1391 (
            .O(N__13314),
            .I(N__13311));
    Span4Mux_v I__1390 (
            .O(N__13311),
            .I(N__13308));
    Span4Mux_v I__1389 (
            .O(N__13308),
            .I(N__13303));
    InMux I__1388 (
            .O(N__13307),
            .I(N__13300));
    InMux I__1387 (
            .O(N__13306),
            .I(N__13297));
    Odrv4 I__1386 (
            .O(N__13303),
            .I(data_in_16_6));
    LocalMux I__1385 (
            .O(N__13300),
            .I(data_in_16_6));
    LocalMux I__1384 (
            .O(N__13297),
            .I(data_in_16_6));
    CascadeMux I__1383 (
            .O(N__13290),
            .I(\c0.n1942_cascade_ ));
    InMux I__1382 (
            .O(N__13287),
            .I(N__13284));
    LocalMux I__1381 (
            .O(N__13284),
            .I(\c0.n18_adj_1938 ));
    CascadeMux I__1380 (
            .O(N__13281),
            .I(\c0.n5578_cascade_ ));
    InMux I__1379 (
            .O(N__13278),
            .I(N__13275));
    LocalMux I__1378 (
            .O(N__13275),
            .I(\c0.n30 ));
    CascadeMux I__1377 (
            .O(N__13272),
            .I(\c0.n6123_cascade_ ));
    CascadeMux I__1376 (
            .O(N__13269),
            .I(N__13266));
    InMux I__1375 (
            .O(N__13266),
            .I(N__13263));
    LocalMux I__1374 (
            .O(N__13263),
            .I(\c0.n5752 ));
    InMux I__1373 (
            .O(N__13260),
            .I(N__13256));
    CascadeMux I__1372 (
            .O(N__13259),
            .I(N__13253));
    LocalMux I__1371 (
            .O(N__13256),
            .I(N__13249));
    InMux I__1370 (
            .O(N__13253),
            .I(N__13244));
    InMux I__1369 (
            .O(N__13252),
            .I(N__13244));
    Odrv12 I__1368 (
            .O(N__13249),
            .I(data_in_14_7));
    LocalMux I__1367 (
            .O(N__13244),
            .I(data_in_14_7));
    InMux I__1366 (
            .O(N__13239),
            .I(N__13236));
    LocalMux I__1365 (
            .O(N__13236),
            .I(N__13233));
    Odrv4 I__1364 (
            .O(N__13233),
            .I(\c0.n24_adj_1877 ));
    CascadeMux I__1363 (
            .O(N__13230),
            .I(N__13227));
    InMux I__1362 (
            .O(N__13227),
            .I(N__13224));
    LocalMux I__1361 (
            .O(N__13224),
            .I(N__13220));
    InMux I__1360 (
            .O(N__13223),
            .I(N__13217));
    Span4Mux_v I__1359 (
            .O(N__13220),
            .I(N__13214));
    LocalMux I__1358 (
            .O(N__13217),
            .I(\c0.data_in_frame_19_2 ));
    Odrv4 I__1357 (
            .O(N__13214),
            .I(\c0.data_in_frame_19_2 ));
    InMux I__1356 (
            .O(N__13209),
            .I(N__13206));
    LocalMux I__1355 (
            .O(N__13206),
            .I(\c0.n5381 ));
    CascadeMux I__1354 (
            .O(N__13203),
            .I(\c0.n6159_cascade_ ));
    InMux I__1353 (
            .O(N__13200),
            .I(N__13197));
    LocalMux I__1352 (
            .O(N__13197),
            .I(N__13194));
    Span4Mux_s2_h I__1351 (
            .O(N__13194),
            .I(N__13191));
    Odrv4 I__1350 (
            .O(N__13191),
            .I(\c0.n5737 ));
    InMux I__1349 (
            .O(N__13188),
            .I(N__13185));
    LocalMux I__1348 (
            .O(N__13185),
            .I(\c0.n5743 ));
    InMux I__1347 (
            .O(N__13182),
            .I(N__13179));
    LocalMux I__1346 (
            .O(N__13179),
            .I(\c0.n6141 ));
    InMux I__1345 (
            .O(N__13176),
            .I(N__13171));
    InMux I__1344 (
            .O(N__13175),
            .I(N__13166));
    InMux I__1343 (
            .O(N__13174),
            .I(N__13166));
    LocalMux I__1342 (
            .O(N__13171),
            .I(\c0.tx2.r_Clock_Count_0 ));
    LocalMux I__1341 (
            .O(N__13166),
            .I(\c0.tx2.r_Clock_Count_0 ));
    InMux I__1340 (
            .O(N__13161),
            .I(N__13156));
    InMux I__1339 (
            .O(N__13160),
            .I(N__13151));
    InMux I__1338 (
            .O(N__13159),
            .I(N__13151));
    LocalMux I__1337 (
            .O(N__13156),
            .I(\c0.tx2.r_Clock_Count_1 ));
    LocalMux I__1336 (
            .O(N__13151),
            .I(\c0.tx2.r_Clock_Count_1 ));
    InMux I__1335 (
            .O(N__13146),
            .I(N__13143));
    LocalMux I__1334 (
            .O(N__13143),
            .I(\c0.tx2.n316 ));
    CascadeMux I__1333 (
            .O(N__13140),
            .I(N__13137));
    InMux I__1332 (
            .O(N__13137),
            .I(N__13132));
    InMux I__1331 (
            .O(N__13136),
            .I(N__13129));
    InMux I__1330 (
            .O(N__13135),
            .I(N__13126));
    LocalMux I__1329 (
            .O(N__13132),
            .I(\c0.tx2.r_Clock_Count_5 ));
    LocalMux I__1328 (
            .O(N__13129),
            .I(\c0.tx2.r_Clock_Count_5 ));
    LocalMux I__1327 (
            .O(N__13126),
            .I(\c0.tx2.r_Clock_Count_5 ));
    InMux I__1326 (
            .O(N__13119),
            .I(N__13113));
    InMux I__1325 (
            .O(N__13118),
            .I(N__13110));
    InMux I__1324 (
            .O(N__13117),
            .I(N__13107));
    InMux I__1323 (
            .O(N__13116),
            .I(N__13104));
    LocalMux I__1322 (
            .O(N__13113),
            .I(N__13101));
    LocalMux I__1321 (
            .O(N__13110),
            .I(\c0.tx2.r_Clock_Count_3 ));
    LocalMux I__1320 (
            .O(N__13107),
            .I(\c0.tx2.r_Clock_Count_3 ));
    LocalMux I__1319 (
            .O(N__13104),
            .I(\c0.tx2.r_Clock_Count_3 ));
    Odrv4 I__1318 (
            .O(N__13101),
            .I(\c0.tx2.r_Clock_Count_3 ));
    InMux I__1317 (
            .O(N__13092),
            .I(N__13089));
    LocalMux I__1316 (
            .O(N__13089),
            .I(N__13086));
    Odrv4 I__1315 (
            .O(N__13086),
            .I(\c0.tx2.n14_adj_1867 ));
    InMux I__1314 (
            .O(N__13083),
            .I(N__13080));
    LocalMux I__1313 (
            .O(N__13080),
            .I(N__13077));
    Odrv12 I__1312 (
            .O(N__13077),
            .I(\c0.rx.r_Rx_Data_R ));
    CascadeMux I__1311 (
            .O(N__13074),
            .I(N__13071));
    InMux I__1310 (
            .O(N__13071),
            .I(N__13065));
    InMux I__1309 (
            .O(N__13070),
            .I(N__13062));
    InMux I__1308 (
            .O(N__13069),
            .I(N__13057));
    InMux I__1307 (
            .O(N__13068),
            .I(N__13057));
    LocalMux I__1306 (
            .O(N__13065),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__1305 (
            .O(N__13062),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__1304 (
            .O(N__13057),
            .I(\c0.tx2.r_Clock_Count_7 ));
    InMux I__1303 (
            .O(N__13050),
            .I(N__13042));
    InMux I__1302 (
            .O(N__13049),
            .I(N__13042));
    InMux I__1301 (
            .O(N__13048),
            .I(N__13037));
    InMux I__1300 (
            .O(N__13047),
            .I(N__13037));
    LocalMux I__1299 (
            .O(N__13042),
            .I(r_Clock_Count_8_adj_1994));
    LocalMux I__1298 (
            .O(N__13037),
            .I(r_Clock_Count_8_adj_1994));
    CascadeMux I__1297 (
            .O(N__13032),
            .I(N__13027));
    CascadeMux I__1296 (
            .O(N__13031),
            .I(N__13023));
    CascadeMux I__1295 (
            .O(N__13030),
            .I(N__13020));
    InMux I__1294 (
            .O(N__13027),
            .I(N__13017));
    InMux I__1293 (
            .O(N__13026),
            .I(N__13014));
    InMux I__1292 (
            .O(N__13023),
            .I(N__13009));
    InMux I__1291 (
            .O(N__13020),
            .I(N__13009));
    LocalMux I__1290 (
            .O(N__13017),
            .I(\c0.tx2.r_Clock_Count_6 ));
    LocalMux I__1289 (
            .O(N__13014),
            .I(\c0.tx2.r_Clock_Count_6 ));
    LocalMux I__1288 (
            .O(N__13009),
            .I(\c0.tx2.r_Clock_Count_6 ));
    InMux I__1287 (
            .O(N__13002),
            .I(N__12998));
    InMux I__1286 (
            .O(N__13001),
            .I(N__12995));
    LocalMux I__1285 (
            .O(N__12998),
            .I(\c0.tx2.n31 ));
    LocalMux I__1284 (
            .O(N__12995),
            .I(\c0.tx2.n31 ));
    InMux I__1283 (
            .O(N__12990),
            .I(N__12987));
    LocalMux I__1282 (
            .O(N__12987),
            .I(N__12984));
    Odrv4 I__1281 (
            .O(N__12984),
            .I(\c0.tx2.n9 ));
    CascadeMux I__1280 (
            .O(N__12981),
            .I(\c0.tx2.n5631_cascade_ ));
    InMux I__1279 (
            .O(N__12978),
            .I(N__12974));
    InMux I__1278 (
            .O(N__12977),
            .I(N__12971));
    LocalMux I__1277 (
            .O(N__12974),
            .I(\c0.tx2.n78 ));
    LocalMux I__1276 (
            .O(N__12971),
            .I(\c0.tx2.n78 ));
    InMux I__1275 (
            .O(N__12966),
            .I(N__12953));
    InMux I__1274 (
            .O(N__12965),
            .I(N__12953));
    InMux I__1273 (
            .O(N__12964),
            .I(N__12950));
    InMux I__1272 (
            .O(N__12963),
            .I(N__12947));
    InMux I__1271 (
            .O(N__12962),
            .I(N__12938));
    InMux I__1270 (
            .O(N__12961),
            .I(N__12938));
    InMux I__1269 (
            .O(N__12960),
            .I(N__12938));
    InMux I__1268 (
            .O(N__12959),
            .I(N__12938));
    InMux I__1267 (
            .O(N__12958),
            .I(N__12935));
    LocalMux I__1266 (
            .O(N__12953),
            .I(N__12930));
    LocalMux I__1265 (
            .O(N__12950),
            .I(N__12930));
    LocalMux I__1264 (
            .O(N__12947),
            .I(n4544));
    LocalMux I__1263 (
            .O(N__12938),
            .I(n4544));
    LocalMux I__1262 (
            .O(N__12935),
            .I(n4544));
    Odrv4 I__1261 (
            .O(N__12930),
            .I(n4544));
    CascadeMux I__1260 (
            .O(N__12921),
            .I(N__12917));
    CascadeMux I__1259 (
            .O(N__12920),
            .I(N__12913));
    InMux I__1258 (
            .O(N__12917),
            .I(N__12909));
    InMux I__1257 (
            .O(N__12916),
            .I(N__12906));
    InMux I__1256 (
            .O(N__12913),
            .I(N__12901));
    InMux I__1255 (
            .O(N__12912),
            .I(N__12901));
    LocalMux I__1254 (
            .O(N__12909),
            .I(\c0.tx2.r_Clock_Count_4 ));
    LocalMux I__1253 (
            .O(N__12906),
            .I(\c0.tx2.r_Clock_Count_4 ));
    LocalMux I__1252 (
            .O(N__12901),
            .I(\c0.tx2.r_Clock_Count_4 ));
    CascadeMux I__1251 (
            .O(N__12894),
            .I(N__12888));
    InMux I__1250 (
            .O(N__12893),
            .I(N__12885));
    CascadeMux I__1249 (
            .O(N__12892),
            .I(N__12878));
    InMux I__1248 (
            .O(N__12891),
            .I(N__12873));
    InMux I__1247 (
            .O(N__12888),
            .I(N__12870));
    LocalMux I__1246 (
            .O(N__12885),
            .I(N__12867));
    InMux I__1245 (
            .O(N__12884),
            .I(N__12858));
    InMux I__1244 (
            .O(N__12883),
            .I(N__12858));
    InMux I__1243 (
            .O(N__12882),
            .I(N__12858));
    InMux I__1242 (
            .O(N__12881),
            .I(N__12858));
    InMux I__1241 (
            .O(N__12878),
            .I(N__12853));
    InMux I__1240 (
            .O(N__12877),
            .I(N__12853));
    InMux I__1239 (
            .O(N__12876),
            .I(N__12850));
    LocalMux I__1238 (
            .O(N__12873),
            .I(r_SM_Main_1_adj_1993));
    LocalMux I__1237 (
            .O(N__12870),
            .I(r_SM_Main_1_adj_1993));
    Odrv4 I__1236 (
            .O(N__12867),
            .I(r_SM_Main_1_adj_1993));
    LocalMux I__1235 (
            .O(N__12858),
            .I(r_SM_Main_1_adj_1993));
    LocalMux I__1234 (
            .O(N__12853),
            .I(r_SM_Main_1_adj_1993));
    LocalMux I__1233 (
            .O(N__12850),
            .I(r_SM_Main_1_adj_1993));
    CascadeMux I__1232 (
            .O(N__12837),
            .I(\c0.tx2.r_SM_Main_2_N_1767_1_cascade_ ));
    InMux I__1231 (
            .O(N__12834),
            .I(N__12831));
    LocalMux I__1230 (
            .O(N__12831),
            .I(\c0.tx2.n315 ));
    InMux I__1229 (
            .O(N__12828),
            .I(N__12825));
    LocalMux I__1228 (
            .O(N__12825),
            .I(\c0.tx2.n5824 ));
    InMux I__1227 (
            .O(N__12822),
            .I(N__12819));
    LocalMux I__1226 (
            .O(N__12819),
            .I(\c0.tx2.n5816 ));
    InMux I__1225 (
            .O(N__12816),
            .I(N__12813));
    LocalMux I__1224 (
            .O(N__12813),
            .I(N__12810));
    Odrv4 I__1223 (
            .O(N__12810),
            .I(\c0.tx2.n314 ));
    CascadeMux I__1222 (
            .O(N__12807),
            .I(N__12804));
    InMux I__1221 (
            .O(N__12804),
            .I(N__12801));
    LocalMux I__1220 (
            .O(N__12801),
            .I(\c0.tx2.n319 ));
    InMux I__1219 (
            .O(N__12798),
            .I(N__12793));
    InMux I__1218 (
            .O(N__12797),
            .I(N__12788));
    InMux I__1217 (
            .O(N__12796),
            .I(N__12788));
    LocalMux I__1216 (
            .O(N__12793),
            .I(\c0.tx2.r_Clock_Count_2 ));
    LocalMux I__1215 (
            .O(N__12788),
            .I(\c0.tx2.r_Clock_Count_2 ));
    InMux I__1214 (
            .O(N__12783),
            .I(N__12778));
    InMux I__1213 (
            .O(N__12782),
            .I(N__12775));
    InMux I__1212 (
            .O(N__12781),
            .I(N__12772));
    LocalMux I__1211 (
            .O(N__12778),
            .I(\c0.tx2.r_Bit_Index_2 ));
    LocalMux I__1210 (
            .O(N__12775),
            .I(\c0.tx2.r_Bit_Index_2 ));
    LocalMux I__1209 (
            .O(N__12772),
            .I(\c0.tx2.r_Bit_Index_2 ));
    CascadeMux I__1208 (
            .O(N__12765),
            .I(N__12761));
    InMux I__1207 (
            .O(N__12764),
            .I(N__12758));
    InMux I__1206 (
            .O(N__12761),
            .I(N__12755));
    LocalMux I__1205 (
            .O(N__12758),
            .I(\c0.tx2.n1136 ));
    LocalMux I__1204 (
            .O(N__12755),
            .I(\c0.tx2.n1136 ));
    CascadeMux I__1203 (
            .O(N__12750),
            .I(n4_adj_1973_cascade_));
    InMux I__1202 (
            .O(N__12747),
            .I(N__12742));
    InMux I__1201 (
            .O(N__12746),
            .I(N__12737));
    InMux I__1200 (
            .O(N__12745),
            .I(N__12737));
    LocalMux I__1199 (
            .O(N__12742),
            .I(tx2_active));
    LocalMux I__1198 (
            .O(N__12737),
            .I(tx2_active));
    CascadeMux I__1197 (
            .O(N__12732),
            .I(N__12726));
    CascadeMux I__1196 (
            .O(N__12731),
            .I(N__12723));
    InMux I__1195 (
            .O(N__12730),
            .I(N__12717));
    InMux I__1194 (
            .O(N__12729),
            .I(N__12717));
    InMux I__1193 (
            .O(N__12726),
            .I(N__12710));
    InMux I__1192 (
            .O(N__12723),
            .I(N__12710));
    InMux I__1191 (
            .O(N__12722),
            .I(N__12710));
    LocalMux I__1190 (
            .O(N__12717),
            .I(\c0.r_SM_Main_2_N_1770_0 ));
    LocalMux I__1189 (
            .O(N__12710),
            .I(\c0.r_SM_Main_2_N_1770_0 ));
    IoInMux I__1188 (
            .O(N__12705),
            .I(N__12701));
    InMux I__1187 (
            .O(N__12704),
            .I(N__12698));
    LocalMux I__1186 (
            .O(N__12701),
            .I(N__12695));
    LocalMux I__1185 (
            .O(N__12698),
            .I(N__12692));
    Span4Mux_s1_h I__1184 (
            .O(N__12695),
            .I(N__12688));
    Span4Mux_v I__1183 (
            .O(N__12692),
            .I(N__12685));
    InMux I__1182 (
            .O(N__12691),
            .I(N__12682));
    Odrv4 I__1181 (
            .O(N__12688),
            .I(tx2_o));
    Odrv4 I__1180 (
            .O(N__12685),
            .I(tx2_o));
    LocalMux I__1179 (
            .O(N__12682),
            .I(tx2_o));
    IoInMux I__1178 (
            .O(N__12675),
            .I(N__12672));
    LocalMux I__1177 (
            .O(N__12672),
            .I(N__12669));
    Odrv4 I__1176 (
            .O(N__12669),
            .I(tx2_enable));
    CascadeMux I__1175 (
            .O(N__12666),
            .I(N__12663));
    InMux I__1174 (
            .O(N__12663),
            .I(N__12660));
    LocalMux I__1173 (
            .O(N__12660),
            .I(N__12657));
    Odrv12 I__1172 (
            .O(N__12657),
            .I(\c0.n6117 ));
    CascadeMux I__1171 (
            .O(N__12654),
            .I(\c0.n5536_cascade_ ));
    CascadeMux I__1170 (
            .O(N__12651),
            .I(\c0.n5570_cascade_ ));
    InMux I__1169 (
            .O(N__12648),
            .I(N__12645));
    LocalMux I__1168 (
            .O(N__12645),
            .I(\c0.n27_adj_1910 ));
    CascadeMux I__1167 (
            .O(N__12642),
            .I(\c0.n3689_cascade_ ));
    InMux I__1166 (
            .O(N__12639),
            .I(N__12636));
    LocalMux I__1165 (
            .O(N__12636),
            .I(\c0.tx2.n12 ));
    InMux I__1164 (
            .O(N__12633),
            .I(N__12630));
    LocalMux I__1163 (
            .O(N__12630),
            .I(\c0.n3689 ));
    InMux I__1162 (
            .O(N__12627),
            .I(N__12624));
    LocalMux I__1161 (
            .O(N__12624),
            .I(N__12619));
    InMux I__1160 (
            .O(N__12623),
            .I(N__12614));
    InMux I__1159 (
            .O(N__12622),
            .I(N__12614));
    Odrv4 I__1158 (
            .O(N__12619),
            .I(\c0.n3703 ));
    LocalMux I__1157 (
            .O(N__12614),
            .I(\c0.n3703 ));
    CascadeMux I__1156 (
            .O(N__12609),
            .I(\c0.n6282_cascade_ ));
    InMux I__1155 (
            .O(N__12606),
            .I(N__12603));
    LocalMux I__1154 (
            .O(N__12603),
            .I(N__12600));
    Span4Mux_v I__1153 (
            .O(N__12600),
            .I(N__12597));
    Odrv4 I__1152 (
            .O(N__12597),
            .I(\c0.n6132 ));
    InMux I__1151 (
            .O(N__12594),
            .I(N__12591));
    LocalMux I__1150 (
            .O(N__12591),
            .I(\c0.tx2.r_Tx_Data_3 ));
    CascadeMux I__1149 (
            .O(N__12588),
            .I(N__12585));
    InMux I__1148 (
            .O(N__12585),
            .I(N__12582));
    LocalMux I__1147 (
            .O(N__12582),
            .I(\c0.n6069 ));
    CascadeMux I__1146 (
            .O(N__12579),
            .I(\c0.n6249_cascade_ ));
    InMux I__1145 (
            .O(N__12576),
            .I(N__12573));
    LocalMux I__1144 (
            .O(N__12573),
            .I(N__12570));
    Odrv4 I__1143 (
            .O(N__12570),
            .I(\c0.n28 ));
    CascadeMux I__1142 (
            .O(N__12567),
            .I(\c0.n3703_cascade_ ));
    InMux I__1141 (
            .O(N__12564),
            .I(N__12561));
    LocalMux I__1140 (
            .O(N__12561),
            .I(\c0.n47 ));
    CascadeMux I__1139 (
            .O(N__12558),
            .I(\c0.n52_cascade_ ));
    InMux I__1138 (
            .O(N__12555),
            .I(N__12552));
    LocalMux I__1137 (
            .O(N__12552),
            .I(\c0.n31 ));
    InMux I__1136 (
            .O(N__12549),
            .I(N__12546));
    LocalMux I__1135 (
            .O(N__12546),
            .I(N__12543));
    Odrv4 I__1134 (
            .O(N__12543),
            .I(\c0.n32 ));
    CascadeMux I__1133 (
            .O(N__12540),
            .I(\c0.n24_adj_1879_cascade_ ));
    InMux I__1132 (
            .O(N__12537),
            .I(N__12534));
    LocalMux I__1131 (
            .O(N__12534),
            .I(N__12531));
    Odrv12 I__1130 (
            .O(N__12531),
            .I(\c0.n6102 ));
    InMux I__1129 (
            .O(N__12528),
            .I(N__12525));
    LocalMux I__1128 (
            .O(N__12525),
            .I(\c0.tx2.r_Tx_Data_2 ));
    InMux I__1127 (
            .O(N__12522),
            .I(N__12519));
    LocalMux I__1126 (
            .O(N__12519),
            .I(N__12516));
    Odrv4 I__1125 (
            .O(N__12516),
            .I(\c0.tx2.n6045 ));
    InMux I__1124 (
            .O(N__12513),
            .I(N__12510));
    LocalMux I__1123 (
            .O(N__12510),
            .I(N__12506));
    InMux I__1122 (
            .O(N__12509),
            .I(N__12503));
    Span4Mux_v I__1121 (
            .O(N__12506),
            .I(N__12500));
    LocalMux I__1120 (
            .O(N__12503),
            .I(\c0.data_in_frame_18_2 ));
    Odrv4 I__1119 (
            .O(N__12500),
            .I(\c0.data_in_frame_18_2 ));
    CascadeMux I__1118 (
            .O(N__12495),
            .I(\c0.n6297_cascade_ ));
    CascadeMux I__1117 (
            .O(N__12492),
            .I(N__12489));
    InMux I__1116 (
            .O(N__12489),
            .I(N__12486));
    LocalMux I__1115 (
            .O(N__12486),
            .I(\c0.n6300 ));
    InMux I__1114 (
            .O(N__12483),
            .I(N__12480));
    LocalMux I__1113 (
            .O(N__12480),
            .I(N__12476));
    InMux I__1112 (
            .O(N__12479),
            .I(N__12473));
    Span4Mux_v I__1111 (
            .O(N__12476),
            .I(N__12470));
    LocalMux I__1110 (
            .O(N__12473),
            .I(\c0.data_in_frame_18_3 ));
    Odrv4 I__1109 (
            .O(N__12470),
            .I(\c0.data_in_frame_18_3 ));
    CascadeMux I__1108 (
            .O(N__12465),
            .I(\c0.n6279_cascade_ ));
    CascadeMux I__1107 (
            .O(N__12462),
            .I(\c0.n6075_cascade_ ));
    InMux I__1106 (
            .O(N__12459),
            .I(N__12456));
    LocalMux I__1105 (
            .O(N__12456),
            .I(\c0.n5773 ));
    CascadeMux I__1104 (
            .O(N__12453),
            .I(\c0.n5454_cascade_ ));
    CascadeMux I__1103 (
            .O(N__12450),
            .I(\c0.n27_cascade_ ));
    CascadeMux I__1102 (
            .O(N__12447),
            .I(N__12444));
    InMux I__1101 (
            .O(N__12444),
            .I(N__12441));
    LocalMux I__1100 (
            .O(N__12441),
            .I(\c0.n6063 ));
    InMux I__1099 (
            .O(N__12438),
            .I(N__12435));
    LocalMux I__1098 (
            .O(N__12435),
            .I(\c0.n5776 ));
    InMux I__1097 (
            .O(N__12432),
            .I(N__12429));
    LocalMux I__1096 (
            .O(N__12429),
            .I(\c0.n6099 ));
    InMux I__1095 (
            .O(N__12426),
            .I(N__12423));
    LocalMux I__1094 (
            .O(N__12423),
            .I(N__12420));
    Span4Mux_v I__1093 (
            .O(N__12420),
            .I(N__12417));
    Odrv4 I__1092 (
            .O(N__12417),
            .I(\c0.tx2.n6006 ));
    CascadeMux I__1091 (
            .O(N__12414),
            .I(\c0.n5375_cascade_ ));
    InMux I__1090 (
            .O(N__12411),
            .I(N__12408));
    LocalMux I__1089 (
            .O(N__12408),
            .I(N__12405));
    Odrv4 I__1088 (
            .O(N__12405),
            .I(\c0.n5755 ));
    CascadeMux I__1087 (
            .O(N__12402),
            .I(\c0.n6135_cascade_ ));
    CascadeMux I__1086 (
            .O(N__12399),
            .I(\c0.n5746_cascade_ ));
    CascadeMux I__1085 (
            .O(N__12396),
            .I(\c0.n6153_cascade_ ));
    CascadeMux I__1084 (
            .O(N__12393),
            .I(\c0.n5740_cascade_ ));
    InMux I__1083 (
            .O(N__12390),
            .I(N__12387));
    LocalMux I__1082 (
            .O(N__12387),
            .I(\c0.n6129 ));
    InMux I__1081 (
            .O(N__12384),
            .I(\c0.tx2.n4779 ));
    InMux I__1080 (
            .O(N__12381),
            .I(\c0.tx2.n4780 ));
    InMux I__1079 (
            .O(N__12378),
            .I(N__12375));
    LocalMux I__1078 (
            .O(N__12375),
            .I(\c0.tx2.n318 ));
    InMux I__1077 (
            .O(N__12372),
            .I(\c0.tx2.n4781 ));
    InMux I__1076 (
            .O(N__12369),
            .I(N__12366));
    LocalMux I__1075 (
            .O(N__12366),
            .I(\c0.tx2.n317 ));
    InMux I__1074 (
            .O(N__12363),
            .I(\c0.tx2.n4782 ));
    InMux I__1073 (
            .O(N__12360),
            .I(\c0.tx2.n4783 ));
    InMux I__1072 (
            .O(N__12357),
            .I(\c0.tx2.n4784 ));
    InMux I__1071 (
            .O(N__12354),
            .I(\c0.tx2.n4785 ));
    InMux I__1070 (
            .O(N__12351),
            .I(bfn_1_30_0_));
    InMux I__1069 (
            .O(N__12348),
            .I(N__12345));
    LocalMux I__1068 (
            .O(N__12345),
            .I(n313_adj_1997));
    CascadeMux I__1067 (
            .O(N__12342),
            .I(\c0.tx2.o_Tx_Serial_N_1798_cascade_ ));
    InMux I__1066 (
            .O(N__12339),
            .I(bfn_1_29_0_));
    CascadeMux I__1065 (
            .O(N__12336),
            .I(\c0.n6027_cascade_ ));
    CascadeMux I__1064 (
            .O(N__12333),
            .I(\c0.n5794_cascade_ ));
    InMux I__1063 (
            .O(N__12330),
            .I(N__12327));
    LocalMux I__1062 (
            .O(N__12327),
            .I(\c0.n6015 ));
    CascadeMux I__1061 (
            .O(N__12324),
            .I(\c0.n6072_cascade_ ));
    InMux I__1060 (
            .O(N__12321),
            .I(N__12318));
    LocalMux I__1059 (
            .O(N__12318),
            .I(\c0.n6018 ));
    InMux I__1058 (
            .O(N__12315),
            .I(N__12312));
    LocalMux I__1057 (
            .O(N__12312),
            .I(N__12309));
    Span4Mux_v I__1056 (
            .O(N__12309),
            .I(N__12306));
    Odrv4 I__1055 (
            .O(N__12306),
            .I(\c0.tx2.r_Tx_Data_1 ));
    CascadeMux I__1054 (
            .O(N__12303),
            .I(N__12300));
    InMux I__1053 (
            .O(N__12300),
            .I(N__12297));
    LocalMux I__1052 (
            .O(N__12297),
            .I(N__12294));
    Odrv4 I__1051 (
            .O(N__12294),
            .I(\c0.tx2.r_Tx_Data_0 ));
    CascadeMux I__1050 (
            .O(N__12291),
            .I(\c0.tx2.n6048_cascade_ ));
    CascadeMux I__1049 (
            .O(N__12288),
            .I(\c0.n6057_cascade_ ));
    InMux I__1048 (
            .O(N__12285),
            .I(N__12282));
    LocalMux I__1047 (
            .O(N__12282),
            .I(\c0.n6306 ));
    CascadeMux I__1046 (
            .O(N__12279),
            .I(\c0.n6060_cascade_ ));
    InMux I__1045 (
            .O(N__12276),
            .I(N__12273));
    LocalMux I__1044 (
            .O(N__12273),
            .I(\c0.n6087 ));
    InMux I__1043 (
            .O(N__12270),
            .I(N__12267));
    LocalMux I__1042 (
            .O(N__12267),
            .I(N__12264));
    Odrv12 I__1041 (
            .O(N__12264),
            .I(\c0.n5770 ));
    CascadeMux I__1040 (
            .O(N__12261),
            .I(\c0.n5788_cascade_ ));
    CascadeMux I__1039 (
            .O(N__12258),
            .I(\c0.n6111_cascade_ ));
    CascadeMux I__1038 (
            .O(N__12255),
            .I(\c0.n5758_cascade_ ));
    InMux I__1037 (
            .O(N__12252),
            .I(N__12249));
    LocalMux I__1036 (
            .O(N__12249),
            .I(\c0.n5761 ));
    InMux I__1035 (
            .O(N__12246),
            .I(N__12242));
    InMux I__1034 (
            .O(N__12245),
            .I(N__12239));
    LocalMux I__1033 (
            .O(N__12242),
            .I(N__12236));
    LocalMux I__1032 (
            .O(N__12239),
            .I(\c0.data_in_frame_18_1 ));
    Odrv4 I__1031 (
            .O(N__12236),
            .I(\c0.data_in_frame_18_1 ));
    CascadeMux I__1030 (
            .O(N__12231),
            .I(N__12228));
    InMux I__1029 (
            .O(N__12228),
            .I(N__12224));
    InMux I__1028 (
            .O(N__12227),
            .I(N__12221));
    LocalMux I__1027 (
            .O(N__12224),
            .I(N__12218));
    LocalMux I__1026 (
            .O(N__12221),
            .I(\c0.data_in_frame_19_1 ));
    Odrv4 I__1025 (
            .O(N__12218),
            .I(\c0.data_in_frame_19_1 ));
    CascadeMux I__1024 (
            .O(N__12213),
            .I(\c0.n6303_cascade_ ));
    IoInMux I__1023 (
            .O(N__12210),
            .I(N__12207));
    LocalMux I__1022 (
            .O(N__12207),
            .I(N__12204));
    IoSpan4Mux I__1021 (
            .O(N__12204),
            .I(N__12201));
    IoSpan4Mux I__1020 (
            .O(N__12201),
            .I(N__12198));
    IoSpan4Mux I__1019 (
            .O(N__12198),
            .I(N__12195));
    Odrv4 I__1018 (
            .O(N__12195),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_1_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_29_0_));
    defparam IN_MUX_bfv_1_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_30_0_ (
            .carryinitin(\c0.tx2.n4786 ),
            .carryinitout(bfn_1_30_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\c0.tx.n4771 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_4_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_27_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\c0.n4761 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_15_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_27_0_ (
            .carryinitin(\c0.n4746 ),
            .carryinitout(bfn_15_27_0_));
    defparam IN_MUX_bfv_3_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_26_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(n4717),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_14_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_27_0_ (
            .carryinitin(n4725),
            .carryinitout(bfn_14_27_0_));
    defparam IN_MUX_bfv_14_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_28_0_ (
            .carryinitin(n4733),
            .carryinitout(bfn_14_28_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__12210),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.data_in_0___i16_LC_1_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i16_LC_1_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i16_LC_1_17_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i16_LC_1_17_0  (
            .in0(N__35977),
            .in1(N__18121),
            .in2(_gnd_net_),
            .in3(N__16430),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37462),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i146_LC_1_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i146_LC_1_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i146_LC_1_17_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i146_LC_1_17_4  (
            .in0(N__12245),
            .in1(N__15161),
            .in2(N__33217),
            .in3(N__32111),
            .lcout(\c0.data_in_frame_18_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37462),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i154_LC_1_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i154_LC_1_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i154_LC_1_18_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i154_LC_1_18_6  (
            .in0(N__12227),
            .in1(N__32144),
            .in2(N__26730),
            .in3(N__33083),
            .lcout(\c0.data_in_frame_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37464),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5749_LC_1_19_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5749_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5749_LC_1_19_0 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5749_LC_1_19_0  (
            .in0(N__27756),
            .in1(N__19593),
            .in2(N__30175),
            .in3(N__23310),
            .lcout(),
            .ltout(\c0.n6111_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6111_bdd_4_lut_LC_1_19_1 .C_ON=1'b0;
    defparam \c0.n6111_bdd_4_lut_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.n6111_bdd_4_lut_LC_1_19_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6111_bdd_4_lut_LC_1_19_1  (
            .in0(N__30105),
            .in1(N__31014),
            .in2(N__12258),
            .in3(N__20958),
            .lcout(),
            .ltout(\c0.n5758_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5759_LC_1_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5759_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5759_LC_1_19_2 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5759_LC_1_19_2  (
            .in0(N__25257),
            .in1(N__25382),
            .in2(N__12255),
            .in3(N__12252),
            .lcout(\c0.n6099 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1047_2_lut_LC_1_19_5 .C_ON=1'b0;
    defparam \c0.i1047_2_lut_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1047_2_lut_LC_1_19_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1047_2_lut_LC_1_19_5  (
            .in0(N__25381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25256),
            .lcout(\c0.n1081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6105_bdd_4_lut_LC_1_19_7 .C_ON=1'b0;
    defparam \c0.n6105_bdd_4_lut_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.n6105_bdd_4_lut_LC_1_19_7 .LUT_INIT=16'b1010101011100100;
    LogicCell40 \c0.n6105_bdd_4_lut_LC_1_19_7  (
            .in0(N__13458),
            .in1(N__28310),
            .in2(N__27299),
            .in3(N__30101),
            .lcout(\c0.n5761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_20_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_20_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_20_0  (
            .in0(N__12246),
            .in1(N__30110),
            .in2(N__12231),
            .in3(N__27719),
            .lcout(),
            .ltout(\c0.n6303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6303_bdd_4_lut_LC_1_20_1 .C_ON=1'b0;
    defparam \c0.n6303_bdd_4_lut_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.n6303_bdd_4_lut_LC_1_20_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6303_bdd_4_lut_LC_1_20_1  (
            .in0(N__30111),
            .in1(N__30896),
            .in2(N__12213),
            .in3(N__17133),
            .lcout(\c0.n6306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5734_LC_1_20_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5734_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5734_LC_1_20_2 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5734_LC_1_20_2  (
            .in0(N__25260),
            .in1(N__12459),
            .in2(N__25407),
            .in3(N__12438),
            .lcout(),
            .ltout(\c0.n6057_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6057_bdd_4_lut_LC_1_20_3 .C_ON=1'b0;
    defparam \c0.n6057_bdd_4_lut_LC_1_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6057_bdd_4_lut_LC_1_20_3 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n6057_bdd_4_lut_LC_1_20_3  (
            .in0(N__15927),
            .in1(N__25390),
            .in2(N__12288),
            .in3(N__12270),
            .lcout(),
            .ltout(\c0.n6060_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i1_LC_1_20_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i1_LC_1_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i1_LC_1_20_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.tx2.r_Tx_Data_i1_LC_1_20_4  (
            .in0(N__12285),
            .in1(N__14226),
            .in2(N__12279),
            .in3(N__13766),
            .lcout(\c0.tx2.r_Tx_Data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37469),
            .ce(N__13736),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5729_LC_1_21_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5729_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5729_LC_1_21_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5729_LC_1_21_2  (
            .in0(N__27716),
            .in1(N__24316),
            .in2(N__30176),
            .in3(N__13485),
            .lcout(\c0.n6087 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6081_bdd_4_lut_LC_1_21_4 .C_ON=1'b0;
    defparam \c0.n6081_bdd_4_lut_LC_1_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.n6081_bdd_4_lut_LC_1_21_4 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6081_bdd_4_lut_LC_1_21_4  (
            .in0(N__30109),
            .in1(N__27098),
            .in2(N__13842),
            .in3(N__17289),
            .lcout(\c0.n6084 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_LC_1_21_5 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_1_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i20_4_lut_LC_1_21_5  (
            .in0(N__15657),
            .in1(N__29433),
            .in2(N__14511),
            .in3(N__24918),
            .lcout(\c0.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6087_bdd_4_lut_LC_1_22_1 .C_ON=1'b0;
    defparam \c0.n6087_bdd_4_lut_LC_1_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.n6087_bdd_4_lut_LC_1_22_1 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n6087_bdd_4_lut_LC_1_22_1  (
            .in0(N__29949),
            .in1(N__16869),
            .in2(N__18921),
            .in3(N__12276),
            .lcout(\c0.n5770 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6039_bdd_4_lut_LC_1_22_2 .C_ON=1'b0;
    defparam \c0.n6039_bdd_4_lut_LC_1_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.n6039_bdd_4_lut_LC_1_22_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6039_bdd_4_lut_LC_1_22_2  (
            .in0(N__29947),
            .in1(N__22242),
            .in2(N__27414),
            .in3(N__15300),
            .lcout(),
            .ltout(\c0.n5788_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6015_bdd_4_lut_LC_1_22_3 .C_ON=1'b0;
    defparam \c0.n6015_bdd_4_lut_LC_1_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6015_bdd_4_lut_LC_1_22_3 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n6015_bdd_4_lut_LC_1_22_3  (
            .in0(N__25392),
            .in1(N__26751),
            .in2(N__12261),
            .in3(N__12330),
            .lcout(\c0.n6018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5680_LC_1_22_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5680_LC_1_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5680_LC_1_22_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5680_LC_1_22_4  (
            .in0(N__27717),
            .in1(N__28356),
            .in2(N__30070),
            .in3(N__21984),
            .lcout(),
            .ltout(\c0.n6027_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6027_bdd_4_lut_LC_1_22_5 .C_ON=1'b0;
    defparam \c0.n6027_bdd_4_lut_LC_1_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.n6027_bdd_4_lut_LC_1_22_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6027_bdd_4_lut_LC_1_22_5  (
            .in0(N__29948),
            .in1(N__25803),
            .in2(N__12336),
            .in3(N__16794),
            .lcout(),
            .ltout(\c0.n5794_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5699_LC_1_22_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5699_LC_1_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5699_LC_1_22_6 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5699_LC_1_22_6  (
            .in0(N__25391),
            .in1(N__25247),
            .in2(N__12333),
            .in3(N__14895),
            .lcout(\c0.n6015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6069_bdd_4_lut_LC_1_23_1 .C_ON=1'b0;
    defparam \c0.n6069_bdd_4_lut_LC_1_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.n6069_bdd_4_lut_LC_1_23_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6069_bdd_4_lut_LC_1_23_1  (
            .in0(N__29999),
            .in1(N__28065),
            .in2(N__12588),
            .in3(N__30573),
            .lcout(),
            .ltout(\c0.n6072_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i0_LC_1_23_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i0_LC_1_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i0_LC_1_23_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i0_LC_1_23_2  (
            .in0(N__14225),
            .in1(N__13798),
            .in2(N__12324),
            .in3(N__12321),
            .lcout(\c0.tx2.r_Tx_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37485),
            .ce(N__13728),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i123_LC_1_24_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i123_LC_1_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i123_LC_1_24_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i123_LC_1_24_5  (
            .in0(N__35682),
            .in1(N__19294),
            .in2(_gnd_net_),
            .in3(N__15914),
            .lcout(data_in_15_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37490),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i107_LC_1_25_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i107_LC_1_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i107_LC_1_25_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i107_LC_1_25_0  (
            .in0(N__35683),
            .in1(N__13388),
            .in2(_gnd_net_),
            .in3(N__28367),
            .lcout(data_in_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37500),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n6045_bdd_4_lut_LC_1_25_3 .C_ON=1'b0;
    defparam \c0.tx2.n6045_bdd_4_lut_LC_1_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n6045_bdd_4_lut_LC_1_25_3 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.tx2.n6045_bdd_4_lut_LC_1_25_3  (
            .in0(N__12315),
            .in1(N__13645),
            .in2(N__12303),
            .in3(N__12522),
            .lcout(),
            .ltout(\c0.tx2.n6048_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i367224_i1_3_lut_LC_1_25_4 .C_ON=1'b0;
    defparam \c0.tx2.i367224_i1_3_lut_LC_1_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i367224_i1_3_lut_LC_1_25_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.tx2.i367224_i1_3_lut_LC_1_25_4  (
            .in0(_gnd_net_),
            .in1(N__12781),
            .in2(N__12291),
            .in3(N__12426),
            .lcout(),
            .ltout(\c0.tx2.o_Tx_Serial_N_1798_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i26_3_lut_LC_1_25_5 .C_ON=1'b0;
    defparam \c0.tx2.i26_3_lut_LC_1_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i26_3_lut_LC_1_25_5 .LUT_INIT=16'b0000001111001100;
    LogicCell40 \c0.tx2.i26_3_lut_LC_1_25_5  (
            .in0(_gnd_net_),
            .in1(N__14024),
            .in2(N__12342),
            .in3(N__12893),
            .lcout(\c0.tx2.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i2_LC_1_26_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i2_LC_1_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i2_LC_1_26_0 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \c0.tx2.r_Bit_Index_i2_LC_1_26_0  (
            .in0(N__13929),
            .in1(_gnd_net_),
            .in2(N__13659),
            .in3(N__12783),
            .lcout(\c0.tx2.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37509),
            .ce(N__13971),
            .sr(N__13947));
    defparam \c0.tx2.r_Bit_Index_i1_LC_1_26_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i1_LC_1_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i1_LC_1_26_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.tx2.r_Bit_Index_i1_LC_1_26_1  (
            .in0(_gnd_net_),
            .in1(N__13646),
            .in2(_gnd_net_),
            .in3(N__13928),
            .lcout(\c0.tx2.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37509),
            .ce(N__13971),
            .sr(N__13947));
    defparam \c0.data_in_0___i143_LC_1_27_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i143_LC_1_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i143_LC_1_27_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i143_LC_1_27_1  (
            .in0(N__35509),
            .in1(N__18976),
            .in2(_gnd_net_),
            .in3(N__16145),
            .lcout(data_in_17_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37520),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i135_LC_1_27_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i135_LC_1_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i135_LC_1_27_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i135_LC_1_27_4  (
            .in0(N__18977),
            .in1(N__35510),
            .in2(_gnd_net_),
            .in3(N__13306),
            .lcout(data_in_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37520),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i3_LC_1_28_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i3_LC_1_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i3_LC_1_28_0 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i3_LC_1_28_0  (
            .in0(N__12965),
            .in1(N__12378),
            .in2(N__14128),
            .in3(N__13118),
            .lcout(\c0.tx2.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i4_LC_1_28_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i4_LC_1_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i4_LC_1_28_1 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i4_LC_1_28_1  (
            .in0(N__12369),
            .in1(N__14104),
            .in2(N__12921),
            .in3(N__12966),
            .lcout(\c0.tx2.r_Clock_Count_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i2_LC_1_28_2 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i2_LC_1_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i2_LC_1_28_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.tx2.r_SM_Main_i2_LC_1_28_2  (
            .in0(N__14025),
            .in1(N__12891),
            .in2(N__14127),
            .in3(N__13881),
            .lcout(r_SM_Main_2_adj_1992),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i127_LC_1_28_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i127_LC_1_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i127_LC_1_28_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i127_LC_1_28_5  (
            .in0(N__35500),
            .in1(N__13307),
            .in2(_gnd_net_),
            .in3(N__17708),
            .lcout(data_in_15_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37532),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_2_lut_LC_1_29_0 .C_ON=1'b1;
    defparam \c0.tx2.add_59_2_lut_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_2_lut_LC_1_29_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_2_lut_LC_1_29_0  (
            .in0(N__12964),
            .in1(N__13176),
            .in2(_gnd_net_),
            .in3(N__12339),
            .lcout(\c0.tx2.n5824 ),
            .ltout(),
            .carryin(bfn_1_29_0_),
            .carryout(\c0.tx2.n4779 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_3_lut_LC_1_29_1 .C_ON=1'b1;
    defparam \c0.tx2.add_59_3_lut_LC_1_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_3_lut_LC_1_29_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_3_lut_LC_1_29_1  (
            .in0(N__12958),
            .in1(N__13161),
            .in2(_gnd_net_),
            .in3(N__12384),
            .lcout(\c0.tx2.n5816 ),
            .ltout(),
            .carryin(\c0.tx2.n4779 ),
            .carryout(\c0.tx2.n4780 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_4_lut_LC_1_29_2 .C_ON=1'b1;
    defparam \c0.tx2.add_59_4_lut_LC_1_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_4_lut_LC_1_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_4_lut_LC_1_29_2  (
            .in0(_gnd_net_),
            .in1(N__12798),
            .in2(_gnd_net_),
            .in3(N__12381),
            .lcout(\c0.tx2.n319 ),
            .ltout(),
            .carryin(\c0.tx2.n4780 ),
            .carryout(\c0.tx2.n4781 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_5_lut_LC_1_29_3 .C_ON=1'b1;
    defparam \c0.tx2.add_59_5_lut_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_5_lut_LC_1_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_5_lut_LC_1_29_3  (
            .in0(_gnd_net_),
            .in1(N__13117),
            .in2(_gnd_net_),
            .in3(N__12372),
            .lcout(\c0.tx2.n318 ),
            .ltout(),
            .carryin(\c0.tx2.n4781 ),
            .carryout(\c0.tx2.n4782 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_6_lut_LC_1_29_4 .C_ON=1'b1;
    defparam \c0.tx2.add_59_6_lut_LC_1_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_6_lut_LC_1_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_6_lut_LC_1_29_4  (
            .in0(_gnd_net_),
            .in1(N__12916),
            .in2(_gnd_net_),
            .in3(N__12363),
            .lcout(\c0.tx2.n317 ),
            .ltout(),
            .carryin(\c0.tx2.n4782 ),
            .carryout(\c0.tx2.n4783 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_7_lut_LC_1_29_5 .C_ON=1'b1;
    defparam \c0.tx2.add_59_7_lut_LC_1_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_7_lut_LC_1_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_7_lut_LC_1_29_5  (
            .in0(_gnd_net_),
            .in1(N__13136),
            .in2(_gnd_net_),
            .in3(N__12360),
            .lcout(\c0.tx2.n316 ),
            .ltout(),
            .carryin(\c0.tx2.n4783 ),
            .carryout(\c0.tx2.n4784 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_8_lut_LC_1_29_6 .C_ON=1'b1;
    defparam \c0.tx2.add_59_8_lut_LC_1_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_8_lut_LC_1_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_8_lut_LC_1_29_6  (
            .in0(_gnd_net_),
            .in1(N__13026),
            .in2(_gnd_net_),
            .in3(N__12357),
            .lcout(\c0.tx2.n315 ),
            .ltout(),
            .carryin(\c0.tx2.n4784 ),
            .carryout(\c0.tx2.n4785 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_9_lut_LC_1_29_7 .C_ON=1'b1;
    defparam \c0.tx2.add_59_9_lut_LC_1_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_9_lut_LC_1_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_9_lut_LC_1_29_7  (
            .in0(_gnd_net_),
            .in1(N__13070),
            .in2(_gnd_net_),
            .in3(N__12354),
            .lcout(\c0.tx2.n314 ),
            .ltout(),
            .carryin(\c0.tx2.n4785 ),
            .carryout(\c0.tx2.n4786 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_10_lut_LC_1_30_0 .C_ON=1'b0;
    defparam \c0.tx2.add_59_10_lut_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_10_lut_LC_1_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_10_lut_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(N__13049),
            .in2(_gnd_net_),
            .in3(N__12351),
            .lcout(n313_adj_1997),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_30_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_30_3 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i8_LC_1_30_3  (
            .in0(N__13050),
            .in1(N__12348),
            .in2(N__14132),
            .in3(N__12963),
            .lcout(r_Clock_Count_8_adj_1994),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37554),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i124_LC_2_16_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i124_LC_2_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i124_LC_2_16_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i124_LC_2_16_3  (
            .in0(N__35976),
            .in1(N__14320),
            .in2(_gnd_net_),
            .in3(N__15200),
            .lcout(data_in_15_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37466),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i116_LC_2_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i116_LC_2_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i116_LC_2_17_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i116_LC_2_17_0  (
            .in0(N__35975),
            .in1(N__26353),
            .in2(_gnd_net_),
            .in3(N__14321),
            .lcout(data_in_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37463),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5769_LC_2_17_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5769_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5769_LC_2_17_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5769_LC_2_17_4  (
            .in0(N__27748),
            .in1(N__20619),
            .in2(N__30185),
            .in3(N__14277),
            .lcout(),
            .ltout(\c0.n6135_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6135_bdd_4_lut_LC_2_17_5 .C_ON=1'b0;
    defparam \c0.n6135_bdd_4_lut_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.n6135_bdd_4_lut_LC_2_17_5 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n6135_bdd_4_lut_LC_2_17_5  (
            .in0(N__17223),
            .in1(N__30132),
            .in2(N__12402),
            .in3(N__22966),
            .lcout(),
            .ltout(\c0.n5746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5789_LC_2_17_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5789_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5789_LC_2_17_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5789_LC_2_17_6  (
            .in0(N__13188),
            .in1(N__25406),
            .in2(N__12399),
            .in3(N__25258),
            .lcout(\c0.n6129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5784_LC_2_18_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5784_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5784_LC_2_18_1 .LUT_INIT=16'b1011100011001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5784_LC_2_18_1  (
            .in0(N__14301),
            .in1(N__27747),
            .in2(N__18750),
            .in3(N__30144),
            .lcout(),
            .ltout(\c0.n6153_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6153_bdd_4_lut_LC_2_18_2 .C_ON=1'b0;
    defparam \c0.n6153_bdd_4_lut_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.n6153_bdd_4_lut_LC_2_18_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6153_bdd_4_lut_LC_2_18_2  (
            .in0(N__30145),
            .in1(N__19110),
            .in2(N__12396),
            .in3(N__18471),
            .lcout(),
            .ltout(\c0.n5740_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6129_bdd_4_lut_LC_2_18_3 .C_ON=1'b0;
    defparam \c0.n6129_bdd_4_lut_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6129_bdd_4_lut_LC_2_18_3 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \c0.n6129_bdd_4_lut_LC_2_18_3  (
            .in0(N__13200),
            .in1(N__25403),
            .in2(N__12393),
            .in3(N__12390),
            .lcout(\c0.n6132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i132_LC_2_18_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i132_LC_2_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i132_LC_2_18_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i132_LC_2_18_5  (
            .in0(N__35974),
            .in1(N__21128),
            .in2(_gnd_net_),
            .in3(N__15193),
            .lcout(data_in_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37467),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5709_LC_2_18_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5709_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5709_LC_2_18_6 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5709_LC_2_18_6  (
            .in0(N__27746),
            .in1(N__24365),
            .in2(N__30193),
            .in3(N__28196),
            .lcout(\c0.n6063 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i148_LC_2_18_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i148_LC_2_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i148_LC_2_18_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0___i148_LC_2_18_7  (
            .in0(N__32142),
            .in1(N__12479),
            .in2(N__33273),
            .in3(N__14714),
            .lcout(\c0.data_in_frame_18_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37467),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6063_bdd_4_lut_LC_2_19_0 .C_ON=1'b0;
    defparam \c0.n6063_bdd_4_lut_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.n6063_bdd_4_lut_LC_2_19_0 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n6063_bdd_4_lut_LC_2_19_0  (
            .in0(N__19392),
            .in1(N__29943),
            .in2(N__12447),
            .in3(N__19884),
            .lcout(\c0.n5776 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i54_LC_2_19_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i54_LC_2_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i54_LC_2_19_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_in_0___i54_LC_2_19_2  (
            .in0(N__18488),
            .in1(_gnd_net_),
            .in2(N__21032),
            .in3(N__35942),
            .lcout(data_in_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37470),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6099_bdd_4_lut_LC_2_19_4 .C_ON=1'b0;
    defparam \c0.n6099_bdd_4_lut_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.n6099_bdd_4_lut_LC_2_19_4 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n6099_bdd_4_lut_LC_2_19_4  (
            .in0(N__25386),
            .in1(N__12411),
            .in2(N__13269),
            .in3(N__12432),
            .lcout(\c0.n6102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i62_LC_2_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i62_LC_2_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i62_LC_2_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i62_LC_2_19_5  (
            .in0(N__35941),
            .in1(N__26575),
            .in2(_gnd_net_),
            .in3(N__18487),
            .lcout(data_in_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37470),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n6003_bdd_4_lut_LC_2_19_7 .C_ON=1'b0;
    defparam \c0.tx2.n6003_bdd_4_lut_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n6003_bdd_4_lut_LC_2_19_7 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.tx2.n6003_bdd_4_lut_LC_2_19_7  (
            .in0(N__13542),
            .in1(N__13663),
            .in2(N__13524),
            .in3(N__13605),
            .lcout(\c0.tx2.n6006 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_916_LC_2_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_916_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_916_LC_2_20_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_916_LC_2_20_0  (
            .in0(N__17219),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24605),
            .lcout(),
            .ltout(\c0.n5375_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_2_20_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_2_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_LC_2_20_1  (
            .in0(N__13239),
            .in1(N__13209),
            .in2(N__12414),
            .in3(N__13278),
            .lcout(\c0.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6117_bdd_4_lut_LC_2_20_3 .C_ON=1'b0;
    defparam \c0.n6117_bdd_4_lut_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6117_bdd_4_lut_LC_2_20_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6117_bdd_4_lut_LC_2_20_3  (
            .in0(N__30146),
            .in1(N__25842),
            .in2(N__12666),
            .in3(N__20559),
            .lcout(\c0.n5755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i147_LC_2_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i147_LC_2_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i147_LC_2_20_5 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0___i147_LC_2_20_5  (
            .in0(N__12509),
            .in1(N__33250),
            .in2(N__32235),
            .in3(N__25734),
            .lcout(\c0.data_in_frame_18_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37474),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i80_LC_2_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i80_LC_2_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i80_LC_2_20_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i80_LC_2_20_7  (
            .in0(N__31341),
            .in1(N__32143),
            .in2(N__20925),
            .in3(N__33251),
            .lcout(\c0.data_in_field_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37474),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5719_LC_2_21_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5719_LC_2_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5719_LC_2_21_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5719_LC_2_21_1  (
            .in0(N__27718),
            .in1(N__23340),
            .in2(N__30069),
            .in3(N__14532),
            .lcout(),
            .ltout(\c0.n6075_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6075_bdd_4_lut_LC_2_21_2 .C_ON=1'b0;
    defparam \c0.n6075_bdd_4_lut_LC_2_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.n6075_bdd_4_lut_LC_2_21_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6075_bdd_4_lut_LC_2_21_2  (
            .in0(N__30053),
            .in1(N__17166),
            .in2(N__12462),
            .in3(N__15459),
            .lcout(\c0.n5773 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_866_LC_2_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_866_LC_2_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_866_LC_2_21_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_866_LC_2_21_4  (
            .in0(_gnd_net_),
            .in1(N__20913),
            .in2(_gnd_net_),
            .in3(N__13477),
            .lcout(\c0.n5454 ),
            .ltout(\c0.n5454_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_851_LC_2_21_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_851_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_851_LC_2_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_851_LC_2_21_5  (
            .in0(N__16789),
            .in1(N__26959),
            .in2(N__12453),
            .in3(N__25112),
            .lcout(\c0.n1892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_932_LC_2_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_932_LC_2_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_932_LC_2_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_932_LC_2_21_6  (
            .in0(_gnd_net_),
            .in1(N__19641),
            .in2(_gnd_net_),
            .in3(N__21001),
            .lcout(\c0.n2009 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_811_LC_2_22_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_811_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_811_LC_2_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_811_LC_2_22_0  (
            .in0(N__21447),
            .in1(N__29514),
            .in2(N__14713),
            .in3(N__15512),
            .lcout(),
            .ltout(\c0.n27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_2_22_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_2_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_LC_2_22_1  (
            .in0(N__13494),
            .in1(N__30614),
            .in2(N__12450),
            .in3(N__17284),
            .lcout(\c0.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i25_4_lut_LC_2_22_2 .C_ON=1'b0;
    defparam \c0.i25_4_lut_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i25_4_lut_LC_2_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i25_4_lut_LC_2_22_2  (
            .in0(N__17043),
            .in1(N__20874),
            .in2(N__15858),
            .in3(N__13440),
            .lcout(),
            .ltout(\c0.n52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_812_LC_2_22_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_812_LC_2_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_812_LC_2_22_3 .LUT_INIT=16'b1111111110010110;
    LogicCell40 \c0.i8_4_lut_adj_812_LC_2_22_3  (
            .in0(N__12564),
            .in1(N__21933),
            .in2(N__12558),
            .in3(N__13422),
            .lcout(),
            .ltout(\c0.n24_adj_1879_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_839_LC_2_22_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_839_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_839_LC_2_22_4 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \c0.i12_4_lut_adj_839_LC_2_22_4  (
            .in0(N__12555),
            .in1(N__12549),
            .in2(N__12540),
            .in3(N__13359),
            .lcout(\c0.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i2_LC_2_23_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i2_LC_2_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i2_LC_2_23_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i2_LC_2_23_0  (
            .in0(N__14217),
            .in1(N__13796),
            .in2(N__12492),
            .in3(N__12537),
            .lcout(\c0.tx2.r_Tx_Data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37491),
            .ce(N__13727),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_23_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_23_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_2_23_1  (
            .in0(N__12594),
            .in1(N__12528),
            .in2(N__13664),
            .in3(N__13927),
            .lcout(\c0.tx2.n6045 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5903_LC_2_23_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5903_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5903_LC_2_23_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5903_LC_2_23_2  (
            .in0(N__12513),
            .in1(N__29823),
            .in2(N__13230),
            .in3(N__27635),
            .lcout(),
            .ltout(\c0.n6297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6297_bdd_4_lut_LC_2_23_3 .C_ON=1'b0;
    defparam \c0.n6297_bdd_4_lut_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6297_bdd_4_lut_LC_2_23_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6297_bdd_4_lut_LC_2_23_3  (
            .in0(N__29824),
            .in1(N__15493),
            .in2(N__12495),
            .in3(N__15540),
            .lcout(\c0.n6300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5898_LC_2_23_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5898_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5898_LC_2_23_4 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5898_LC_2_23_4  (
            .in0(N__12483),
            .in1(N__29825),
            .in2(N__27702),
            .in3(N__13505),
            .lcout(),
            .ltout(\c0.n6279_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6279_bdd_4_lut_LC_2_23_5 .C_ON=1'b0;
    defparam \c0.n6279_bdd_4_lut_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.n6279_bdd_4_lut_LC_2_23_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6279_bdd_4_lut_LC_2_23_5  (
            .in0(N__29826),
            .in1(N__16392),
            .in2(N__12465),
            .in3(N__22551),
            .lcout(),
            .ltout(\c0.n6282_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i3_LC_2_23_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i3_LC_2_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i3_LC_2_23_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i3_LC_2_23_6  (
            .in0(N__14218),
            .in1(N__13797),
            .in2(N__12609),
            .in3(N__12606),
            .lcout(\c0.tx2.r_Tx_Data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37491),
            .ce(N__13727),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_940_LC_2_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_940_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_940_LC_2_23_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_940_LC_2_23_7  (
            .in0(_gnd_net_),
            .in1(N__15492),
            .in2(_gnd_net_),
            .in3(N__15539),
            .lcout(\c0.n2056 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i131_LC_2_24_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i131_LC_2_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i131_LC_2_24_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i131_LC_2_24_0  (
            .in0(N__32474),
            .in1(N__32234),
            .in2(N__15508),
            .in3(N__15915),
            .lcout(\c0.data_in_field_130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37501),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5714_LC_2_24_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5714_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5714_LC_2_24_1 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5714_LC_2_24_1  (
            .in0(N__23205),
            .in1(N__27684),
            .in2(N__30148),
            .in3(N__15962),
            .lcout(\c0.n6069 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5864_LC_2_24_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5864_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5864_LC_2_24_2 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5864_LC_2_24_2  (
            .in0(N__27683),
            .in1(N__30055),
            .in2(N__24543),
            .in3(N__18380),
            .lcout(),
            .ltout(\c0.n6249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6249_bdd_4_lut_LC_2_24_3 .C_ON=1'b0;
    defparam \c0.n6249_bdd_4_lut_LC_2_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6249_bdd_4_lut_LC_2_24_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6249_bdd_4_lut_LC_2_24_3  (
            .in0(N__30054),
            .in1(N__30615),
            .in2(N__12579),
            .in3(N__28005),
            .lcout(\c0.n5695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i115_LC_2_24_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i115_LC_2_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i115_LC_2_24_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i115_LC_2_24_6  (
            .in0(N__35501),
            .in1(N__13387),
            .in2(_gnd_net_),
            .in3(N__19301),
            .lcout(data_in_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37501),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i64_LC_2_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i64_LC_2_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i64_LC_2_24_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i64_LC_2_24_7  (
            .in0(N__15611),
            .in1(N__35502),
            .in2(_gnd_net_),
            .in3(N__23249),
            .lcout(data_in_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37501),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3459_4_lut_LC_2_25_0 .C_ON=1'b0;
    defparam \c0.i3459_4_lut_LC_2_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3459_4_lut_LC_2_25_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3459_4_lut_LC_2_25_0  (
            .in0(N__32233),
            .in1(N__12648),
            .in2(N__15378),
            .in3(N__12576),
            .lcout(\c0.n3703 ),
            .ltout(\c0.n3703_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5628_2_lut_LC_2_25_1 .C_ON=1'b0;
    defparam \c0.i5628_2_lut_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5628_2_lut_LC_2_25_1 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \c0.i5628_2_lut_LC_2_25_1  (
            .in0(N__32372),
            .in1(_gnd_net_),
            .in2(N__12567),
            .in3(_gnd_net_),
            .lcout(\c0.n2325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5754_LC_2_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5754_LC_2_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5754_LC_2_25_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5754_LC_2_25_2  (
            .in0(N__27546),
            .in1(N__14598),
            .in2(N__29924),
            .in3(N__24806),
            .lcout(\c0.n6117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_846_LC_2_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_846_LC_2_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_846_LC_2_25_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_846_LC_2_25_3  (
            .in0(_gnd_net_),
            .in1(N__29562),
            .in2(_gnd_net_),
            .in3(N__18381),
            .lcout(\c0.n5536 ),
            .ltout(\c0.n5536_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_827_LC_2_25_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_827_LC_2_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_827_LC_2_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_827_LC_2_25_4  (
            .in0(N__17058),
            .in1(N__14433),
            .in2(N__12654),
            .in3(N__16992),
            .lcout(),
            .ltout(\c0.n5570_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_840_LC_2_25_5 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_840_LC_2_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_840_LC_2_25_5 .LUT_INIT=16'b1111111101101111;
    LogicCell40 \c0.i11_4_lut_adj_840_LC_2_25_5  (
            .in0(N__19356),
            .in1(N__20448),
            .in2(N__12651),
            .in3(N__22380),
            .lcout(\c0.n27_adj_1910 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i489_3_lut_4_lut_LC_2_26_0 .C_ON=1'b0;
    defparam \c0.i489_3_lut_4_lut_LC_2_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i489_3_lut_4_lut_LC_2_26_0 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \c0.i489_3_lut_4_lut_LC_2_26_0  (
            .in0(N__12746),
            .in1(N__12730),
            .in2(N__32437),
            .in3(N__12622),
            .lcout(\c0.n195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3445_2_lut_LC_2_26_2 .C_ON=1'b0;
    defparam \c0.i3445_2_lut_LC_2_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3445_2_lut_LC_2_26_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i3445_2_lut_LC_2_26_2  (
            .in0(N__12745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12729),
            .lcout(\c0.n3689 ),
            .ltout(\c0.n3689_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_2_26_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_2_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_2_26_3 .LUT_INIT=16'b1111101000110011;
    LogicCell40 \c0.FRAME_MATCHER_wait_for_transmission_1803_LC_2_26_3  (
            .in0(N__13591),
            .in1(N__12627),
            .in2(N__12642),
            .in3(N__32379),
            .lcout(\c0.FRAME_MATCHER_wait_for_transmission ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_45_LC_2_26_4 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_45_LC_2_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.o_Tx_Serial_45_LC_2_26_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \c0.tx2.o_Tx_Serial_45_LC_2_26_4  (
            .in0(N__14126),
            .in1(N__12691),
            .in2(_gnd_net_),
            .in3(N__12639),
            .lcout(tx2_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_1801_LC_2_26_6 .C_ON=1'b0;
    defparam \c0.tx2_transmit_1801_LC_2_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2_transmit_1801_LC_2_26_6 .LUT_INIT=16'b0100000001001111;
    LogicCell40 \c0.tx2_transmit_1801_LC_2_26_6  (
            .in0(N__12633),
            .in1(N__13592),
            .in2(N__32438),
            .in3(N__12623),
            .lcout(\c0.r_SM_Main_2_N_1770_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37521),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i895_2_lut_LC_2_26_7 .C_ON=1'b0;
    defparam \c0.tx2.i895_2_lut_LC_2_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i895_2_lut_LC_2_26_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx2.i895_2_lut_LC_2_26_7  (
            .in0(_gnd_net_),
            .in1(N__12782),
            .in2(_gnd_net_),
            .in3(N__13644),
            .lcout(\c0.tx2.n1136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i28_4_lut_LC_2_27_0 .C_ON=1'b0;
    defparam \c0.tx2.i28_4_lut_LC_2_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i28_4_lut_LC_2_27_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.tx2.i28_4_lut_LC_2_27_0  (
            .in0(N__12764),
            .in1(N__12722),
            .in2(N__12894),
            .in3(N__13854),
            .lcout(\c0.tx2.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2088_4_lut_LC_2_27_1 .C_ON=1'b0;
    defparam \c0.tx2.i2088_4_lut_LC_2_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2088_4_lut_LC_2_27_1 .LUT_INIT=16'b1101010100000000;
    LogicCell40 \c0.tx2.i2088_4_lut_LC_2_27_1  (
            .in0(N__12882),
            .in1(N__13914),
            .in2(N__12765),
            .in3(N__13963),
            .lcout(n2339),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5614_4_lut_4_lut_LC_2_27_5 .C_ON=1'b0;
    defparam \c0.tx2.i5614_4_lut_4_lut_LC_2_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5614_4_lut_4_lut_LC_2_27_5 .LUT_INIT=16'b1001100000010000;
    LogicCell40 \c0.tx2.i5614_4_lut_4_lut_LC_2_27_5  (
            .in0(N__12883),
            .in1(N__14011),
            .in2(N__12731),
            .in3(N__13879),
            .lcout(),
            .ltout(n4_adj_1973_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_47_LC_2_27_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_47_LC_2_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_47_LC_2_27_6 .LUT_INIT=16'b1000110011011100;
    LogicCell40 \c0.tx2.r_Tx_Active_47_LC_2_27_6  (
            .in0(N__14100),
            .in1(N__12747),
            .in2(N__12750),
            .in3(N__12884),
            .lcout(tx2_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37533),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_3_lut_4_lut_LC_2_27_7 .C_ON=1'b0;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_2_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_2_27_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx2.i2_3_lut_4_lut_LC_2_27_7  (
            .in0(N__12881),
            .in1(N__14099),
            .in2(N__12732),
            .in3(N__14012),
            .lcout(\c0.tx2.n1624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_28_0 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_28_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_2_28_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12704),
            .lcout(tx2_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_2_28_1 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_2_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_2_28_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_2_28_1  (
            .in0(N__16305),
            .in1(N__17695),
            .in2(N__18023),
            .in3(N__17645),
            .lcout(r_SM_Main_2_adj_1989),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37544),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i1_LC_2_28_3 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_28_3 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \c0.tx2.r_SM_Main_i1_LC_2_28_3  (
            .in0(N__14115),
            .in1(N__14007),
            .in2(N__12892),
            .in3(N__13880),
            .lcout(r_SM_Main_1_adj_1993),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37544),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i3_4_lut_adj_799_LC_2_28_4 .C_ON=1'b0;
    defparam \c0.tx2.i3_4_lut_adj_799_LC_2_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i3_4_lut_adj_799_LC_2_28_4 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \c0.tx2.i3_4_lut_adj_799_LC_2_28_4  (
            .in0(N__12876),
            .in1(N__12912),
            .in2(N__14017),
            .in3(N__13116),
            .lcout(\c0.tx2.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i7_4_lut_LC_2_28_5 .C_ON=1'b0;
    defparam \c0.tx2.i7_4_lut_LC_2_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i7_4_lut_LC_2_28_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx2.i7_4_lut_LC_2_28_5  (
            .in0(N__12977),
            .in1(N__13092),
            .in2(N__12920),
            .in3(N__13001),
            .lcout(\c0.tx2.r_SM_Main_2_N_1767_1 ),
            .ltout(\c0.tx2.r_SM_Main_2_N_1767_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_4_lut_LC_2_28_6 .C_ON=1'b0;
    defparam \c0.tx2.i2_4_lut_LC_2_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_4_lut_LC_2_28_6 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \c0.tx2.i2_4_lut_LC_2_28_6  (
            .in0(N__14006),
            .in1(N__12877),
            .in2(N__12837),
            .in3(N__14114),
            .lcout(n2208),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_793_LC_2_28_7 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_793_LC_2_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_793_LC_2_28_7 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \c0.rx.i1_4_lut_adj_793_LC_2_28_7  (
            .in0(N__13848),
            .in1(N__16286),
            .in2(N__18022),
            .in3(N__20300),
            .lcout(\c0.rx.n359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i6_LC_2_29_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i6_LC_2_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i6_LC_2_29_0 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i6_LC_2_29_0  (
            .in0(N__12834),
            .in1(N__12961),
            .in2(N__13032),
            .in3(N__14125),
            .lcout(\c0.tx2.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i0_LC_2_29_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i0_LC_2_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i0_LC_2_29_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx2.r_Clock_Count__i0_LC_2_29_1  (
            .in0(N__13175),
            .in1(N__12828),
            .in2(_gnd_net_),
            .in3(N__14111),
            .lcout(\c0.tx2.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_29_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_29_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx2.r_Clock_Count__i1_LC_2_29_2  (
            .in0(N__12822),
            .in1(N__14123),
            .in2(_gnd_net_),
            .in3(N__13160),
            .lcout(\c0.tx2.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i7_LC_2_29_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i7_LC_2_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i7_LC_2_29_3 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i7_LC_2_29_3  (
            .in0(N__12960),
            .in1(N__12816),
            .in2(N__13074),
            .in3(N__14113),
            .lcout(\c0.tx2.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i2_LC_2_29_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i2_LC_2_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i2_LC_2_29_4 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i2_LC_2_29_4  (
            .in0(N__12797),
            .in1(N__12962),
            .in2(N__12807),
            .in3(N__14124),
            .lcout(\c0.tx2.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i85_2_lut_LC_2_29_5 .C_ON=1'b0;
    defparam \c0.tx2.i85_2_lut_LC_2_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i85_2_lut_LC_2_29_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx2.i85_2_lut_LC_2_29_5  (
            .in0(_gnd_net_),
            .in1(N__12796),
            .in2(_gnd_net_),
            .in3(N__13135),
            .lcout(\c0.tx2.n78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_2_lut_LC_2_29_6 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_LC_2_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_LC_2_29_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx2.i1_2_lut_LC_2_29_6  (
            .in0(_gnd_net_),
            .in1(N__13174),
            .in2(_gnd_net_),
            .in3(N__13159),
            .lcout(\c0.tx2.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i5_LC_2_29_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i5_LC_2_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i5_LC_2_29_7 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i5_LC_2_29_7  (
            .in0(N__12959),
            .in1(N__13146),
            .in2(N__13140),
            .in3(N__14112),
            .lcout(\c0.tx2.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37555),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i6_4_lut_LC_2_30_2 .C_ON=1'b0;
    defparam \c0.tx2.i6_4_lut_LC_2_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i6_4_lut_LC_2_30_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx2.i6_4_lut_LC_2_30_2  (
            .in0(N__13068),
            .in1(N__13119),
            .in2(N__13030),
            .in3(N__13047),
            .lcout(\c0.tx2.n14_adj_1867 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_2_30_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_2_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_2_30_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_2_30_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13083),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37564),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5285_4_lut_LC_2_30_6 .C_ON=1'b0;
    defparam \c0.tx2.i5285_4_lut_LC_2_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5285_4_lut_LC_2_30_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx2.i5285_4_lut_LC_2_30_6  (
            .in0(N__13069),
            .in1(N__13048),
            .in2(N__13031),
            .in3(N__13002),
            .lcout(),
            .ltout(\c0.tx2.n5631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_adj_800_LC_2_30_7 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_adj_800_LC_2_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_adj_800_LC_2_30_7 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \c0.tx2.i1_4_lut_adj_800_LC_2_30_7  (
            .in0(N__14119),
            .in1(N__12990),
            .in2(N__12981),
            .in3(N__12978),
            .lcout(n4544),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i44_LC_3_16_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i44_LC_3_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i44_LC_3_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i44_LC_3_16_1  (
            .in0(N__35943),
            .in1(N__16469),
            .in2(_gnd_net_),
            .in3(N__16694),
            .lcout(data_in_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37471),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i60_LC_3_16_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i60_LC_3_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i60_LC_3_16_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i60_LC_3_16_2  (
            .in0(N__32063),
            .in1(N__33138),
            .in2(N__14247),
            .in3(N__14297),
            .lcout(\c0.data_in_field_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37471),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i60_LC_3_16_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i60_LC_3_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i60_LC_3_16_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i60_LC_3_16_3  (
            .in0(N__35944),
            .in1(N__14242),
            .in2(_gnd_net_),
            .in3(N__14390),
            .lcout(data_in_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37471),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5794_LC_3_16_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5794_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5794_LC_3_16_5 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5794_LC_3_16_5  (
            .in0(N__27749),
            .in1(N__18609),
            .in2(N__30208),
            .in3(N__22593),
            .lcout(),
            .ltout(\c0.n6159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6159_bdd_4_lut_LC_3_16_6 .C_ON=1'b0;
    defparam \c0.n6159_bdd_4_lut_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.n6159_bdd_4_lut_LC_3_16_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6159_bdd_4_lut_LC_3_16_6  (
            .in0(N__30186),
            .in1(N__18654),
            .in2(N__13203),
            .in3(N__14414),
            .lcout(\c0.n5737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6141_bdd_4_lut_LC_3_16_7 .C_ON=1'b0;
    defparam \c0.n6141_bdd_4_lut_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.n6141_bdd_4_lut_LC_3_16_7 .LUT_INIT=16'b1010110110101000;
    LogicCell40 \c0.n6141_bdd_4_lut_LC_3_16_7  (
            .in0(N__13182),
            .in1(N__19026),
            .in2(N__30207),
            .in3(N__14365),
            .lcout(\c0.n5743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5774_LC_3_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5774_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5774_LC_3_17_0 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5774_LC_3_17_0  (
            .in0(N__27608),
            .in1(N__18572),
            .in2(N__30059),
            .in3(N__27957),
            .lcout(\c0.n6141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_850_LC_3_17_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_850_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_850_LC_3_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_850_LC_3_17_1  (
            .in0(N__18466),
            .in1(N__14773),
            .in2(_gnd_net_),
            .in3(N__14364),
            .lcout(\c0.n2095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i24_LC_3_17_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i24_LC_3_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i24_LC_3_17_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i24_LC_3_17_2  (
            .in0(N__16416),
            .in1(N__18194),
            .in2(_gnd_net_),
            .in3(N__35939),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37465),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i120_LC_3_17_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i120_LC_3_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i120_LC_3_17_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i120_LC_3_17_3  (
            .in0(N__21872),
            .in1(_gnd_net_),
            .in2(N__36023),
            .in3(N__13252),
            .lcout(data_in_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37465),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i120_LC_3_17_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i120_LC_3_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i120_LC_3_17_4 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i120_LC_3_17_4  (
            .in0(N__14774),
            .in1(N__33026),
            .in2(N__13259),
            .in3(N__31850),
            .lcout(\c0.data_in_field_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37465),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i104_LC_3_17_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i104_LC_3_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i104_LC_3_17_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i104_LC_3_17_5  (
            .in0(N__35935),
            .in1(N__13346),
            .in2(_gnd_net_),
            .in3(N__18841),
            .lcout(data_in_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37465),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i68_LC_3_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i68_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i68_LC_3_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i68_LC_3_18_0  (
            .in0(N__35933),
            .in1(N__18671),
            .in2(_gnd_net_),
            .in3(N__14383),
            .lcout(data_in_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37472),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5764_LC_3_18_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5764_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5764_LC_3_18_2 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5764_LC_3_18_2  (
            .in0(N__27753),
            .in1(N__23025),
            .in2(N__30060),
            .in3(N__16827),
            .lcout(),
            .ltout(\c0.n6123_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6123_bdd_4_lut_LC_3_18_3 .C_ON=1'b0;
    defparam \c0.n6123_bdd_4_lut_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6123_bdd_4_lut_LC_3_18_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6123_bdd_4_lut_LC_3_18_3  (
            .in0(N__30147),
            .in1(N__27261),
            .in2(N__13272),
            .in3(N__16905),
            .lcout(\c0.n5752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i112_LC_3_18_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i112_LC_3_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i112_LC_3_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i112_LC_3_18_4  (
            .in0(N__35932),
            .in1(N__13260),
            .in2(_gnd_net_),
            .in3(N__13339),
            .lcout(data_in_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37472),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_adj_983_LC_3_18_5 .C_ON=1'b0;
    defparam \c0.i7_3_lut_adj_983_LC_3_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_adj_983_LC_3_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i7_3_lut_adj_983_LC_3_18_5  (
            .in0(N__28195),
            .in1(N__24119),
            .in2(_gnd_net_),
            .in3(N__22968),
            .lcout(\c0.n24_adj_1877 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i84_LC_3_18_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i84_LC_3_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i84_LC_3_18_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i84_LC_3_18_7  (
            .in0(N__16944),
            .in1(N__35934),
            .in2(_gnd_net_),
            .in3(N__14464),
            .lcout(data_in_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37472),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i140_LC_3_19_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i140_LC_3_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i140_LC_3_19_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i140_LC_3_19_0  (
            .in0(N__35681),
            .in1(N__21127),
            .in2(_gnd_net_),
            .in3(N__14715),
            .lcout(data_in_17_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37475),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i155_LC_3_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i155_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i155_LC_3_19_2 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i155_LC_3_19_2  (
            .in0(N__32071),
            .in1(N__13223),
            .in2(N__25908),
            .in3(N__32978),
            .lcout(\c0.data_in_frame_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37475),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_854_LC_3_19_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_854_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_854_LC_3_19_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_854_LC_3_19_4  (
            .in0(N__20614),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27097),
            .lcout(\c0.n5381 ),
            .ltout(\c0.n5381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_3_19_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_3_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_LC_3_19_5  (
            .in0(N__20679),
            .in1(N__15777),
            .in2(N__13353),
            .in3(N__16381),
            .lcout(\c0.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_902_LC_3_19_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_902_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_902_LC_3_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_902_LC_3_19_6  (
            .in0(N__15267),
            .in1(N__24870),
            .in2(N__28311),
            .in3(N__26799),
            .lcout(\c0.n18_adj_1938 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i112_LC_3_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i112_LC_3_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i112_LC_3_19_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i112_LC_3_19_7  (
            .in0(N__32977),
            .in1(N__32072),
            .in2(N__13350),
            .in3(N__14753),
            .lcout(\c0.data_in_field_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37475),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_3_20_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_3_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_LC_3_20_0  (
            .in0(N__20171),
            .in1(N__13323),
            .in2(N__24355),
            .in3(N__27042),
            .lcout(\c0.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i82_LC_3_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i82_LC_3_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i82_LC_3_20_1 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i82_LC_3_20_1  (
            .in0(N__32064),
            .in1(N__17844),
            .in2(N__32778),
            .in3(N__14531),
            .lcout(\c0.data_in_field_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37479),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i135_LC_3_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i135_LC_3_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i135_LC_3_20_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i135_LC_3_20_2  (
            .in0(N__17031),
            .in1(N__13317),
            .in2(N__32217),
            .in3(N__32598),
            .lcout(\c0.data_in_field_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37479),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i96_LC_3_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i96_LC_3_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i96_LC_3_20_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i96_LC_3_20_3  (
            .in0(N__20843),
            .in1(N__26163),
            .in2(N__32779),
            .in3(N__32076),
            .lcout(\c0.data_in_field_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37479),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_921_LC_3_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_921_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_921_LC_3_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_921_LC_3_20_5  (
            .in0(N__20842),
            .in1(N__20811),
            .in2(_gnd_net_),
            .in3(N__14530),
            .lcout(\c0.n1942 ),
            .ltout(\c0.n1942_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_920_LC_3_20_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_920_LC_3_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_920_LC_3_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_920_LC_3_20_6  (
            .in0(N__25148),
            .in1(N__18577),
            .in2(N__13290),
            .in3(N__19879),
            .lcout(\c0.n5578 ),
            .ltout(\c0.n5578_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_984_LC_3_20_7 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_984_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_984_LC_3_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_984_LC_3_20_7  (
            .in0(N__13287),
            .in1(N__17106),
            .in2(N__13281),
            .in3(N__20892),
            .lcout(\c0.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_972_LC_3_21_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_972_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_972_LC_3_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_972_LC_3_21_0  (
            .in0(N__23238),
            .in1(N__25517),
            .in2(N__15351),
            .in3(N__13404),
            .lcout(\c0.n5488 ),
            .ltout(\c0.n5488_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_2_lut_3_lut_LC_3_21_1 .C_ON=1'b0;
    defparam \c0.i9_2_lut_3_lut_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_2_lut_3_lut_LC_3_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i9_2_lut_3_lut_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(N__14418),
            .in2(N__13446),
            .in3(N__16391),
            .lcout(),
            .ltout(\c0.n36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_3_21_2 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_3_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_LC_3_21_2  (
            .in0(N__24263),
            .in1(N__15840),
            .in2(N__13443),
            .in3(N__21769),
            .lcout(\c0.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_810_LC_3_21_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_810_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_810_LC_3_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_810_LC_3_21_3  (
            .in0(N__13434),
            .in1(N__13416),
            .in2(N__15165),
            .in3(N__13428),
            .lcout(\c0.n5489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_909_LC_3_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_909_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_909_LC_3_21_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_909_LC_3_21_5  (
            .in0(_gnd_net_),
            .in1(N__18578),
            .in2(_gnd_net_),
            .in3(N__19880),
            .lcout(\c0.n1886 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_970_LC_3_21_6 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_970_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_970_LC_3_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_970_LC_3_21_6  (
            .in0(N__13410),
            .in1(N__16967),
            .in2(N__15762),
            .in3(N__14486),
            .lcout(\c0.n12_adj_1951 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i115_LC_3_22_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i115_LC_3_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i115_LC_3_22_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i115_LC_3_22_0  (
            .in0(N__32982),
            .in1(N__32067),
            .in2(N__13398),
            .in3(N__17086),
            .lcout(\c0.data_in_field_114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37492),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_3_22_1 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_3_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_3_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_LC_3_22_1  (
            .in0(N__13371),
            .in1(N__15630),
            .in2(N__14637),
            .in3(N__14538),
            .lcout(\c0.n5586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i156_LC_3_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i156_LC_3_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i156_LC_3_22_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i156_LC_3_22_3  (
            .in0(N__32065),
            .in1(N__15747),
            .in2(N__13509),
            .in3(N__32985),
            .lcout(\c0.data_in_frame_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37492),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i72_LC_3_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i72_LC_3_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i72_LC_3_22_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i72_LC_3_22_4  (
            .in0(N__36024),
            .in1(N__31337),
            .in2(_gnd_net_),
            .in3(N__15598),
            .lcout(data_in_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37492),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_3_22_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_3_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_LC_3_22_5  (
            .in0(N__16904),
            .in1(N__18431),
            .in2(_gnd_net_),
            .in3(N__18743),
            .lcout(\c0.n22_adj_1876 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i139_LC_3_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i139_LC_3_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i139_LC_3_22_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i139_LC_3_22_6  (
            .in0(N__32983),
            .in1(N__32068),
            .in2(N__15551),
            .in3(N__25695),
            .lcout(\c0.data_in_field_138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37492),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i50_LC_3_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i50_LC_3_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i50_LC_3_22_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i50_LC_3_22_7  (
            .in0(N__32066),
            .in1(N__32984),
            .in2(N__22484),
            .in3(N__13481),
            .lcout(\c0.data_in_field_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37492),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5652_LC_3_23_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5652_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5652_LC_3_23_0 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5652_LC_3_23_0  (
            .in0(N__28130),
            .in1(N__27647),
            .in2(N__20859),
            .in3(N__29802),
            .lcout(),
            .ltout(\c0.n5991_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5991_bdd_4_lut_LC_3_23_1 .C_ON=1'b0;
    defparam \c0.n5991_bdd_4_lut_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.n5991_bdd_4_lut_LC_3_23_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n5991_bdd_4_lut_LC_3_23_1  (
            .in0(N__29803),
            .in1(N__30779),
            .in2(N__13461),
            .in3(N__20924),
            .lcout(\c0.n5994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i119_LC_3_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i119_LC_3_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i119_LC_3_23_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i119_LC_3_23_2  (
            .in0(N__32756),
            .in1(N__19818),
            .in2(N__18791),
            .in3(N__32070),
            .lcout(\c0.data_in_field_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5744_LC_3_23_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5744_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5744_LC_3_23_3 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5744_LC_3_23_3  (
            .in0(N__27646),
            .in1(N__17085),
            .in2(N__29938),
            .in3(N__24606),
            .lcout(\c0.n6105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i79_LC_3_23_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i79_LC_3_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i79_LC_3_23_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i79_LC_3_23_4  (
            .in0(N__36043),
            .in1(N__31183),
            .in2(_gnd_net_),
            .in3(N__17474),
            .lcout(data_in_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i96_LC_3_23_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i96_LC_3_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i96_LC_3_23_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i96_LC_3_23_5  (
            .in0(N__26158),
            .in1(N__36044),
            .in2(_gnd_net_),
            .in3(N__18854),
            .lcout(data_in_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i150_LC_3_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i150_LC_3_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i150_LC_3_23_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i150_LC_3_23_7  (
            .in0(N__32069),
            .in1(N__13560),
            .in2(N__21399),
            .in3(N__32757),
            .lcout(\c0.data_in_frame_18_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37502),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5849_LC_3_24_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5849_LC_3_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5849_LC_3_24_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5849_LC_3_24_0  (
            .in0(N__27633),
            .in1(N__19839),
            .in2(N__30126),
            .in3(N__13559),
            .lcout(),
            .ltout(\c0.n6225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6225_bdd_4_lut_LC_3_24_1 .C_ON=1'b0;
    defparam \c0.n6225_bdd_4_lut_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.n6225_bdd_4_lut_LC_3_24_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n6225_bdd_4_lut_LC_3_24_1  (
            .in0(N__20175),
            .in1(N__30025),
            .in2(N__13548),
            .in3(N__27168),
            .lcout(),
            .ltout(\c0.n6228_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i5_LC_3_24_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i5_LC_3_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i5_LC_3_24_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i5_LC_3_24_2  (
            .in0(N__14220),
            .in1(N__13789),
            .in2(N__13545),
            .in3(N__23589),
            .lcout(\c0.tx2.r_Tx_Data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37510),
            .ce(N__13737),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5879_LC_3_24_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5879_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5879_LC_3_24_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5879_LC_3_24_4  (
            .in0(N__27634),
            .in1(N__17544),
            .in2(N__30127),
            .in3(N__14829),
            .lcout(),
            .ltout(\c0.n6267_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6267_bdd_4_lut_LC_3_24_5 .C_ON=1'b0;
    defparam \c0.n6267_bdd_4_lut_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n6267_bdd_4_lut_LC_3_24_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6267_bdd_4_lut_LC_3_24_5  (
            .in0(N__29827),
            .in1(N__20742),
            .in2(N__13530),
            .in3(N__18888),
            .lcout(),
            .ltout(\c0.n6270_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i4_LC_3_24_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i4_LC_3_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i4_LC_3_24_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \c0.tx2.r_Tx_Data_i4_LC_3_24_6  (
            .in0(N__14219),
            .in1(N__13788),
            .in2(N__13527),
            .in3(N__14649),
            .lcout(\c0.tx2.r_Tx_Data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37510),
            .ce(N__13737),
            .sr(_gnd_net_));
    defparam \c0.i5622_4_lut_LC_3_24_7 .C_ON=1'b0;
    defparam \c0.i5622_4_lut_LC_3_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5622_4_lut_LC_3_24_7 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \c0.i5622_4_lut_LC_3_24_7  (
            .in0(N__13787),
            .in1(N__30018),
            .in2(N__14221),
            .in3(N__27632),
            .lcout(\c0.FRAME_MATCHER_wait_for_transmission_N_909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5724_LC_3_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5724_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5724_LC_3_25_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5724_LC_3_25_0  (
            .in0(N__16095),
            .in1(N__29782),
            .in2(N__19752),
            .in3(N__27557),
            .lcout(\c0.n6081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i7_LC_3_25_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i7_LC_3_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i7_LC_3_25_2 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \c0.tx2.r_Tx_Data_i7_LC_3_25_2  (
            .in0(N__13827),
            .in1(N__14207),
            .in2(N__13803),
            .in3(N__14721),
            .lcout(\c0.tx2.r_Tx_Data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(N__13732),
            .sr(_gnd_net_));
    defparam \c0.n6231_bdd_4_lut_LC_3_25_3 .C_ON=1'b0;
    defparam \c0.n6231_bdd_4_lut_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6231_bdd_4_lut_LC_3_25_3 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n6231_bdd_4_lut_LC_3_25_3  (
            .in0(N__13812),
            .in1(N__25306),
            .in2(N__14790),
            .in3(N__17523),
            .lcout(),
            .ltout(\c0.n6234_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i6_LC_3_25_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i6_LC_3_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i6_LC_3_25_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.tx2.r_Tx_Data_i6_LC_3_25_4  (
            .in0(N__14847),
            .in1(N__14206),
            .in2(N__13806),
            .in3(N__13802),
            .lcout(\c0.tx2.r_Tx_Data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37522),
            .ce(N__13732),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_5690_LC_3_25_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_5690_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_5690_LC_3_25_5 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_5690_LC_3_25_5  (
            .in0(N__13680),
            .in1(N__13674),
            .in2(N__13668),
            .in3(N__13918),
            .lcout(\c0.tx2.n6003 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_525_526__i1_LC_3_26_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_525_526__i1_LC_3_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i1_LC_3_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i1_LC_3_26_0  (
            .in0(_gnd_net_),
            .in1(N__27568),
            .in2(N__13593),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter2_0 ),
            .ltout(),
            .carryin(bfn_3_26_0_),
            .carryout(\c0.n4735 ),
            .clk(N__37534),
            .ce(N__14157),
            .sr(N__14148));
    defparam \c0.byte_transmit_counter2_525_526__i2_LC_3_26_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_525_526__i2_LC_3_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i2_LC_3_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i2_LC_3_26_1  (
            .in0(_gnd_net_),
            .in1(N__29792),
            .in2(_gnd_net_),
            .in3(N__13569),
            .lcout(\c0.byte_transmit_counter2_1 ),
            .ltout(),
            .carryin(\c0.n4735 ),
            .carryout(\c0.n4736 ),
            .clk(N__37534),
            .ce(N__14157),
            .sr(N__14148));
    defparam \c0.byte_transmit_counter2_525_526__i3_LC_3_26_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_525_526__i3_LC_3_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i3_LC_3_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i3_LC_3_26_2  (
            .in0(_gnd_net_),
            .in1(N__25238),
            .in2(_gnd_net_),
            .in3(N__13566),
            .lcout(\c0.byte_transmit_counter2_2 ),
            .ltout(),
            .carryin(\c0.n4736 ),
            .carryout(\c0.n4737 ),
            .clk(N__37534),
            .ce(N__14157),
            .sr(N__14148));
    defparam \c0.byte_transmit_counter2_525_526__i4_LC_3_26_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_525_526__i4_LC_3_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i4_LC_3_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i4_LC_3_26_3  (
            .in0(_gnd_net_),
            .in1(N__25305),
            .in2(_gnd_net_),
            .in3(N__13563),
            .lcout(\c0.byte_transmit_counter2_3 ),
            .ltout(),
            .carryin(\c0.n4737 ),
            .carryout(\c0.n4738 ),
            .clk(N__37534),
            .ce(N__14157),
            .sr(N__14148));
    defparam \c0.byte_transmit_counter2_525_526__i5_LC_3_26_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_525_526__i5_LC_3_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_525_526__i5_LC_3_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_525_526__i5_LC_3_26_4  (
            .in0(_gnd_net_),
            .in1(N__14205),
            .in2(_gnd_net_),
            .in3(N__14229),
            .lcout(\c0.byte_transmit_counter2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37534),
            .ce(N__14157),
            .sr(N__14148));
    defparam \c0.tx2.r_SM_Main_i0_LC_3_27_0 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i0_LC_3_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i0_LC_3_27_0 .LUT_INIT=16'b0000011100000010;
    LogicCell40 \c0.tx2.r_SM_Main_i0_LC_3_27_0  (
            .in0(N__14016),
            .in1(N__13878),
            .in2(N__14136),
            .in3(N__14031),
            .lcout(\c0.tx2.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37545),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i0_LC_3_27_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i0_LC_3_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i0_LC_3_27_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \c0.tx2.r_Bit_Index_i0_LC_3_27_1  (
            .in0(N__13913),
            .in1(N__13964),
            .in2(_gnd_net_),
            .in3(N__13940),
            .lcout(r_Bit_Index_0_adj_1995),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37545),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i1_LC_3_27_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i1_LC_3_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_3_27_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_3_27_3  (
            .in0(N__16208),
            .in1(N__14997),
            .in2(_gnd_net_),
            .in3(N__14880),
            .lcout(\c0.rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37545),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5567_2_lut_LC_3_27_4 .C_ON=1'b0;
    defparam \c0.tx2.i5567_2_lut_LC_3_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5567_2_lut_LC_3_27_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx2.i5567_2_lut_LC_3_27_4  (
            .in0(_gnd_net_),
            .in1(N__13912),
            .in2(_gnd_net_),
            .in3(N__13877),
            .lcout(\c0.tx2.n5847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i3_LC_3_27_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i3_LC_3_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_3_27_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_3_27_5  (
            .in0(N__16209),
            .in1(N__14868),
            .in2(_gnd_net_),
            .in3(N__15069),
            .lcout(\c0.rx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37545),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i16_4_lut_LC_3_27_7 .C_ON=1'b0;
    defparam \c0.rx.i16_4_lut_LC_3_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i16_4_lut_LC_3_27_7 .LUT_INIT=16'b1011101010111111;
    LogicCell40 \c0.rx.i16_4_lut_LC_3_27_7  (
            .in0(N__16293),
            .in1(N__17630),
            .in2(N__18024),
            .in3(N__14334),
            .lcout(\c0.rx.n36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5570_2_lut_3_lut_LC_3_28_1 .C_ON=1'b0;
    defparam \c0.rx.i5570_2_lut_3_lut_LC_3_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5570_2_lut_3_lut_LC_3_28_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.rx.i5570_2_lut_3_lut_LC_3_28_1  (
            .in0(N__15014),
            .in1(N__14994),
            .in2(_gnd_net_),
            .in3(N__14955),
            .lcout(\c0.rx.n5823 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_4_lut_adj_794_LC_3_28_4 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_4_lut_adj_794_LC_3_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_4_lut_adj_794_LC_3_28_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \c0.rx.i1_2_lut_4_lut_adj_794_LC_3_28_4  (
            .in0(N__14993),
            .in1(N__14953),
            .in2(N__17697),
            .in3(N__15015),
            .lcout(\c0.rx.n3589 ),
            .ltout(\c0.rx.n3589_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5560_2_lut_LC_3_28_5 .C_ON=1'b0;
    defparam \c0.rx.i5560_2_lut_LC_3_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5560_2_lut_LC_3_28_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \c0.rx.i5560_2_lut_LC_3_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14340),
            .in3(N__20299),
            .lcout(\c0.rx.n5815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_4_lut_LC_3_28_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_4_lut_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_4_lut_LC_3_28_6 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \c0.rx.i1_2_lut_4_lut_LC_3_28_6  (
            .in0(N__14992),
            .in1(N__14952),
            .in2(N__20316),
            .in3(N__15012),
            .lcout(),
            .ltout(\c0.rx.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5574_4_lut_LC_3_28_7 .C_ON=1'b0;
    defparam \c0.rx.i5574_4_lut_LC_3_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5574_4_lut_LC_3_28_7 .LUT_INIT=16'b0111001100110011;
    LogicCell40 \c0.rx.i5574_4_lut_LC_3_28_7  (
            .in0(N__15013),
            .in1(N__17691),
            .in2(N__14337),
            .in3(N__15087),
            .lcout(\c0.rx.n5817 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i59_LC_4_15_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i59_LC_4_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i59_LC_4_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i59_LC_4_15_6  (
            .in0(N__35641),
            .in1(N__14614),
            .in2(_gnd_net_),
            .in3(N__16736),
            .lcout(data_in_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37480),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i124_LC_4_15_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i124_LC_4_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i124_LC_4_15_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i124_LC_4_15_7  (
            .in0(N__33077),
            .in1(N__32125),
            .in2(N__14328),
            .in3(N__14271),
            .lcout(\c0.data_in_field_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37480),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i51_LC_4_16_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i51_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i51_LC_4_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i51_LC_4_16_1  (
            .in0(N__36070),
            .in1(N__14621),
            .in2(_gnd_net_),
            .in3(N__25643),
            .lcout(data_in_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37476),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_939_LC_4_16_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_939_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_939_LC_4_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_939_LC_4_16_3  (
            .in0(N__14273),
            .in1(N__14293),
            .in2(_gnd_net_),
            .in3(N__18653),
            .lcout(\c0.n1979 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_980_LC_4_16_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_980_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_980_LC_4_16_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_980_LC_4_16_5  (
            .in0(N__14272),
            .in1(N__14409),
            .in2(N__14367),
            .in3(N__16361),
            .lcout(\c0.n1926 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i52_LC_4_16_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i52_LC_4_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i52_LC_4_16_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i52_LC_4_16_6  (
            .in0(N__14246),
            .in1(N__36071),
            .in2(_gnd_net_),
            .in3(N__16462),
            .lcout(data_in_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37476),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i12_LC_4_16_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i12_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i12_LC_4_16_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i12_LC_4_16_7  (
            .in0(N__16497),
            .in1(N__32124),
            .in2(N__33219),
            .in3(N__14410),
            .lcout(\c0.data_in_field_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37476),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i105_LC_4_17_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i105_LC_4_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i105_LC_4_17_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i105_LC_4_17_0  (
            .in0(N__33174),
            .in1(N__31847),
            .in2(N__14922),
            .in3(N__19671),
            .lcout(\c0.data_in_field_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37468),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i24_LC_4_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i24_LC_4_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i24_LC_4_17_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i24_LC_4_17_1  (
            .in0(N__31845),
            .in1(N__33175),
            .in2(N__16426),
            .in3(N__15266),
            .lcout(\c0.data_in_field_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37468),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6183_bdd_4_lut_LC_4_17_3 .C_ON=1'b0;
    defparam \c0.n6183_bdd_4_lut_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6183_bdd_4_lut_LC_4_17_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6183_bdd_4_lut_LC_4_17_3  (
            .in0(N__30172),
            .in1(N__24897),
            .in2(N__16680),
            .in3(N__19640),
            .lcout(\c0.n5725 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i138_LC_4_17_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i138_LC_4_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i138_LC_4_17_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i138_LC_4_17_4  (
            .in0(N__36069),
            .in1(N__15568),
            .in2(_gnd_net_),
            .in3(N__15148),
            .lcout(data_in_17_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37468),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i76_LC_4_17_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i76_LC_4_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i76_LC_4_17_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i76_LC_4_17_5  (
            .in0(N__35962),
            .in1(N__18670),
            .in2(_gnd_net_),
            .in3(N__14465),
            .lcout(data_in_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37468),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i16_LC_4_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i16_LC_4_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i16_LC_4_17_6 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i16_LC_4_17_6  (
            .in0(N__18133),
            .in1(N__31848),
            .in2(N__33245),
            .in3(N__15315),
            .lcout(\c0.data_in_field_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37468),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i68_LC_4_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i68_LC_4_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i68_LC_4_17_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i68_LC_4_17_7  (
            .in0(N__31846),
            .in1(N__33176),
            .in2(N__14391),
            .in3(N__14366),
            .lcout(\c0.data_in_field_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37468),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i66_LC_4_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i66_LC_4_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i66_LC_4_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i66_LC_4_18_0  (
            .in0(N__35940),
            .in1(N__17820),
            .in2(_gnd_net_),
            .in3(N__16510),
            .lcout(data_in_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i122_LC_4_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i122_LC_4_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i122_LC_4_18_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i122_LC_4_18_1  (
            .in0(N__36064),
            .in1(N__19519),
            .in2(_gnd_net_),
            .in3(N__15815),
            .lcout(data_in_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_883_LC_4_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_883_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_883_LC_4_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_883_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(N__14914),
            .in2(_gnd_net_),
            .in3(N__16641),
            .lcout(\c0.n2143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i26_LC_4_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i26_LC_4_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i26_LC_4_18_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i26_LC_4_18_3  (
            .in0(N__22316),
            .in1(N__32211),
            .in2(N__30828),
            .in3(N__33081),
            .lcout(\c0.data_in_field_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_adj_815_LC_4_18_4 .C_ON=1'b0;
    defparam \c0.i3_2_lut_adj_815_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_adj_815_LC_4_18_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_adj_815_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(N__17212),
            .in2(_gnd_net_),
            .in3(N__16790),
            .lcout(\c0.n16_adj_1880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i84_LC_4_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i84_LC_4_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i84_LC_4_18_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i84_LC_4_18_5  (
            .in0(N__14466),
            .in1(N__32212),
            .in2(N__18579),
            .in3(N__33082),
            .lcout(\c0.data_in_field_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i18_LC_4_18_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i18_LC_4_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i18_LC_4_18_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i18_LC_4_18_6  (
            .in0(N__22317),
            .in1(N__36068),
            .in2(_gnd_net_),
            .in3(N__18279),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i58_LC_4_18_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i58_LC_4_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i58_LC_4_18_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i58_LC_4_18_7  (
            .in0(N__16511),
            .in1(_gnd_net_),
            .in2(N__36075),
            .in3(N__16066),
            .lcout(data_in_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37477),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_915_LC_4_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_915_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_915_LC_4_19_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_915_LC_4_19_0  (
            .in0(N__27285),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27327),
            .lcout(),
            .ltout(\c0.n5412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_816_LC_4_19_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_816_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_816_LC_4_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_816_LC_4_19_1  (
            .in0(N__15276),
            .in1(N__28188),
            .in2(N__14448),
            .in3(N__18430),
            .lcout(),
            .ltout(\c0.n22_adj_1881_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_818_LC_4_19_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_818_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_818_LC_4_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_818_LC_4_19_2  (
            .in0(N__14445),
            .in1(N__24807),
            .in2(N__14436),
            .in3(N__25524),
            .lcout(\c0.n24_adj_1884 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_872_LC_4_19_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_872_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_872_LC_4_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_872_LC_4_19_3  (
            .in0(N__29607),
            .in1(N__14749),
            .in2(_gnd_net_),
            .in3(N__14529),
            .lcout(\c0.n2134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i107_LC_4_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i107_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i107_LC_4_19_4 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i107_LC_4_19_4  (
            .in0(N__27286),
            .in1(N__32868),
            .in2(N__28395),
            .in3(N__32227),
            .lcout(\c0.data_in_field_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37481),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_879_LC_4_19_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_879_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_879_LC_4_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_879_LC_4_19_5  (
            .in0(N__17010),
            .in1(N__27284),
            .in2(_gnd_net_),
            .in3(N__14806),
            .lcout(\c0.n5554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i15_LC_4_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i15_LC_4_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i15_LC_4_19_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i15_LC_4_19_6  (
            .in0(N__14807),
            .in1(N__32869),
            .in2(N__18162),
            .in3(N__32228),
            .lcout(\c0.data_in_field_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37481),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i130_LC_4_19_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i130_LC_4_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i130_LC_4_19_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i130_LC_4_19_7  (
            .in0(N__36072),
            .in1(N__15575),
            .in2(_gnd_net_),
            .in3(N__15808),
            .lcout(data_in_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37481),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_960_LC_4_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_960_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_960_LC_4_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_960_LC_4_20_0  (
            .in0(N__24536),
            .in1(N__22364),
            .in2(_gnd_net_),
            .in3(N__29608),
            .lcout(\c0.n5551 ),
            .ltout(\c0.n5551_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_1007_LC_4_20_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_1007_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_1007_LC_4_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_1007_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(N__24344),
            .in2(N__14496),
            .in3(N__24299),
            .lcout(\c0.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i48_LC_4_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i48_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i48_LC_4_20_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0___i48_LC_4_20_3  (
            .in0(N__32860),
            .in1(N__29612),
            .in2(N__32284),
            .in3(N__27195),
            .lcout(\c0.data_in_field_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37486),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_4_20_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_4_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_4_20_4  (
            .in0(N__22793),
            .in1(N__20523),
            .in2(N__19731),
            .in3(N__14493),
            .lcout(),
            .ltout(\c0.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_836_LC_4_20_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_836_LC_4_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_836_LC_4_20_5 .LUT_INIT=16'b1001011011111111;
    LogicCell40 \c0.i4_4_lut_adj_836_LC_4_20_5  (
            .in0(N__14475),
            .in1(N__21147),
            .in2(N__14469),
            .in3(N__15699),
            .lcout(\c0.n20_adj_1905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i114_LC_4_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i114_LC_4_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i114_LC_4_20_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i114_LC_4_20_6  (
            .in0(N__24345),
            .in1(N__32861),
            .in2(N__19503),
            .in3(N__32226),
            .lcout(\c0.data_in_field_113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37486),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_LC_4_20_7 .C_ON=1'b0;
    defparam \c0.i6_3_lut_LC_4_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_LC_4_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i6_3_lut_LC_4_20_7  (
            .in0(N__14556),
            .in1(N__25463),
            .in2(_gnd_net_),
            .in3(N__28131),
            .lcout(\c0.n18_adj_1904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5804_LC_4_21_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5804_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5804_LC_4_21_0 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5804_LC_4_21_0  (
            .in0(N__19206),
            .in1(N__27667),
            .in2(N__30171),
            .in3(N__29558),
            .lcout(),
            .ltout(\c0.n6177_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6177_bdd_4_lut_LC_4_21_1 .C_ON=1'b0;
    defparam \c0.n6177_bdd_4_lut_LC_4_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.n6177_bdd_4_lut_LC_4_21_1 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n6177_bdd_4_lut_LC_4_21_1  (
            .in0(N__15687),
            .in1(N__17577),
            .in2(N__14547),
            .in3(N__30089),
            .lcout(),
            .ltout(\c0.n5728_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5814_LC_4_21_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5814_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5814_LC_4_21_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5814_LC_4_21_2  (
            .in0(N__25372),
            .in1(N__25248),
            .in2(N__14544),
            .in3(N__21501),
            .lcout(\c0.n6165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_946_LC_4_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_946_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_946_LC_4_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_946_LC_4_21_4  (
            .in0(N__17285),
            .in1(N__25995),
            .in2(N__19209),
            .in3(N__17241),
            .lcout(\c0.n1973 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i58_LC_4_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i58_LC_4_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i58_LC_4_21_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i58_LC_4_21_7  (
            .in0(N__32240),
            .in1(N__32643),
            .in2(N__16080),
            .in3(N__24309),
            .lcout(\c0.data_in_field_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37493),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_LC_4_22_0 .C_ON=1'b0;
    defparam \c0.i3_2_lut_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_LC_4_22_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_LC_4_22_0  (
            .in0(_gnd_net_),
            .in1(N__16131),
            .in2(_gnd_net_),
            .in3(N__15544),
            .lcout(),
            .ltout(\c0.n16_adj_1873_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_4_22_1 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_4_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_LC_4_22_1  (
            .in0(N__15441),
            .in1(N__15882),
            .in2(N__14541),
            .in3(N__17445),
            .lcout(\c0.n24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6165_bdd_4_lut_LC_4_22_2 .C_ON=1'b0;
    defparam \c0.n6165_bdd_4_lut_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.n6165_bdd_4_lut_LC_4_22_2 .LUT_INIT=16'b1111110000001010;
    LogicCell40 \c0.n6165_bdd_4_lut_LC_4_22_2  (
            .in0(N__21717),
            .in1(N__14667),
            .in2(N__25408),
            .in3(N__14658),
            .lcout(\c0.n6168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_LC_4_22_3 .C_ON=1'b0;
    defparam \c0.i2_4_lut_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_LC_4_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_LC_4_22_3  (
            .in0(N__15440),
            .in1(N__30518),
            .in2(N__30882),
            .in3(N__15872),
            .lcout(\c0.n2012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i159_LC_4_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i159_LC_4_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i159_LC_4_22_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0___i159_LC_4_22_5  (
            .in0(N__32201),
            .in1(N__14570),
            .in2(N__32988),
            .in3(N__15983),
            .lcout(\c0.data_in_frame_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37503),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i74_LC_4_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i74_LC_4_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i74_LC_4_22_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i74_LC_4_22_6  (
            .in0(N__17819),
            .in1(N__32202),
            .in2(N__15457),
            .in3(N__32777),
            .lcout(\c0.data_in_field_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37503),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6213_bdd_4_lut_LC_4_22_7 .C_ON=1'b0;
    defparam \c0.n6213_bdd_4_lut_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.n6213_bdd_4_lut_LC_4_22_7 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6213_bdd_4_lut_LC_4_22_7  (
            .in0(N__29939),
            .in1(N__21228),
            .in2(N__15474),
            .in3(N__23237),
            .lcout(\c0.n5710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i86_LC_4_23_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i86_LC_4_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i86_LC_4_23_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i86_LC_4_23_1  (
            .in0(N__32705),
            .in1(N__32219),
            .in2(N__28857),
            .in3(N__25134),
            .lcout(\c0.data_in_field_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37511),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_LC_4_23_2 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_LC_4_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_3_lut_4_lut_LC_4_23_2  (
            .in0(N__28239),
            .in1(N__28349),
            .in2(N__14594),
            .in3(N__16826),
            .lcout(\c0.n20_adj_1878 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i59_LC_4_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i59_LC_4_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i59_LC_4_23_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i59_LC_4_23_3  (
            .in0(N__32704),
            .in1(N__32218),
            .in2(N__14628),
            .in3(N__14590),
            .lcout(\c0.data_in_field_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37511),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1009_LC_4_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1009_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1009_LC_4_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1009_LC_4_23_4  (
            .in0(N__14586),
            .in1(N__28348),
            .in2(N__17087),
            .in3(N__26848),
            .lcout(\c0.n5575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5779_LC_4_23_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5779_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5779_LC_4_23_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5779_LC_4_23_5  (
            .in0(N__16110),
            .in1(N__29970),
            .in2(N__14571),
            .in3(N__27648),
            .lcout(),
            .ltout(\c0.n6147_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6147_bdd_4_lut_LC_4_23_6 .C_ON=1'b0;
    defparam \c0.n6147_bdd_4_lut_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.n6147_bdd_4_lut_LC_4_23_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6147_bdd_4_lut_LC_4_23_6  (
            .in0(N__29971),
            .in1(N__18963),
            .in2(N__14850),
            .in3(N__17026),
            .lcout(\c0.n6150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i157_LC_4_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i157_LC_4_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i157_LC_4_23_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i157_LC_4_23_7  (
            .in0(N__14828),
            .in1(N__20657),
            .in2(N__32916),
            .in3(N__32220),
            .lcout(\c0.data_in_frame_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37511),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5874_LC_4_24_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5874_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5874_LC_4_24_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5874_LC_4_24_1  (
            .in0(N__27666),
            .in1(N__17354),
            .in2(N__30128),
            .in3(N__19281),
            .lcout(),
            .ltout(\c0.n6255_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6255_bdd_4_lut_LC_4_24_2 .C_ON=1'b0;
    defparam \c0.n6255_bdd_4_lut_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.n6255_bdd_4_lut_LC_4_24_2 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6255_bdd_4_lut_LC_4_24_2  (
            .in0(N__29929),
            .in1(N__14814),
            .in2(N__14793),
            .in3(N__16650),
            .lcout(\c0.n5692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5884_LC_4_24_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5884_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5884_LC_4_24_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5884_LC_4_24_4  (
            .in0(N__27665),
            .in1(N__14781),
            .in2(N__30061),
            .in3(N__19473),
            .lcout(),
            .ltout(\c0.n6273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6273_bdd_4_lut_LC_4_24_5 .C_ON=1'b0;
    defparam \c0.n6273_bdd_4_lut_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n6273_bdd_4_lut_LC_4_24_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6273_bdd_4_lut_LC_4_24_5  (
            .in0(N__30029),
            .in1(N__19143),
            .in2(N__14760),
            .in3(N__14757),
            .lcout(),
            .ltout(\c0.n5686_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_4_24_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_4_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_4_24_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_LC_4_24_6  (
            .in0(N__14733),
            .in1(N__25404),
            .in2(N__14727),
            .in3(N__25231),
            .lcout(),
            .ltout(\c0.n6261_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6261_bdd_4_lut_LC_4_24_7 .C_ON=1'b0;
    defparam \c0.n6261_bdd_4_lut_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.n6261_bdd_4_lut_LC_4_24_7 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6261_bdd_4_lut_LC_4_24_7  (
            .in0(N__25405),
            .in1(N__15327),
            .in2(N__14724),
            .in3(N__29580),
            .lcout(\c0.n6264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i148_LC_4_25_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i148_LC_4_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i148_LC_4_25_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i148_LC_4_25_2  (
            .in0(N__15746),
            .in1(N__35384),
            .in2(_gnd_net_),
            .in3(N__14694),
            .lcout(data_in_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37535),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5675_LC_4_25_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5675_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5675_LC_4_25_5 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5675_LC_4_25_5  (
            .in0(N__27607),
            .in1(N__17372),
            .in2(N__29925),
            .in3(N__25572),
            .lcout(),
            .ltout(\c0.n6021_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6021_bdd_4_lut_LC_4_25_6 .C_ON=1'b0;
    defparam \c0.n6021_bdd_4_lut_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.n6021_bdd_4_lut_LC_4_25_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6021_bdd_4_lut_LC_4_25_6  (
            .in0(N__29786),
            .in1(N__14921),
            .in2(N__14898),
            .in3(N__20809),
            .lcout(\c0.n5797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_2_lut_LC_4_27_0 .C_ON=1'b1;
    defparam \c0.rx.add_62_2_lut_LC_4_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_2_lut_LC_4_27_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_2_lut_LC_4_27_0  (
            .in0(N__15122),
            .in1(N__14954),
            .in2(_gnd_net_),
            .in3(N__14883),
            .lcout(\c0.rx.n5855 ),
            .ltout(),
            .carryin(bfn_4_27_0_),
            .carryout(\c0.rx.n4772 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_3_lut_LC_4_27_1 .C_ON=1'b1;
    defparam \c0.rx.add_62_3_lut_LC_4_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_3_lut_LC_4_27_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_3_lut_LC_4_27_1  (
            .in0(N__15108),
            .in1(N__14996),
            .in2(_gnd_net_),
            .in3(N__14874),
            .lcout(\c0.rx.n5860 ),
            .ltout(),
            .carryin(\c0.rx.n4772 ),
            .carryout(\c0.rx.n4773 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_4_lut_LC_4_27_2 .C_ON=1'b1;
    defparam \c0.rx.add_62_4_lut_LC_4_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_4_lut_LC_4_27_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_4_lut_LC_4_27_2  (
            .in0(N__15121),
            .in1(N__16009),
            .in2(_gnd_net_),
            .in3(N__14871),
            .lcout(\c0.rx.n5822 ),
            .ltout(),
            .carryin(\c0.rx.n4773 ),
            .carryout(\c0.rx.n4774 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_5_lut_LC_4_27_3 .C_ON=1'b1;
    defparam \c0.rx.add_62_5_lut_LC_4_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_5_lut_LC_4_27_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_5_lut_LC_4_27_3  (
            .in0(N__15107),
            .in1(N__15068),
            .in2(_gnd_net_),
            .in3(N__14862),
            .lcout(\c0.rx.n5856 ),
            .ltout(),
            .carryin(\c0.rx.n4774 ),
            .carryout(\c0.rx.n4775 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_6_lut_LC_4_27_4 .C_ON=1'b1;
    defparam \c0.rx.add_62_6_lut_LC_4_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_6_lut_LC_4_27_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_6_lut_LC_4_27_4  (
            .in0(N__15120),
            .in1(_gnd_net_),
            .in2(N__15234),
            .in3(N__14859),
            .lcout(\c0.rx.n5857 ),
            .ltout(),
            .carryin(\c0.rx.n4775 ),
            .carryout(\c0.rx.n4776 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_7_lut_LC_4_27_5 .C_ON=1'b1;
    defparam \c0.rx.add_62_7_lut_LC_4_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_7_lut_LC_4_27_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_7_lut_LC_4_27_5  (
            .in0(N__15109),
            .in1(N__15035),
            .in2(_gnd_net_),
            .in3(N__14856),
            .lcout(\c0.rx.n5858 ),
            .ltout(),
            .carryin(\c0.rx.n4776 ),
            .carryout(\c0.rx.n4777 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_8_lut_LC_4_27_6 .C_ON=1'b1;
    defparam \c0.rx.add_62_8_lut_LC_4_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_8_lut_LC_4_27_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_8_lut_LC_4_27_6  (
            .in0(N__15123),
            .in1(N__15051),
            .in2(_gnd_net_),
            .in3(N__14853),
            .lcout(\c0.rx.n5854 ),
            .ltout(),
            .carryin(\c0.rx.n4777 ),
            .carryout(\c0.rx.n4778 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_9_lut_LC_4_27_7 .C_ON=1'b0;
    defparam \c0.rx.add_62_9_lut_LC_4_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_9_lut_LC_4_27_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_9_lut_LC_4_27_7  (
            .in0(N__15110),
            .in1(N__16172),
            .in2(_gnd_net_),
            .in3(N__15090),
            .lcout(\c0.rx.n5859 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_LC_4_28_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_4_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_4_28_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.i1_2_lut_LC_4_28_0  (
            .in0(_gnd_net_),
            .in1(N__14991),
            .in2(_gnd_net_),
            .in3(N__14949),
            .lcout(\c0.rx.n5361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i5_LC_4_28_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i5_LC_4_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_4_28_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_4_28_1  (
            .in0(N__15036),
            .in1(N__16212),
            .in2(_gnd_net_),
            .in3(N__15081),
            .lcout(\c0.rx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i6_LC_4_28_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i6_LC_4_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_4_28_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_4_28_2  (
            .in0(N__15050),
            .in1(_gnd_net_),
            .in2(N__16222),
            .in3(N__15075),
            .lcout(\c0.rx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_3_lut_LC_4_28_3 .C_ON=1'b0;
    defparam \c0.rx.i3_3_lut_LC_4_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_3_lut_LC_4_28_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.rx.i3_3_lut_LC_4_28_3  (
            .in0(N__15067),
            .in1(N__15229),
            .in2(_gnd_net_),
            .in3(N__15049),
            .lcout(),
            .ltout(\c0.rx.n8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5277_4_lut_LC_4_28_4 .C_ON=1'b0;
    defparam \c0.rx.i5277_4_lut_LC_4_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5277_4_lut_LC_4_28_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.rx.i5277_4_lut_LC_4_28_4  (
            .in0(N__15034),
            .in1(N__16011),
            .in2(N__15018),
            .in3(N__16171),
            .lcout(\c0.rx.n1724 ),
            .ltout(\c0.rx.n1724_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_3_lut_LC_4_28_5 .C_ON=1'b0;
    defparam \c0.rx.i1_3_lut_LC_4_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_3_lut_LC_4_28_5 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \c0.rx.i1_3_lut_LC_4_28_5  (
            .in0(N__14950),
            .in1(_gnd_net_),
            .in2(N__15000),
            .in3(N__14995),
            .lcout(r_SM_Main_2_N_1824_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_4_28_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i0_LC_4_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_4_28_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_4_28_6  (
            .in0(N__16210),
            .in1(N__14951),
            .in2(_gnd_net_),
            .in3(N__14961),
            .lcout(\c0.rx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i4_LC_4_28_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i4_LC_4_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_4_28_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_4_28_7  (
            .in0(N__15233),
            .in1(N__15240),
            .in2(_gnd_net_),
            .in3(N__16211),
            .lcout(\c0.rx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37565),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i8_1_lut_LC_4_32_0 .C_ON=1'b0;
    defparam \c0.tx.i8_1_lut_LC_4_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i8_1_lut_LC_4_32_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.i8_1_lut_LC_4_32_0  (
            .in0(N__28883),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i9_LC_5_15_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i9_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i9_LC_5_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i9_LC_5_15_0  (
            .in0(N__35640),
            .in1(N__28437),
            .in2(_gnd_net_),
            .in3(N__18236),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37487),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i156_LC_5_16_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i156_LC_5_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i156_LC_5_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i156_LC_5_16_1  (
            .in0(N__35478),
            .in1(N__15173),
            .in2(_gnd_net_),
            .in3(N__15735),
            .lcout(data_in_19_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37482),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i132_LC_5_16_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i132_LC_5_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i132_LC_5_16_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i132_LC_5_16_2  (
            .in0(N__33246),
            .in1(N__32024),
            .in2(N__15207),
            .in3(N__16371),
            .lcout(\c0.data_in_field_131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37482),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_5_16_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_5_16_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_5_16_4  (
            .in0(N__19443),
            .in1(N__20360),
            .in2(N__15177),
            .in3(N__17769),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37482),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i146_LC_5_16_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i146_LC_5_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i146_LC_5_16_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i146_LC_5_16_5  (
            .in0(N__35477),
            .in1(N__15147),
            .in2(_gnd_net_),
            .in3(N__26726),
            .lcout(data_in_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37482),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i10_LC_5_17_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i10_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i10_LC_5_17_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i10_LC_5_17_1  (
            .in0(N__16335),
            .in1(N__18286),
            .in2(_gnd_net_),
            .in3(N__35450),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37473),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i100_LC_5_17_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i100_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i100_LC_5_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i100_LC_5_17_2  (
            .in0(N__35449),
            .in1(N__26333),
            .in2(_gnd_net_),
            .in3(N__16444),
            .lcout(data_in_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37473),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i122_LC_5_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i122_LC_5_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i122_LC_5_17_3 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i122_LC_5_17_3  (
            .in0(N__28169),
            .in1(N__33006),
            .in2(N__19529),
            .in3(N__31849),
            .lcout(\c0.data_in_field_121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37473),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5670_LC_5_17_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5670_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5670_LC_5_17_4 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5670_LC_5_17_4  (
            .in0(N__27745),
            .in1(N__15265),
            .in2(N__30204),
            .in3(N__30529),
            .lcout(),
            .ltout(\c0.n6009_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6009_bdd_4_lut_LC_5_17_5 .C_ON=1'b0;
    defparam \c0.n6009_bdd_4_lut_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.n6009_bdd_4_lut_LC_5_17_5 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n6009_bdd_4_lut_LC_5_17_5  (
            .in0(N__16598),
            .in1(N__15314),
            .in2(N__15330),
            .in3(N__30170),
            .lcout(\c0.n6012 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i7_LC_5_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i7_LC_5_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i7_LC_5_17_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i7_LC_5_17_6  (
            .in0(N__31915),
            .in1(N__18219),
            .in2(N__33155),
            .in3(N__16645),
            .lcout(\c0.data_in_field_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37473),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_922_LC_5_17_7 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_922_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_922_LC_5_17_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_922_LC_5_17_7  (
            .in0(N__28168),
            .in1(N__15313),
            .in2(N__30967),
            .in3(N__22949),
            .lcout(\c0.n2080 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i69_LC_5_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i69_LC_5_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i69_LC_5_18_0 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i69_LC_5_18_0  (
            .in0(N__33253),
            .in1(N__23457),
            .in2(N__32283),
            .in3(N__15676),
            .lcout(\c0.data_in_field_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37483),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i9_LC_5_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i9_LC_5_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i9_LC_5_18_1 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0___i9_LC_5_18_1  (
            .in0(N__15290),
            .in1(N__33254),
            .in2(N__32282),
            .in3(N__18252),
            .lcout(\c0.data_in_field_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37483),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_953_LC_5_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_953_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_953_LC_5_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_953_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__15675),
            .in2(_gnd_net_),
            .in3(N__15289),
            .lcout(\c0.n2039 ),
            .ltout(\c0.n2039_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_954_LC_5_18_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_954_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_954_LC_5_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_954_LC_5_18_3  (
            .in0(N__15411),
            .in1(N__16587),
            .in2(N__15270),
            .in3(N__15261),
            .lcout(\c0.n5458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i54_LC_5_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i54_LC_5_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i54_LC_5_18_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i54_LC_5_18_4  (
            .in0(N__33252),
            .in1(N__32207),
            .in2(N__21051),
            .in3(N__15412),
            .lcout(\c0.data_in_field_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37483),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_945_LC_5_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_945_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_945_LC_5_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_945_LC_5_18_5  (
            .in0(N__21975),
            .in1(N__15552),
            .in2(N__15516),
            .in3(N__20857),
            .lcout(\c0.n1835 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_989_LC_5_18_6 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_989_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_989_LC_5_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_989_LC_5_18_6  (
            .in0(N__25568),
            .in1(N__24942),
            .in2(N__30821),
            .in3(N__15341),
            .lcout(\c0.n41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5834_LC_5_19_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5834_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5834_LC_5_19_0 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5834_LC_5_19_0  (
            .in0(N__15414),
            .in1(N__27720),
            .in2(N__30153),
            .in3(N__22363),
            .lcout(\c0.n6213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_LC_5_19_1 .C_ON=1'b0;
    defparam \c0.i8_3_lut_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_LC_5_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i8_3_lut_LC_5_19_1  (
            .in0(N__15458),
            .in1(N__15876),
            .in2(_gnd_net_),
            .in3(N__15360),
            .lcout(\c0.n28_adj_1955 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_LC_5_19_2 .C_ON=1'b0;
    defparam \c0.i2_2_lut_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_LC_5_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i2_2_lut_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__24317),
            .in2(_gnd_net_),
            .in3(N__22202),
            .lcout(),
            .ltout(\c0.n14_adj_1957_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1003_LC_5_19_3 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1003_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1003_LC_5_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1003_LC_5_19_3  (
            .in0(N__21391),
            .in1(N__16665),
            .in2(N__15417),
            .in3(N__15413),
            .lcout(),
            .ltout(\c0.n22_adj_1903_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_835_LC_5_19_4 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_835_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_835_LC_5_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_835_LC_5_19_4  (
            .in0(N__15894),
            .in1(N__30735),
            .in2(N__15396),
            .in3(N__15393),
            .lcout(),
            .ltout(\c0.n5589_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_LC_5_19_5 .C_ON=1'b0;
    defparam \c0.i13_4_lut_LC_5_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_LC_5_19_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i13_4_lut_LC_5_19_5  (
            .in0(N__15636),
            .in1(N__15387),
            .in2(N__15381),
            .in3(N__24621),
            .lcout(\c0.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_955_LC_5_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_955_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_955_LC_5_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_955_LC_5_19_7  (
            .in0(_gnd_net_),
            .in1(N__19388),
            .in2(_gnd_net_),
            .in3(N__15359),
            .lcout(\c0.n1994 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_971_LC_5_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_971_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_971_LC_5_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_971_LC_5_20_0  (
            .in0(N__21699),
            .in1(N__20741),
            .in2(N__26675),
            .in3(N__20555),
            .lcout(\c0.n5557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_807_LC_5_20_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_807_LC_5_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_807_LC_5_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_807_LC_5_20_1  (
            .in0(N__29408),
            .in1(N__16982),
            .in2(N__16602),
            .in3(N__22896),
            .lcout(),
            .ltout(\c0.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_837_LC_5_20_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_837_LC_5_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_837_LC_5_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_837_LC_5_20_2  (
            .in0(N__15653),
            .in1(N__15623),
            .in2(N__15639),
            .in3(N__16950),
            .lcout(\c0.n5574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_845_LC_5_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_845_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_845_LC_5_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_845_LC_5_20_4  (
            .in0(_gnd_net_),
            .in1(N__18789),
            .in2(_gnd_net_),
            .in3(N__18877),
            .lcout(\c0.n5572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_860_LC_5_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_860_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_860_LC_5_20_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_860_LC_5_20_5  (
            .in0(N__21974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20847),
            .lcout(\c0.n2000 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i152_LC_5_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i152_LC_5_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i152_LC_5_20_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i152_LC_5_20_6  (
            .in0(N__19791),
            .in1(N__35348),
            .in2(_gnd_net_),
            .in3(N__23136),
            .lcout(data_in_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37494),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i32_LC_5_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i32_LC_5_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i32_LC_5_21_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i32_LC_5_21_0  (
            .in0(N__18198),
            .in1(N__32239),
            .in2(N__32838),
            .in3(N__30522),
            .lcout(\c0.data_in_field_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37504),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i72_LC_5_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i72_LC_5_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i72_LC_5_21_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i72_LC_5_21_1  (
            .in0(N__32237),
            .in1(N__32639),
            .in2(N__30775),
            .in3(N__15612),
            .lcout(\c0.data_in_field_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37504),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i138_LC_5_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i138_LC_5_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i138_LC_5_21_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i138_LC_5_21_2  (
            .in0(N__32637),
            .in1(N__32238),
            .in2(N__15582),
            .in3(N__30881),
            .lcout(\c0.data_in_field_137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37504),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1006_LC_5_21_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1006_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1006_LC_5_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1006_LC_5_21_4  (
            .in0(N__21178),
            .in1(N__28126),
            .in2(N__27260),
            .in3(N__15758),
            .lcout(),
            .ltout(\c0.n18_adj_1959_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1008_LC_5_21_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1008_LC_5_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1008_LC_5_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1008_LC_5_21_5  (
            .in0(N__22712),
            .in1(N__15736),
            .in2(N__15714),
            .in3(N__19101),
            .lcout(),
            .ltout(\c0.n20_adj_1870_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_5_21_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_5_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_LC_5_21_6  (
            .in0(N__19323),
            .in1(N__15711),
            .in2(N__15702),
            .in3(N__17394),
            .lcout(\c0.n5577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i125_LC_5_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i125_LC_5_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i125_LC_5_21_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i125_LC_5_21_7  (
            .in0(N__32236),
            .in1(N__32638),
            .in2(N__30324),
            .in3(N__21537),
            .lcout(\c0.data_in_field_124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37504),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i42_LC_5_22_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i42_LC_5_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i42_LC_5_22_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i42_LC_5_22_0  (
            .in0(N__16867),
            .in1(N__22452),
            .in2(N__32987),
            .in3(N__32292),
            .lcout(\c0.data_in_field_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i13_LC_5_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i13_LC_5_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i13_LC_5_22_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i13_LC_5_22_1  (
            .in0(N__32290),
            .in1(N__23062),
            .in2(N__21765),
            .in3(N__32773),
            .lcout(\c0.data_in_field_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i103_LC_5_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i103_LC_5_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i103_LC_5_22_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i103_LC_5_22_2  (
            .in0(N__32769),
            .in1(N__32291),
            .in2(N__17793),
            .in3(N__17504),
            .lcout(\c0.data_in_field_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37512),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_LC_5_22_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_5_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_5_22_3  (
            .in0(N__21527),
            .in1(N__17500),
            .in2(N__16868),
            .in3(N__21743),
            .lcout(\c0.n2101 ),
            .ltout(\c0.n2101_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_901_LC_5_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_901_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_901_LC_5_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_901_LC_5_22_4  (
            .in0(N__28306),
            .in1(N__24868),
            .in2(N__15693),
            .in3(N__26801),
            .lcout(),
            .ltout(\c0.n6_adj_1917_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_848_LC_5_22_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_848_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_848_LC_5_22_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_848_LC_5_22_5  (
            .in0(N__17211),
            .in1(N__28020),
            .in2(N__15690),
            .in3(N__15683),
            .lcout(\c0.n5512 ),
            .ltout(\c0.n5512_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_808_LC_5_22_6 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_808_LC_5_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_808_LC_5_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_808_LC_5_22_6  (
            .in0(N__17318),
            .in1(N__19074),
            .in2(N__15885),
            .in3(N__19557),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_929_LC_5_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_929_LC_5_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_929_LC_5_22_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_929_LC_5_22_7  (
            .in0(N__21528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17499),
            .lcout(\c0.n2026 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_924_LC_5_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_924_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_924_LC_5_23_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_924_LC_5_23_0  (
            .in0(_gnd_net_),
            .in1(N__15943),
            .in2(_gnd_net_),
            .in3(N__17124),
            .lcout(\c0.n2155 ),
            .ltout(\c0.n2155_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_LC_5_23_1 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_5_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i16_4_lut_LC_5_23_1  (
            .in0(N__16545),
            .in1(N__19589),
            .in2(N__15861),
            .in3(N__15792),
            .lcout(\c0.n43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i18_LC_5_23_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i18_LC_5_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i18_LC_5_23_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i18_LC_5_23_2  (
            .in0(N__18290),
            .in1(N__32295),
            .in2(N__33068),
            .in3(N__15944),
            .lcout(\c0.data_in_field_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_991_LC_5_23_3 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_991_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_991_LC_5_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_991_LC_5_23_3  (
            .in0(N__22763),
            .in1(N__15833),
            .in2(N__15984),
            .in3(N__29382),
            .lcout(\c0.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i130_LC_5_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i130_LC_5_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i130_LC_5_23_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i130_LC_5_23_4  (
            .in0(N__32839),
            .in1(N__32294),
            .in2(N__15822),
            .in3(N__17125),
            .lcout(\c0.data_in_field_129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i159_LC_5_23_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i159_LC_5_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i159_LC_5_23_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i159_LC_5_23_5  (
            .in0(N__15981),
            .in1(N__35347),
            .in2(_gnd_net_),
            .in3(N__16032),
            .lcout(data_in_19_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_903_LC_5_23_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_903_LC_5_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_903_LC_5_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_903_LC_5_23_6  (
            .in0(N__15791),
            .in1(N__17588),
            .in2(N__17353),
            .in3(N__15773),
            .lcout(\c0.n5491 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i151_LC_5_23_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i151_LC_5_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i151_LC_5_23_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i151_LC_5_23_7  (
            .in0(N__15982),
            .in1(N__35346),
            .in2(_gnd_net_),
            .in3(N__16138),
            .lcout(data_in_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37523),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i113_LC_5_24_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i113_LC_5_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i113_LC_5_24_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i113_LC_5_24_0  (
            .in0(N__32587),
            .in1(N__32286),
            .in2(N__19695),
            .in3(N__17373),
            .lcout(\c0.data_in_field_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i153_LC_5_24_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i153_LC_5_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i153_LC_5_24_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i153_LC_5_24_1  (
            .in0(N__32285),
            .in1(N__32588),
            .in2(N__15963),
            .in3(N__21910),
            .lcout(\c0.data_in_frame_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i158_LC_5_24_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i158_LC_5_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i158_LC_5_24_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i158_LC_5_24_2  (
            .in0(N__35343),
            .in1(N__16047),
            .in2(_gnd_net_),
            .in3(N__19714),
            .lcout(data_in_19_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5739_LC_5_24_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5739_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5739_LC_5_24_3 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5739_LC_5_24_3  (
            .in0(N__27664),
            .in1(N__30016),
            .in2(N__30845),
            .in3(N__15945),
            .lcout(),
            .ltout(\c0.n6093_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6093_bdd_4_lut_LC_5_24_4 .C_ON=1'b0;
    defparam \c0.n6093_bdd_4_lut_LC_5_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.n6093_bdd_4_lut_LC_5_24_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6093_bdd_4_lut_LC_5_24_4  (
            .in0(N__30017),
            .in1(N__30975),
            .in2(N__15930),
            .in3(N__18432),
            .lcout(\c0.n5767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i97_LC_5_24_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i97_LC_5_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i97_LC_5_24_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i97_LC_5_24_5  (
            .in0(N__25756),
            .in1(N__35345),
            .in2(_gnd_net_),
            .in3(N__19670),
            .lcout(data_in_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i131_LC_5_24_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i131_LC_5_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i131_LC_5_24_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i131_LC_5_24_6  (
            .in0(N__35342),
            .in1(N__25691),
            .in2(_gnd_net_),
            .in3(N__15907),
            .lcout(data_in_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i23_LC_5_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i23_LC_5_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i23_LC_5_24_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i23_LC_5_24_7  (
            .in0(N__20249),
            .in1(N__35344),
            .in2(_gnd_net_),
            .in3(N__27795),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37536),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i151_LC_5_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i151_LC_5_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i151_LC_5_25_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i151_LC_5_25_0  (
            .in0(N__16109),
            .in1(N__32296),
            .in2(N__16146),
            .in3(N__32590),
            .lcout(\c0.data_in_frame_18_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i152_LC_5_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i152_LC_5_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i152_LC_5_25_5 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i152_LC_5_25_5  (
            .in0(N__32589),
            .in1(N__16094),
            .in2(N__23156),
            .in3(N__32304),
            .lcout(\c0.data_in_frame_18_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i50_LC_5_25_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i50_LC_5_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i50_LC_5_25_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i50_LC_5_25_7  (
            .in0(N__36047),
            .in1(N__16079),
            .in2(_gnd_net_),
            .in3(N__22463),
            .lcout(data_in_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37546),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_791_LC_5_26_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_791_LC_5_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_791_LC_5_26_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.rx.i1_2_lut_adj_791_LC_5_26_0  (
            .in0(_gnd_net_),
            .in1(N__20404),
            .in2(_gnd_net_),
            .in3(N__19951),
            .lcout(n1764),
            .ltout(n1764_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_5_26_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_5_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_5_26_1 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_5_26_1  (
            .in0(N__20344),
            .in1(N__16043),
            .in2(N__16050),
            .in3(N__15990),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37556),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5854_LC_5_26_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5854_LC_5_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5854_LC_5_26_2 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5854_LC_5_26_2  (
            .in0(N__27613),
            .in1(N__18790),
            .in2(N__30093),
            .in3(N__18828),
            .lcout(\c0.n6237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_5_26_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_5_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_5_26_3 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_5_26_3  (
            .in0(N__20093),
            .in1(N__18057),
            .in2(N__20361),
            .in3(N__16028),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37556),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i2_LC_5_26_4 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i2_LC_5_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_5_26_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_5_26_4  (
            .in0(N__16224),
            .in1(N__16010),
            .in2(_gnd_net_),
            .in3(N__16017),
            .lcout(\c0.rx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37556),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_26_i4_2_lut_LC_5_26_5 .C_ON=1'b0;
    defparam \c0.rx.equal_26_i4_2_lut_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_26_i4_2_lut_LC_5_26_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.rx.equal_26_i4_2_lut_LC_5_26_5  (
            .in0(N__20044),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20004),
            .lcout(n4_adj_1980),
            .ltout(n4_adj_1980_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_5_26_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_5_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_5_26_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_5_26_6  (
            .in0(N__16236),
            .in1(N__20345),
            .in2(N__16239),
            .in3(N__20092),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37556),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i157_LC_5_26_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i157_LC_5_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i157_LC_5_26_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i157_LC_5_26_7  (
            .in0(N__35349),
            .in1(N__16235),
            .in2(_gnd_net_),
            .in3(N__20646),
            .lcout(data_in_19_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37556),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i5287_3_lut_4_lut_LC_5_27_1 .C_ON=1'b0;
    defparam \c0.rx.i5287_3_lut_4_lut_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i5287_3_lut_4_lut_LC_5_27_1 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \c0.rx.i5287_3_lut_4_lut_LC_5_27_1  (
            .in0(N__17638),
            .in1(N__16307),
            .in2(N__18017),
            .in3(N__17690),
            .lcout(\c0.rx.n5633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_3_lut_4_lut_4_lut_LC_5_27_3.C_ON=1'b0;
    defparam i13_3_lut_4_lut_4_lut_LC_5_27_3.SEQ_MODE=4'b0000;
    defparam i13_3_lut_4_lut_4_lut_LC_5_27_3.LUT_INIT=16'b0010000000001111;
    LogicCell40 i13_3_lut_4_lut_4_lut_LC_5_27_3 (
            .in0(N__17637),
            .in1(N__16306),
            .in2(N__18018),
            .in3(N__17689),
            .lcout(),
            .ltout(n2198_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_5_27_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_5_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_5_27_4 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_5_27_4  (
            .in0(N__16308),
            .in1(N__35261),
            .in2(N__16227),
            .in3(N__18003),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37566),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i7_LC_5_27_5 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_5_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_5_27_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_5_27_5  (
            .in0(N__16223),
            .in1(N__16173),
            .in2(_gnd_net_),
            .in3(N__16179),
            .lcout(\c0.rx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37566),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i87_LC_5_27_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i87_LC_5_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i87_LC_5_27_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i87_LC_5_27_6  (
            .in0(N__35255),
            .in1(N__19043),
            .in2(_gnd_net_),
            .in3(N__17461),
            .lcout(data_in_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37566),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_3_lut_4_lut_LC_5_28_0 .C_ON=1'b0;
    defparam \c0.rx.i1_3_lut_4_lut_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_3_lut_4_lut_LC_5_28_0 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.rx.i1_3_lut_4_lut_LC_5_28_0  (
            .in0(N__16295),
            .in1(N__17684),
            .in2(N__18006),
            .in3(N__17635),
            .lcout(\c0.rx.n2259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.n6291_bdd_4_lut_LC_5_28_1 .C_ON=1'b0;
    defparam \c0.rx.n6291_bdd_4_lut_LC_5_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.n6291_bdd_4_lut_LC_5_28_1 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.rx.n6291_bdd_4_lut_LC_5_28_1  (
            .in0(N__16155),
            .in1(N__17983),
            .in2(N__20359),
            .in3(N__17598),
            .lcout(),
            .ltout(\c0.rx.n6294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_5_28_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_5_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_5_28_2 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_5_28_2  (
            .in0(N__16296),
            .in1(_gnd_net_),
            .in2(N__16311),
            .in3(_gnd_net_),
            .lcout(r_SM_Main_0_adj_1991),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_LC_5_28_4 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_LC_5_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_LC_5_28_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.rx.i2_4_lut_LC_5_28_4  (
            .in0(N__16294),
            .in1(N__17683),
            .in2(N__18005),
            .in3(N__17634),
            .lcout(\c0.rx.n1706 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i90_2_lut_LC_5_28_5 .C_ON=1'b0;
    defparam \c0.rx.i90_2_lut_LC_5_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i90_2_lut_LC_5_28_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \c0.rx.i90_2_lut_LC_5_28_5  (
            .in0(N__17636),
            .in1(_gnd_net_),
            .in2(N__17696),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.rx.n75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_5_28_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_5_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_5_28_6 .LUT_INIT=16'b0001010100000100;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_5_28_6  (
            .in0(N__16297),
            .in1(N__18004),
            .in2(N__16251),
            .in3(N__16248),
            .lcout(r_SM_Main_1_adj_1990),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_5_28_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_5_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_5_28_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_5_28_7  (
            .in0(N__33570),
            .in1(N__23862),
            .in2(_gnd_net_),
            .in3(N__21638),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37574),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_5_29_2 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_5_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_5_29_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_5_29_2  (
            .in0(N__20043),
            .in1(N__20417),
            .in2(_gnd_net_),
            .in3(N__19999),
            .lcout(\c0.rx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37581),
            .ce(N__17927),
            .sr(N__17898));
    defparam \c0.data_in_0___i67_LC_6_15_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i67_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i67_LC_6_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i67_LC_6_15_0  (
            .in0(N__35634),
            .in1(N__23897),
            .in2(_gnd_net_),
            .in3(N__16729),
            .lcout(data_in_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i36_LC_6_15_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i36_LC_6_15_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i36_LC_6_15_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i36_LC_6_15_2  (
            .in0(N__35633),
            .in1(N__22108),
            .in2(_gnd_net_),
            .in3(N__16713),
            .lcout(data_in_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_886_LC_6_15_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_886_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_886_LC_6_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i9_4_lut_adj_886_LC_6_15_3  (
            .in0(N__16488),
            .in1(N__18235),
            .in2(N__23069),
            .in3(N__22055),
            .lcout(\c0.n25_adj_1929 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i12_LC_6_15_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i12_LC_6_15_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i12_LC_6_15_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i12_LC_6_15_6  (
            .in0(N__35632),
            .in1(N__21101),
            .in2(_gnd_net_),
            .in3(N__16489),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i4_LC_6_15_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i4_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i4_LC_6_15_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i4_LC_6_15_7  (
            .in0(N__16490),
            .in1(N__35635),
            .in2(_gnd_net_),
            .in3(N__18329),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37495),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i52_LC_6_16_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i52_LC_6_16_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i52_LC_6_16_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i52_LC_6_16_0  (
            .in0(N__33268),
            .in1(N__31715),
            .in2(N__16473),
            .in3(N__18726),
            .lcout(\c0.data_in_field_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37488),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i92_LC_6_16_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i92_LC_6_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i92_LC_6_16_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i92_LC_6_16_2  (
            .in0(N__35827),
            .in1(N__16933),
            .in2(_gnd_net_),
            .in3(N__16445),
            .lcout(data_in_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37488),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i2_LC_6_16_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i2_LC_6_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i2_LC_6_16_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i2_LC_6_16_3  (
            .in0(N__16565),
            .in1(N__16330),
            .in2(_gnd_net_),
            .in3(N__35829),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37488),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i100_LC_6_16_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i100_LC_6_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i100_LC_6_16_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i100_LC_6_16_4  (
            .in0(N__33267),
            .in1(N__31714),
            .in2(N__17209),
            .in3(N__16446),
            .lcout(\c0.data_in_field_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37488),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i5_LC_6_16_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i5_LC_6_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i5_LC_6_16_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i5_LC_6_16_5  (
            .in0(N__18509),
            .in1(N__23070),
            .in2(_gnd_net_),
            .in3(N__35828),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37488),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i14_LC_6_16_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i14_LC_6_16_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i14_LC_6_16_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i14_LC_6_16_6  (
            .in0(N__35826),
            .in1(N__17869),
            .in2(_gnd_net_),
            .in3(N__25045),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37488),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_885_LC_6_16_7 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_885_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_885_LC_6_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i11_4_lut_adj_885_LC_6_16_7  (
            .in0(N__18508),
            .in1(N__16329),
            .in2(N__16431),
            .in3(N__16561),
            .lcout(\c0.n27_adj_1928 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_985_LC_6_17_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_985_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_985_LC_6_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_985_LC_6_17_0  (
            .in0(N__20164),
            .in1(N__19639),
            .in2(N__19790),
            .in3(N__16362),
            .lcout(\c0.n22_adj_1886 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i10_LC_6_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i10_LC_6_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i10_LC_6_17_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i10_LC_6_17_1  (
            .in0(N__31705),
            .in1(N__16331),
            .in2(N__18423),
            .in3(N__33163),
            .lcout(\c0.data_in_field_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37478),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i8_LC_6_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i8_LC_6_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i8_LC_6_17_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i8_LC_6_17_2  (
            .in0(N__18105),
            .in1(N__31709),
            .in2(N__33242),
            .in3(N__16594),
            .lcout(\c0.data_in_field_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37478),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i2_LC_6_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i2_LC_6_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i2_LC_6_17_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i2_LC_6_17_3  (
            .in0(N__31706),
            .in1(N__33159),
            .in2(N__16566),
            .in3(N__30966),
            .lcout(\c0.data_in_field_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37478),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i6_LC_6_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i6_LC_6_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i6_LC_6_17_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i6_LC_6_17_5  (
            .in0(N__31707),
            .in1(N__20211),
            .in2(N__22823),
            .in3(N__33164),
            .lcout(\c0.data_in_field_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37478),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i108_LC_6_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i108_LC_6_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i108_LC_6_17_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i108_LC_6_17_6  (
            .in0(N__33158),
            .in1(N__31708),
            .in2(N__26337),
            .in3(N__22959),
            .lcout(\c0.data_in_field_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37478),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i32_LC_6_17_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i32_LC_6_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i32_LC_6_17_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i32_LC_6_17_7  (
            .in0(N__18186),
            .in1(N__35830),
            .in2(_gnd_net_),
            .in3(N__31443),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37478),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i22_LC_6_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i22_LC_6_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i22_LC_6_18_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i22_LC_6_18_0  (
            .in0(N__31710),
            .in1(N__33086),
            .in2(N__17877),
            .in3(N__27131),
            .lcout(\c0.data_in_field_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37489),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_967_LC_6_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_967_LC_6_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_967_LC_6_18_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_967_LC_6_18_1  (
            .in0(N__22813),
            .in1(_gnd_net_),
            .in2(N__21798),
            .in3(N__17154),
            .lcout(\c0.n2104 ),
            .ltout(\c0.n2104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_871_LC_6_18_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_871_LC_6_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_871_LC_6_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_871_LC_6_18_2  (
            .in0(N__16533),
            .in1(N__16611),
            .in2(N__16527),
            .in3(N__20688),
            .lcout(\c0.n5497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i66_LC_6_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i66_LC_6_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i66_LC_6_18_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i66_LC_6_18_3  (
            .in0(N__33085),
            .in1(N__31712),
            .in2(N__16524),
            .in3(N__17155),
            .lcout(\c0.data_in_field_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37489),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i81_LC_6_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i81_LC_6_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i81_LC_6_18_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i81_LC_6_18_4  (
            .in0(N__31711),
            .in1(N__33087),
            .in2(N__21982),
            .in3(N__30452),
            .lcout(\c0.data_in_field_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37489),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_966_LC_6_18_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_966_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_966_LC_6_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_966_LC_6_18_5  (
            .in0(N__22812),
            .in1(N__17153),
            .in2(N__27137),
            .in3(N__16617),
            .lcout(\c0.n5521 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_896_LC_6_18_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_896_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_896_LC_6_18_6 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_896_LC_6_18_6  (
            .in0(N__17311),
            .in1(N__18464),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n5476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_1002_LC_6_18_7 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_1002_LC_6_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_1002_LC_6_18_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_1002_LC_6_18_7  (
            .in0(N__18585),
            .in1(N__20740),
            .in2(N__26645),
            .in3(N__22544),
            .lcout(\c0.n20_adj_1958 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_6_19_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_6_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_6_19_0  (
            .in0(N__16767),
            .in1(N__26611),
            .in2(N__21227),
            .in3(N__24437),
            .lcout(),
            .ltout(\c0.n31_adj_1896_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_adj_829_LC_6_19_1 .C_ON=1'b0;
    defparam \c0.i21_4_lut_adj_829_LC_6_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_adj_829_LC_6_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_adj_829_LC_6_19_1  (
            .in0(N__21693),
            .in1(N__22350),
            .in2(N__16659),
            .in3(N__16656),
            .lcout(\c0.n47_adj_1897 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_843_LC_6_19_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_843_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_843_LC_6_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_843_LC_6_19_2  (
            .in0(N__16646),
            .in1(N__20516),
            .in2(N__19021),
            .in3(N__24707),
            .lcout(\c0.n10_adj_1915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i110_LC_6_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i110_LC_6_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i110_LC_6_19_3 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i110_LC_6_19_3  (
            .in0(N__26612),
            .in1(N__32763),
            .in2(N__34491),
            .in3(N__31887),
            .lcout(\c0.data_in_field_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i126_LC_6_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i126_LC_6_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i126_LC_6_19_4 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i126_LC_6_19_4  (
            .in0(N__31882),
            .in1(N__21309),
            .in2(N__32986),
            .in3(N__17310),
            .lcout(\c0.data_in_field_125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_944_LC_6_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_944_LC_6_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_944_LC_6_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_944_LC_6_19_5  (
            .in0(N__17309),
            .in1(N__18470),
            .in2(_gnd_net_),
            .in3(N__16766),
            .lcout(\c0.n1913 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i65_LC_6_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i65_LC_6_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i65_LC_6_19_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0___i65_LC_6_19_6  (
            .in0(N__32762),
            .in1(N__16788),
            .in2(N__32100),
            .in3(N__31062),
            .lcout(\c0.data_in_field_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i136_LC_6_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i136_LC_6_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i136_LC_6_19_7 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i136_LC_6_19_7  (
            .in0(N__22425),
            .in1(N__31883),
            .in2(N__17283),
            .in3(N__32767),
            .lcout(\c0.data_in_field_135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37496),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i11_LC_6_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i11_LC_6_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i11_LC_6_20_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i11_LC_6_20_0  (
            .in0(N__22020),
            .in1(N__32054),
            .in2(N__33276),
            .in3(N__16897),
            .lcout(\c0.data_in_field_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i67_LC_6_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i67_LC_6_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i67_LC_6_20_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i67_LC_6_20_1  (
            .in0(N__32053),
            .in1(N__33263),
            .in2(N__16743),
            .in3(N__20950),
            .lcout(\c0.data_in_field_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i141_LC_6_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i141_LC_6_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i141_LC_6_20_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i141_LC_6_20_2  (
            .in0(N__33261),
            .in1(N__32055),
            .in2(N__27395),
            .in3(N__18881),
            .lcout(\c0.data_in_field_140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i44_LC_6_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i44_LC_6_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i44_LC_6_20_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i44_LC_6_20_3  (
            .in0(N__32052),
            .in1(N__33262),
            .in2(N__16712),
            .in3(N__19106),
            .lcout(\c0.data_in_field_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37505),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5839_LC_6_20_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5839_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5839_LC_6_20_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5839_LC_6_20_4  (
            .in0(N__27686),
            .in1(N__19338),
            .in2(N__30149),
            .in3(N__27133),
            .lcout(\c0.n6219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5809_LC_6_20_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5809_LC_6_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5809_LC_6_20_5 .LUT_INIT=16'b1011100011001100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5809_LC_6_20_5  (
            .in0(N__22650),
            .in1(N__27687),
            .in2(N__19164),
            .in3(N__30065),
            .lcout(\c0.n6183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_936_LC_6_20_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_936_LC_6_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_936_LC_6_20_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_936_LC_6_20_6  (
            .in0(_gnd_net_),
            .in1(N__30607),
            .in2(_gnd_net_),
            .in3(N__27132),
            .lcout(),
            .ltout(\c0.n2062_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_LC_6_20_7 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_6_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_LC_6_20_7  (
            .in0(N__19260),
            .in1(N__18823),
            .in2(N__17046),
            .in3(N__18624),
            .lcout(\c0.n44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_6_21_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_6_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_LC_6_21_0  (
            .in0(N__24746),
            .in1(N__17027),
            .in2(N__18958),
            .in3(N__16836),
            .lcout(\c0.n5503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_6_21_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_6_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_6_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_LC_6_21_1  (
            .in0(N__16911),
            .in1(N__16971),
            .in2(N__24180),
            .in3(N__17237),
            .lcout(\c0.n16_adj_1871 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i92_LC_6_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i92_LC_6_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i92_LC_6_21_3 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i92_LC_6_21_3  (
            .in0(N__32089),
            .in1(N__16943),
            .in2(N__33275),
            .in3(N__27951),
            .lcout(\c0.data_in_field_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37513),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_863_LC_6_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_863_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_863_LC_6_21_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_863_LC_6_21_4  (
            .in0(_gnd_net_),
            .in1(N__20943),
            .in2(_gnd_net_),
            .in3(N__19159),
            .lcout(\c0.n2021 ),
            .ltout(\c0.n2021_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_864_LC_6_21_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_864_LC_6_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_864_LC_6_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_864_LC_6_21_5  (
            .in0(N__16890),
            .in1(N__16812),
            .in2(N__16872),
            .in3(N__26800),
            .lcout(\c0.n2074 ),
            .ltout(\c0.n2074_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_976_LC_6_21_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_976_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_976_LC_6_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_976_LC_6_21_6  (
            .in0(N__16860),
            .in1(N__22742),
            .in2(N__16839),
            .in3(N__16835),
            .lcout(\c0.n5527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i27_LC_6_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i27_LC_6_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i27_LC_6_21_7 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i27_LC_6_21_7  (
            .in0(N__32088),
            .in1(N__21486),
            .in2(N__33274),
            .in3(N__16813),
            .lcout(\c0.data_in_field_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37513),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i134_LC_6_22_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i134_LC_6_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i134_LC_6_22_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i134_LC_6_22_0  (
            .in0(N__18694),
            .in1(N__21347),
            .in2(_gnd_net_),
            .in3(N__35965),
            .lcout(data_in_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_LC_6_22_1 .C_ON=1'b0;
    defparam \c0.i22_4_lut_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_LC_6_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i22_4_lut_LC_6_22_1  (
            .in0(N__19070),
            .in1(N__27210),
            .in2(N__17409),
            .in3(N__17379),
            .lcout(\c0.n48_adj_1895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_923_LC_6_22_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_923_LC_6_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_923_LC_6_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_923_LC_6_22_2  (
            .in0(N__27940),
            .in1(N__19207),
            .in2(N__19469),
            .in3(N__17273),
            .lcout(\c0.n5418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i75_LC_6_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i75_LC_6_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i75_LC_6_22_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i75_LC_6_22_3  (
            .in0(N__32293),
            .in1(N__32768),
            .in2(N__23910),
            .in3(N__31000),
            .lcout(\c0.data_in_field_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_898_LC_6_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_898_LC_6_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_898_LC_6_22_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_898_LC_6_22_5  (
            .in0(_gnd_net_),
            .in1(N__27941),
            .in2(_gnd_net_),
            .in3(N__19461),
            .lcout(\c0.n1908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_919_LC_6_22_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_919_LC_6_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_919_LC_6_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_919_LC_6_22_6  (
            .in0(N__17441),
            .in1(N__17210),
            .in2(N__30768),
            .in3(N__24581),
            .lcout(\c0.n1889 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i126_LC_6_22_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i126_LC_6_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i126_LC_6_22_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i126_LC_6_22_7  (
            .in0(N__35964),
            .in1(N__18695),
            .in2(_gnd_net_),
            .in3(N__21289),
            .lcout(data_in_15_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37524),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i127_LC_6_23_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i127_LC_6_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i127_LC_6_23_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i127_LC_6_23_0  (
            .in0(N__18813),
            .in1(N__17730),
            .in2(N__32222),
            .in3(N__32602),
            .lcout(\c0.data_in_field_126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_910_LC_6_23_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_910_LC_6_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_910_LC_6_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_910_LC_6_23_1  (
            .in0(N__25947),
            .in1(N__17162),
            .in2(_gnd_net_),
            .in3(N__17126),
            .lcout(\c0.n5569 ),
            .ltout(\c0.n5569_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_LC_6_23_2 .C_ON=1'b0;
    defparam \c0.i7_3_lut_LC_6_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_LC_6_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i7_3_lut_LC_6_23_2  (
            .in0(_gnd_net_),
            .in1(N__25727),
            .in2(N__17094),
            .in3(N__17091),
            .lcout(\c0.n20_adj_1882 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_908_LC_6_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_908_LC_6_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_908_LC_6_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_908_LC_6_23_3  (
            .in0(N__19232),
            .in1(N__30993),
            .in2(N__23013),
            .in3(N__17565),
            .lcout(\c0.n1958 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_938_LC_6_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_938_LC_6_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_938_LC_6_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_938_LC_6_23_4  (
            .in0(N__17566),
            .in1(N__23003),
            .in2(_gnd_net_),
            .in3(N__19233),
            .lcout(\c0.n5388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i79_LC_6_23_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i79_LC_6_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i79_LC_6_23_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i79_LC_6_23_5  (
            .in0(N__19234),
            .in1(N__31193),
            .in2(N__32780),
            .in3(N__32099),
            .lcout(\c0.data_in_field_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37537),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_adj_988_LC_6_23_6 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_988_LC_6_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_988_LC_6_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i18_4_lut_adj_988_LC_6_23_6  (
            .in0(N__17400),
            .in1(N__19245),
            .in2(N__22895),
            .in3(N__17390),
            .lcout(\c0.n44_adj_1894 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_881_LC_6_23_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_881_LC_6_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_881_LC_6_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_881_LC_6_23_7  (
            .in0(N__17371),
            .in1(N__18812),
            .in2(_gnd_net_),
            .in3(N__17564),
            .lcout(\c0.n5524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_926_LC_6_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_926_LC_6_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_926_LC_6_24_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_926_LC_6_24_0  (
            .in0(_gnd_net_),
            .in1(N__17346),
            .in2(_gnd_net_),
            .in3(N__17435),
            .lcout(\c0.n1917 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i160_LC_6_24_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i160_LC_6_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i160_LC_6_24_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i160_LC_6_24_1  (
            .in0(N__19789),
            .in1(N__17748),
            .in2(_gnd_net_),
            .in3(N__36046),
            .lcout(data_in_19_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37547),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i31_LC_6_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i31_LC_6_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i31_LC_6_24_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i31_LC_6_24_2  (
            .in0(N__32847),
            .in1(N__32288),
            .in2(N__17355),
            .in3(N__20250),
            .lcout(\c0.data_in_field_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37547),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5824_LC_6_24_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5824_LC_6_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5824_LC_6_24_3 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5824_LC_6_24_3  (
            .in0(N__27663),
            .in1(N__22206),
            .in2(N__30112),
            .in3(N__17322),
            .lcout(\c0.n6201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_986_LC_6_24_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_986_LC_6_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_986_LC_6_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_986_LC_6_24_4  (
            .in0(N__22674),
            .in1(N__19553),
            .in2(N__30264),
            .in3(N__17592),
            .lcout(\c0.n18_adj_1887 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i77_LC_6_24_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i77_LC_6_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i77_LC_6_24_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i77_LC_6_24_5  (
            .in0(N__32287),
            .in1(N__30390),
            .in2(N__17576),
            .in3(N__32846),
            .lcout(\c0.data_in_field_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37547),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i149_LC_6_24_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i149_LC_6_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i149_LC_6_24_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i149_LC_6_24_6  (
            .in0(N__17543),
            .in1(N__20123),
            .in2(N__33069),
            .in3(N__32289),
            .lcout(\c0.data_in_frame_18_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37547),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i141_LC_6_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i141_LC_6_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i141_LC_6_24_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i141_LC_6_24_7  (
            .in0(N__20122),
            .in1(N__36045),
            .in2(_gnd_net_),
            .in3(N__27379),
            .lcout(data_in_17_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37547),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5859_LC_6_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5859_LC_6_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5859_LC_6_25_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5859_LC_6_25_0  (
            .in0(N__27685),
            .in1(N__21003),
            .in2(N__30184),
            .in3(N__17439),
            .lcout(),
            .ltout(\c0.n6243_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6243_bdd_4_lut_LC_6_25_1 .C_ON=1'b0;
    defparam \c0.n6243_bdd_4_lut_LC_6_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.n6243_bdd_4_lut_LC_6_25_1 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n6243_bdd_4_lut_LC_6_25_1  (
            .in0(N__29513),
            .in1(N__19239),
            .in2(N__17529),
            .in3(N__30125),
            .lcout(),
            .ltout(\c0.n5698_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5869_LC_6_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5869_LC_6_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5869_LC_6_25_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5869_LC_6_25_2  (
            .in0(N__25402),
            .in1(N__25252),
            .in2(N__17526),
            .in3(N__17481),
            .lcout(\c0.n6231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6237_bdd_4_lut_LC_6_25_3 .C_ON=1'b0;
    defparam \c0.n6237_bdd_4_lut_LC_6_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6237_bdd_4_lut_LC_6_25_3 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n6237_bdd_4_lut_LC_6_25_3  (
            .in0(N__17514),
            .in1(N__23691),
            .in2(N__17508),
            .in3(N__30121),
            .lcout(\c0.n5701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i87_LC_6_25_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i87_LC_6_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i87_LC_6_25_5 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i87_LC_6_25_5  (
            .in0(N__17440),
            .in1(N__17475),
            .in2(N__32303),
            .in3(N__32591),
            .lcout(\c0.data_in_field_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i82_LC_6_25_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i82_LC_6_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i82_LC_6_25_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i82_LC_6_25_6  (
            .in0(N__21248),
            .in1(_gnd_net_),
            .in2(N__35684),
            .in3(N__17837),
            .lcout(data_in_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i74_LC_6_25_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i74_LC_6_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i74_LC_6_25_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i74_LC_6_25_7  (
            .in0(N__17836),
            .in1(N__35511),
            .in2(_gnd_net_),
            .in3(N__17804),
            .lcout(data_in_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37557),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i95_LC_6_26_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i95_LC_6_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i95_LC_6_26_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i95_LC_6_26_0  (
            .in0(N__35260),
            .in1(N__19042),
            .in2(_gnd_net_),
            .in3(N__17783),
            .lcout(data_in_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i103_LC_6_26_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i103_LC_6_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i103_LC_6_26_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i103_LC_6_26_4  (
            .in0(N__35259),
            .in1(N__22915),
            .in2(_gnd_net_),
            .in3(N__17782),
            .lcout(data_in_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_6_26_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_6_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_6_26_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_6_26_6  (
            .in0(N__18056),
            .in1(N__20349),
            .in2(N__17747),
            .in3(N__17759),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37567),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_27_i4_2_lut_LC_6_26_7 .C_ON=1'b0;
    defparam \c0.rx.equal_27_i4_2_lut_LC_6_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_27_i4_2_lut_LC_6_26_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.equal_27_i4_2_lut_LC_6_26_7  (
            .in0(_gnd_net_),
            .in1(N__20045),
            .in2(_gnd_net_),
            .in3(N__20000),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i119_LC_6_27_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i119_LC_6_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i119_LC_6_27_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i119_LC_6_27_2  (
            .in0(N__35257),
            .in1(N__19807),
            .in2(_gnd_net_),
            .in3(N__17726),
            .lcout(data_in_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i98_LC_6_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i98_LC_6_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i98_LC_6_27_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i98_LC_6_27_3  (
            .in0(N__19406),
            .in1(N__35258),
            .in2(_gnd_net_),
            .in3(N__19897),
            .lcout(data_in_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i106_LC_6_27_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i106_LC_6_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i106_LC_6_27_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i106_LC_6_27_4  (
            .in0(N__35256),
            .in1(N__19499),
            .in2(_gnd_net_),
            .in3(N__19405),
            .lcout(data_in_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_6_27_5 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_6_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_6_27_5 .LUT_INIT=16'b1101110000111100;
    LogicCell40 \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_6_27_5  (
            .in0(N__18035),
            .in1(N__17688),
            .in2(N__18016),
            .in3(N__17646),
            .lcout(\c0.rx.n6291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_6_27_6 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_6_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_6_27_6 .LUT_INIT=16'b1000100110001000;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_6_27_6  (
            .in0(N__20411),
            .in1(N__18063),
            .in2(N__18039),
            .in3(N__17996),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i90_LC_6_27_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i90_LC_6_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i90_LC_6_27_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i90_LC_6_27_7  (
            .in0(N__35448),
            .in1(N__21241),
            .in2(_gnd_net_),
            .in3(N__19898),
            .lcout(data_in_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37575),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3393_2_lut_LC_6_28_0 .C_ON=1'b0;
    defparam \c0.rx.i3393_2_lut_LC_6_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3393_2_lut_LC_6_28_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i3393_2_lut_LC_6_28_0  (
            .in0(N__19990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20033),
            .lcout(n3636),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_3_lut_LC_6_28_5 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_3_lut_LC_6_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_3_lut_LC_6_28_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i2_2_lut_3_lut_LC_6_28_5  (
            .in0(N__20032),
            .in1(N__20402),
            .in2(_gnd_net_),
            .in3(N__19989),
            .lcout(\c0.rx.n3850 ),
            .ltout(\c0.rx.n3850_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2116_2_lut_3_lut_LC_6_28_6 .C_ON=1'b0;
    defparam \c0.rx.i2116_2_lut_3_lut_LC_6_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2116_2_lut_3_lut_LC_6_28_6 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \c0.rx.i2116_2_lut_3_lut_LC_6_28_6  (
            .in0(_gnd_net_),
            .in1(N__17992),
            .in2(N__17931),
            .in3(N__17914),
            .lcout(\c0.rx.n2367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_6_29_1 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_6_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_6_29_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_6_29_1  (
            .in0(_gnd_net_),
            .in1(N__20416),
            .in2(_gnd_net_),
            .in3(N__19998),
            .lcout(\c0.rx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37590),
            .ce(N__17928),
            .sr(N__17897));
    defparam \c0.i10_4_lut_adj_882_LC_7_15_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_882_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_882_LC_7_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i10_4_lut_adj_882_LC_7_15_1  (
            .in0(N__18328),
            .in1(N__21099),
            .in2(N__17870),
            .in3(N__28432),
            .lcout(\c0.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i20_LC_7_15_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i20_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i20_LC_7_15_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i20_LC_7_15_4  (
            .in0(N__21100),
            .in1(N__35636),
            .in2(_gnd_net_),
            .in3(N__22087),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37506),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i22_LC_7_15_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i22_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i22_LC_7_15_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \c0.data_in_0___i22_LC_7_15_5  (
            .in0(N__17865),
            .in1(N__27896),
            .in2(N__35825),
            .in3(_gnd_net_),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37506),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_877_LC_7_16_0 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_877_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_877_LC_7_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i12_4_lut_adj_877_LC_7_16_0  (
            .in0(N__18211),
            .in1(N__25044),
            .in2(N__18104),
            .in3(N__18134),
            .lcout(),
            .ltout(\c0.n28_adj_1926_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_956_LC_7_16_1 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_956_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_956_LC_7_16_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i15_4_lut_adj_956_LC_7_16_1  (
            .in0(N__18312),
            .in1(N__18306),
            .in2(N__18300),
            .in3(N__18297),
            .lcout(\c0.n4795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i15_LC_7_16_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i15_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i15_LC_7_16_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i15_LC_7_16_2  (
            .in0(N__35928),
            .in1(N__18152),
            .in2(_gnd_net_),
            .in3(N__27819),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_925_LC_7_16_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_925_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_925_LC_7_16_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_925_LC_7_16_3  (
            .in0(N__20236),
            .in1(N__20184),
            .in2(N__18291),
            .in3(N__27771),
            .lcout(\c0.n30_adj_1941 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i1_LC_7_16_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i1_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i1_LC_7_16_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i1_LC_7_16_4  (
            .in0(N__35931),
            .in1(N__22264),
            .in2(_gnd_net_),
            .in3(N__18248),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i7_LC_7_16_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i7_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i7_LC_7_16_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i7_LC_7_16_5  (
            .in0(N__18151),
            .in1(N__35929),
            .in2(_gnd_net_),
            .in3(N__18212),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_912_LC_7_16_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_912_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_912_LC_7_16_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_912_LC_7_16_6  (
            .in0(N__18193),
            .in1(N__18150),
            .in2(N__24680),
            .in3(N__22309),
            .lcout(\c0.n26_adj_1940 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i8_LC_7_16_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i8_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i8_LC_7_16_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i8_LC_7_16_7  (
            .in0(N__18135),
            .in1(N__35930),
            .in2(_gnd_net_),
            .in3(N__18100),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37497),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_958_LC_7_17_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_958_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_958_LC_7_17_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i1_4_lut_adj_958_LC_7_17_0  (
            .in0(N__18084),
            .in1(N__18078),
            .in2(N__18072),
            .in3(N__21015),
            .lcout(\c0.n1729 ),
            .ltout(\c0.n1729_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i36_LC_7_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i36_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i36_LC_7_17_1 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i36_LC_7_17_1  (
            .in0(N__22116),
            .in1(N__33165),
            .in2(N__18474),
            .in3(N__18465),
            .lcout(\c0.data_in_field_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37484),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i28_LC_7_17_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i28_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i28_LC_7_17_2 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i28_LC_7_17_2  (
            .in0(N__22092),
            .in1(N__31700),
            .in2(N__33243),
            .in3(N__18605),
            .lcout(\c0.data_in_field_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37484),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i55_LC_7_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i55_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i55_LC_7_17_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i55_LC_7_17_3  (
            .in0(N__18358),
            .in1(N__24209),
            .in2(N__31944),
            .in3(N__33173),
            .lcout(\c0.data_in_field_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37484),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_934_LC_7_17_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_934_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_934_LC_7_17_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_934_LC_7_17_4  (
            .in0(N__18402),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18718),
            .lcout(),
            .ltout(\c0.n5369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_935_LC_7_17_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_935_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_935_LC_7_17_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_935_LC_7_17_5  (
            .in0(N__18357),
            .in1(N__18914),
            .in2(N__18339),
            .in3(N__26828),
            .lcout(\c0.n2125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i33_LC_7_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i33_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i33_LC_7_17_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i33_LC_7_17_6  (
            .in0(N__26829),
            .in1(N__23496),
            .in2(N__33244),
            .in3(N__31704),
            .lcout(\c0.data_in_field_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37484),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i4_LC_7_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i4_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i4_LC_7_17_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i4_LC_7_17_7  (
            .in0(N__31699),
            .in1(N__33166),
            .in2(N__18336),
            .in3(N__18646),
            .lcout(\c0.data_in_field_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37484),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i56_LC_7_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i56_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i56_LC_7_18_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i56_LC_7_18_0  (
            .in0(N__21070),
            .in1(N__35927),
            .in2(_gnd_net_),
            .in3(N__23267),
            .lcout(data_in_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37498),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i3_LC_7_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i3_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i3_LC_7_18_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i3_LC_7_18_1  (
            .in0(N__35926),
            .in1(N__24670),
            .in2(_gnd_net_),
            .in3(N__22019),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37498),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i76_LC_7_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i76_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i76_LC_7_18_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i76_LC_7_18_2  (
            .in0(N__33084),
            .in1(N__31713),
            .in2(N__18681),
            .in3(N__19020),
            .lcout(\c0.data_in_field_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37498),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_869_LC_7_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_869_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_869_LC_7_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_869_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(N__18640),
            .in2(_gnd_net_),
            .in3(N__18620),
            .lcout(\c0.n6_adj_1923 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_867_LC_7_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_867_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_867_LC_7_18_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_867_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(N__18601),
            .in2(_gnd_net_),
            .in3(N__20471),
            .lcout(\c0.n5469 ),
            .ltout(\c0.n5469_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_870_LC_7_18_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_870_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_870_LC_7_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_870_LC_7_18_5  (
            .in0(N__18573),
            .in1(N__18540),
            .in2(N__18525),
            .in3(N__18522),
            .lcout(\c0.n5548 ),
            .ltout(\c0.n5548_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_7_18_6 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_7_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_LC_7_18_6  (
            .in0(N__22691),
            .in1(N__20495),
            .in2(N__18516),
            .in3(N__24401),
            .lcout(\c0.n45_adj_1892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i5_LC_7_19_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i5_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i5_LC_7_19_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i5_LC_7_19_0  (
            .in0(N__18513),
            .in1(N__32059),
            .in2(N__33233),
            .in3(N__21797),
            .lcout(\c0.data_in_field_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37507),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i62_LC_7_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i62_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i62_LC_7_19_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i62_LC_7_19_1  (
            .in0(N__32056),
            .in1(N__33131),
            .in2(N__18495),
            .in3(N__22346),
            .lcout(\c0.data_in_field_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37507),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i116_LC_7_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i116_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i116_LC_7_19_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i116_LC_7_19_2  (
            .in0(N__33129),
            .in1(N__32057),
            .in2(N__26373),
            .in3(N__20613),
            .lcout(\c0.data_in_field_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37507),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i34_LC_7_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i34_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i34_LC_7_19_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i34_LC_7_19_3  (
            .in0(N__18910),
            .in1(N__23181),
            .in2(N__32216),
            .in3(N__33135),
            .lcout(\c0.data_in_field_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37507),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_893_LC_7_19_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_893_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_893_LC_7_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_893_LC_7_19_4  (
            .in0(N__19190),
            .in1(N__18909),
            .in2(_gnd_net_),
            .in3(N__27952),
            .lcout(\c0.n5403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_892_LC_7_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_892_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_892_LC_7_19_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_892_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__18876),
            .in2(_gnd_net_),
            .in3(N__22345),
            .lcout(\c0.n5391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i41_LC_7_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i41_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i41_LC_7_19_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i41_LC_7_19_6  (
            .in0(N__33130),
            .in1(N__32058),
            .in2(N__23523),
            .in3(N__26789),
            .lcout(\c0.data_in_field_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37507),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_982_LC_7_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_982_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_982_LC_7_19_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_982_LC_7_19_7  (
            .in0(N__27084),
            .in1(N__28058),
            .in2(N__18962),
            .in3(N__28122),
            .lcout(\c0.n5539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i93_LC_7_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i93_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i93_LC_7_20_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i93_LC_7_20_0  (
            .in0(N__33118),
            .in1(N__31932),
            .in2(N__24969),
            .in3(N__19191),
            .lcout(\c0.data_in_field_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i104_LC_7_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i104_LC_7_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i104_LC_7_20_1 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.data_in_frame_0___i104_LC_7_20_1  (
            .in0(N__18855),
            .in1(N__19136),
            .in2(N__32132),
            .in3(N__33120),
            .lcout(\c0.data_in_field_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_820_LC_7_20_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_820_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_820_LC_7_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_820_LC_7_20_2  (
            .in0(N__19116),
            .in1(N__18824),
            .in2(N__18792),
            .in3(N__18736),
            .lcout(\c0.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i19_LC_7_20_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i19_LC_7_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i19_LC_7_20_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i19_LC_7_20_3  (
            .in0(N__22044),
            .in1(_gnd_net_),
            .in2(N__35963),
            .in3(N__21485),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i134_LC_7_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i134_LC_7_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i134_LC_7_20_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i134_LC_7_20_4  (
            .in0(N__33117),
            .in1(N__31931),
            .in2(N__18702),
            .in3(N__27157),
            .lcout(\c0.data_in_field_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i53_LC_7_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i53_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i53_LC_7_20_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i53_LC_7_20_5  (
            .in0(N__31930),
            .in1(N__33119),
            .in2(N__23400),
            .in3(N__19163),
            .lcout(\c0.data_in_field_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37514),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_847_LC_7_20_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_847_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_847_LC_7_20_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_847_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__19132),
            .in2(_gnd_net_),
            .in3(N__27156),
            .lcout(\c0.n2152 ),
            .ltout(\c0.n2152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_849_LC_7_20_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_849_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_849_LC_7_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_849_LC_7_20_7  (
            .in0(N__23079),
            .in1(N__19105),
            .in2(N__19077),
            .in3(N__20739),
            .lcout(\c0.n5397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i30_LC_7_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i30_LC_7_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i30_LC_7_21_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i30_LC_7_21_0  (
            .in0(N__32090),
            .in1(N__19337),
            .in2(N__27900),
            .in3(N__32807),
            .lcout(\c0.data_in_field_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i95_LC_7_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i95_LC_7_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i95_LC_7_21_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i95_LC_7_21_1  (
            .in0(N__32805),
            .in1(N__32092),
            .in2(N__19053),
            .in3(N__21000),
            .lcout(\c0.data_in_field_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_905_LC_7_21_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_905_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_905_LC_7_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_905_LC_7_21_2  (
            .in0(N__23339),
            .in1(N__23306),
            .in2(_gnd_net_),
            .in3(N__19022),
            .lcout(\c0.n2065 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i143_LC_7_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i143_LC_7_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i143_LC_7_21_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i143_LC_7_21_3  (
            .in0(N__32804),
            .in1(N__32091),
            .in2(N__18990),
            .in3(N__18945),
            .lcout(\c0.data_in_field_142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i144_LC_7_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i144_LC_7_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i144_LC_7_21_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i144_LC_7_21_4  (
            .in0(N__27071),
            .in1(N__23109),
            .in2(N__32221),
            .in3(N__32806),
            .lcout(\c0.data_in_field_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37525),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_field_143__I_0_1808_2_lut_LC_7_21_5 .C_ON=1'b0;
    defparam \c0.data_in_field_143__I_0_1808_2_lut_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.data_in_field_143__I_0_1808_2_lut_LC_7_21_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_in_field_143__I_0_1808_2_lut_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__18944),
            .in2(_gnd_net_),
            .in3(N__27070),
            .lcout(),
            .ltout(\c0.tx2_transmit_N_1031_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_927_LC_7_21_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_927_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_927_LC_7_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_927_LC_7_21_6  (
            .in0(N__20163),
            .in1(N__25144),
            .in2(N__19341),
            .in3(N__19336),
            .lcout(\c0.n2030 ),
            .ltout(\c0.n2030_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_7_21_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_7_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_7_21_7  (
            .in0(N__20576),
            .in1(N__22235),
            .in2(N__19314),
            .in3(N__22649),
            .lcout(\c0.n5466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i23_LC_7_22_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i23_LC_7_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i23_LC_7_22_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i23_LC_7_22_0  (
            .in0(N__32084),
            .in1(N__19274),
            .in2(N__27815),
            .in3(N__33124),
            .lcout(\c0.data_in_field_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37538),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i123_LC_7_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i123_LC_7_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i123_LC_7_22_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i123_LC_7_22_1  (
            .in0(N__33121),
            .in1(N__32086),
            .in2(N__24603),
            .in3(N__19311),
            .lcout(\c0.data_in_field_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37538),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i83_LC_7_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i83_LC_7_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i83_LC_7_22_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i83_LC_7_22_2  (
            .in0(N__32085),
            .in1(N__33123),
            .in2(N__30678),
            .in3(N__19582),
            .lcout(\c0.data_in_field_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37538),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_914_LC_7_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_914_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_914_LC_7_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_914_LC_7_22_3  (
            .in0(N__19273),
            .in1(N__19616),
            .in2(_gnd_net_),
            .in3(N__20977),
            .lcout(\c0.n5436 ),
            .ltout(\c0.n5436_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_900_LC_7_22_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_900_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_900_LC_7_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_900_LC_7_22_4  (
            .in0(_gnd_net_),
            .in1(N__19549),
            .in2(N__19248),
            .in3(N__21440),
            .lcout(\c0.n5509 ),
            .ltout(\c0.n5509_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_874_LC_7_22_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_874_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_874_LC_7_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_874_LC_7_22_5  (
            .in0(_gnd_net_),
            .in1(N__19235),
            .in2(N__19212),
            .in3(N__19208),
            .lcout(\c0.n2053 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_918_LC_7_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_918_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_918_LC_7_22_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_918_LC_7_22_6  (
            .in0(N__20978),
            .in1(_gnd_net_),
            .in2(N__21568),
            .in3(_gnd_net_),
            .lcout(\c0.n1779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i37_LC_7_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i37_LC_7_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i37_LC_7_22_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i37_LC_7_22_7  (
            .in0(N__33122),
            .in1(N__32087),
            .in2(N__31230),
            .in3(N__19617),
            .lcout(\c0.data_in_field_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37538),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i117_LC_7_23_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i117_LC_7_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i117_LC_7_23_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i117_LC_7_23_0  (
            .in0(N__31936),
            .in1(N__32760),
            .in2(N__21572),
            .in3(N__26925),
            .lcout(\c0.data_in_field_116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_917_LC_7_23_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_917_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_917_LC_7_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_917_LC_7_23_1  (
            .in0(N__19575),
            .in1(N__19860),
            .in2(_gnd_net_),
            .in3(N__20780),
            .lcout(\c0.n1948 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i114_LC_7_23_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i114_LC_7_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i114_LC_7_23_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i114_LC_7_23_2  (
            .in0(N__35812),
            .in1(N__19486),
            .in2(_gnd_net_),
            .in3(N__19533),
            .lcout(data_in_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i19_LC_7_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i19_LC_7_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i19_LC_7_23_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i19_LC_7_23_4  (
            .in0(N__31937),
            .in1(N__22054),
            .in2(N__23020),
            .in3(N__32761),
            .lcout(\c0.data_in_field_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i128_LC_7_23_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i128_LC_7_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i128_LC_7_23_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i128_LC_7_23_5  (
            .in0(N__32759),
            .in1(N__31939),
            .in2(N__21876),
            .in3(N__19468),
            .lcout(\c0.data_in_field_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_23_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_23_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_7_23_6  (
            .in0(N__19439),
            .in1(N__20364),
            .in2(N__25496),
            .in3(N__20094),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i106_LC_7_23_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i106_LC_7_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i106_LC_7_23_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i106_LC_7_23_7  (
            .in0(N__32758),
            .in1(N__31938),
            .in2(N__19416),
            .in3(N__19376),
            .lcout(\c0.data_in_field_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37548),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_824_LC_7_24_0 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_824_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_824_LC_7_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_824_LC_7_24_0  (
            .in0(N__19362),
            .in1(N__27326),
            .in2(N__20124),
            .in3(N__25464),
            .lcout(\c0.n20_adj_1888 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i98_LC_7_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i98_LC_7_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i98_LC_7_24_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i98_LC_7_24_2  (
            .in0(N__31940),
            .in1(N__32970),
            .in2(N__19905),
            .in3(N__19869),
            .lcout(\c0.data_in_field_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i153_LC_7_24_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i153_LC_7_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i153_LC_7_24_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i153_LC_7_24_3  (
            .in0(N__21895),
            .in1(N__19923),
            .in2(_gnd_net_),
            .in3(N__35516),
            .lcout(data_in_19_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i113_LC_7_24_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i113_LC_7_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i113_LC_7_24_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i113_LC_7_24_6  (
            .in0(N__35515),
            .in1(N__19687),
            .in2(_gnd_net_),
            .in3(N__35069),
            .lcout(data_in_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i97_LC_7_24_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i97_LC_7_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i97_LC_7_24_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i97_LC_7_24_7  (
            .in0(N__32969),
            .in1(N__31941),
            .in2(N__20802),
            .in3(N__25760),
            .lcout(\c0.data_in_field_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37558),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i158_LC_7_25_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i158_LC_7_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i158_LC_7_25_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i158_LC_7_25_0  (
            .in0(N__19832),
            .in1(N__19730),
            .in2(N__33136),
            .in3(N__31943),
            .lcout(\c0.data_in_frame_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37568),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i111_LC_7_25_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i111_LC_7_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i111_LC_7_25_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i111_LC_7_25_3  (
            .in0(N__35629),
            .in1(N__19814),
            .in2(_gnd_net_),
            .in3(N__22916),
            .lcout(data_in_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37568),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i160_LC_7_25_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i160_LC_7_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i160_LC_7_25_4 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.data_in_frame_0___i160_LC_7_25_4  (
            .in0(N__19745),
            .in1(N__31942),
            .in2(N__33137),
            .in3(N__19782),
            .lcout(\c0.data_in_frame_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37568),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i150_LC_7_25_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i150_LC_7_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i150_LC_7_25_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i150_LC_7_25_6  (
            .in0(N__35518),
            .in1(N__21381),
            .in2(_gnd_net_),
            .in3(N__19729),
            .lcout(data_in_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37568),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i105_LC_7_25_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i105_LC_7_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i105_LC_7_25_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i105_LC_7_25_7  (
            .in0(N__35628),
            .in1(N__19688),
            .in2(_gnd_net_),
            .in3(N__19657),
            .lcout(data_in_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37568),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_LC_7_26_0 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_LC_7_26_0 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \c0.tx.i2_4_lut_LC_7_26_0  (
            .in0(N__29200),
            .in1(N__29115),
            .in2(N__29022),
            .in3(N__28495),
            .lcout(\c0.tx.n2247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i149_LC_7_26_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i149_LC_7_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i149_LC_7_26_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i149_LC_7_26_3  (
            .in0(N__35517),
            .in1(N__20118),
            .in2(_gnd_net_),
            .in3(N__20653),
            .lcout(data_in_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37576),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_7_26_4 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_7_26_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx.i1_2_lut_LC_7_26_4  (
            .in0(_gnd_net_),
            .in1(N__33868),
            .in2(_gnd_net_),
            .in3(N__29238),
            .lcout(),
            .ltout(\c0.tx.n40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2105_4_lut_LC_7_26_5 .C_ON=1'b0;
    defparam \c0.tx.i2105_4_lut_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2105_4_lut_LC_7_26_5 .LUT_INIT=16'b1100010001000100;
    LogicCell40 \c0.tx.i2105_4_lut_LC_7_26_5  (
            .in0(N__29116),
            .in1(N__20066),
            .in2(N__20097),
            .in3(N__29327),
            .lcout(\c0.tx.n2356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_792_LC_7_26_7 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_792_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_792_LC_7_26_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.i1_2_lut_adj_792_LC_7_26_7  (
            .in0(N__20403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19956),
            .lcout(n1760),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_7_27_0 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_7_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_7_27_0 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_7_27_0  (
            .in0(N__29334),
            .in1(_gnd_net_),
            .in2(N__33884),
            .in3(N__29239),
            .lcout(\c0.tx.r_Bit_Index_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37582),
            .ce(N__20073),
            .sr(N__20055));
    defparam \c0.tx.r_Bit_Index_i1_LC_7_27_1 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_7_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_7_27_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_7_27_1  (
            .in0(_gnd_net_),
            .in1(N__33869),
            .in2(_gnd_net_),
            .in3(N__29333),
            .lcout(\c0.tx.r_Bit_Index_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37582),
            .ce(N__20073),
            .sr(N__20055));
    defparam \c0.tx.i1_2_lut_3_lut_4_lut_LC_7_28_4 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_3_lut_4_lut_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_3_lut_4_lut_LC_7_28_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx.i1_2_lut_3_lut_4_lut_LC_7_28_4  (
            .in0(N__29005),
            .in1(N__29203),
            .in2(N__28617),
            .in3(N__29121),
            .lcout(n1519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_LC_7_28_6 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_LC_7_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_LC_7_28_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.rx.i2_3_lut_LC_7_28_6  (
            .in0(N__20049),
            .in1(N__19997),
            .in2(_gnd_net_),
            .in3(N__19952),
            .lcout(n1757),
            .ltout(n1757_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_7_28_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_7_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_7_28_7 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_7_28_7  (
            .in0(N__19916),
            .in1(N__20412),
            .in2(N__19926),
            .in3(N__20363),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37591),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_7_29_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_7_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_7_29_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_7_29_0  (
            .in0(N__20418),
            .in1(N__20362),
            .in2(N__26390),
            .in3(N__20256),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37597),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i6_LC_9_15_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i6_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i6_LC_9_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i6_LC_9_15_3  (
            .in0(N__35557),
            .in1(N__25058),
            .in2(_gnd_net_),
            .in3(N__20201),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37526),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i47_LC_9_16_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i47_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i47_LC_9_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i47_LC_9_16_1  (
            .in0(N__35406),
            .in1(N__24210),
            .in2(_gnd_net_),
            .in3(N__23353),
            .lcout(data_in_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37515),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i31_LC_9_16_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i31_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i31_LC_9_16_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i31_LC_9_16_3  (
            .in0(N__30629),
            .in1(_gnd_net_),
            .in2(N__35558),
            .in3(N__20235),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37515),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i39_LC_9_16_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i39_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i39_LC_9_16_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i39_LC_9_16_4  (
            .in0(N__23354),
            .in1(N__35405),
            .in2(_gnd_net_),
            .in3(N__30628),
            .lcout(data_in_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37515),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_LC_9_16_6 .C_ON=1'b0;
    defparam \c0.i6_2_lut_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_LC_9_16_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i6_2_lut_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__20200),
            .in2(_gnd_net_),
            .in3(N__22005),
            .lcout(\c0.n22_adj_1924 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i63_LC_9_16_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i63_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i63_LC_9_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i63_LC_9_16_7  (
            .in0(N__35407),
            .in1(N__31170),
            .in2(_gnd_net_),
            .in3(N__24226),
            .lcout(data_in_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37515),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i142_LC_9_17_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i142_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i142_LC_9_17_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i142_LC_9_17_0  (
            .in0(N__32122),
            .in1(N__33157),
            .in2(N__21354),
            .in3(N__20150),
            .lcout(\c0.data_in_field_141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37499),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_928_LC_9_17_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_928_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_928_LC_9_17_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_928_LC_9_17_1  (
            .in0(N__22222),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22637),
            .lcout(\c0.n5590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_949_LC_9_17_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_949_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_949_LC_9_17_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_949_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__28299),
            .in2(_gnd_net_),
            .in3(N__24861),
            .lcout(),
            .ltout(\c0.n5394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_825_LC_9_17_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_825_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_825_LC_9_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_825_LC_9_17_3  (
            .in0(N__29445),
            .in1(N__20499),
            .in2(N__20478),
            .in3(N__20475),
            .lcout(\c0.n19_adj_1889 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_821_LC_9_17_5 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_821_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_821_LC_9_17_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_821_LC_9_17_5  (
            .in0(N__20891),
            .in1(N__22194),
            .in2(N__20430),
            .in3(N__22170),
            .lcout(\c0.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i118_LC_9_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i118_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i118_LC_9_17_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i118_LC_9_17_7  (
            .in0(N__33156),
            .in1(N__32123),
            .in2(N__31311),
            .in3(N__22195),
            .lcout(\c0.data_in_field_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37499),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i56_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i56_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i56_LC_9_18_0 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i56_LC_9_18_0  (
            .in0(N__33095),
            .in1(N__32205),
            .in2(N__21080),
            .in3(N__26986),
            .lcout(\c0.data_in_field_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i35_LC_9_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i35_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i35_LC_9_18_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i35_LC_9_18_1  (
            .in0(N__32203),
            .in1(N__33097),
            .in2(N__21423),
            .in3(N__20543),
            .lcout(\c0.data_in_field_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i133_LC_9_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i133_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i133_LC_9_18_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i133_LC_9_18_2  (
            .in0(N__33094),
            .in1(N__32204),
            .in2(N__30351),
            .in3(N__20714),
            .lcout(\c0.data_in_field_132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_961_LC_9_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_961_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_961_LC_9_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_961_LC_9_18_3  (
            .in0(N__30829),
            .in1(N__31416),
            .in2(N__26990),
            .in3(N__30892),
            .lcout(\c0.n5515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_828_LC_9_18_4 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_828_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_828_LC_9_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_828_LC_9_18_4  (
            .in0(N__26982),
            .in1(N__23622),
            .in2(N__21915),
            .in3(N__21771),
            .lcout(),
            .ltout(\c0.n40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_LC_9_18_5 .C_ON=1'b0;
    defparam \c0.i23_4_lut_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_LC_9_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i23_4_lut_LC_9_18_5  (
            .in0(N__20760),
            .in1(N__21267),
            .in2(N__20754),
            .in3(N__20751),
            .lcout(\c0.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i61_LC_9_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i61_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i61_LC_9_18_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i61_LC_9_18_6  (
            .in0(N__33096),
            .in1(N__32206),
            .in2(N__23427),
            .in3(N__22642),
            .lcout(\c0.data_in_field_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37516),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_861_LC_9_18_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_861_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_861_LC_9_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_861_LC_9_18_7  (
            .in0(N__20713),
            .in1(N__21680),
            .in2(_gnd_net_),
            .in3(N__20542),
            .lcout(\c0.n1969 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_895_LC_9_19_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_895_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_895_LC_9_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_895_LC_9_19_0  (
            .in0(N__24380),
            .in1(N__20675),
            .in2(_gnd_net_),
            .in3(N__25105),
            .lcout(\c0.n1855 ),
            .ltout(\c0.n1855_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_832_LC_9_19_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_832_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_832_LC_9_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_832_LC_9_19_1  (
            .in0(N__20661),
            .in1(N__20615),
            .in2(N__20586),
            .in3(N__20583),
            .lcout(\c0.n13_adj_1899 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i21_LC_9_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i21_LC_9_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i21_LC_9_19_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0___i21_LC_9_19_2  (
            .in0(N__31104),
            .in1(N__32172),
            .in2(N__21698),
            .in3(N__33271),
            .lcout(\c0.data_in_field_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37527),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i25_LC_9_19_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i25_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i25_LC_9_19_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i25_LC_9_19_3  (
            .in0(N__35853),
            .in1(N__23492),
            .in2(_gnd_net_),
            .in3(N__27843),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37527),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i69_LC_9_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i69_LC_9_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i69_LC_9_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i69_LC_9_19_4  (
            .in0(N__35401),
            .in1(N__30386),
            .in2(_gnd_net_),
            .in3(N__23449),
            .lcout(data_in_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37527),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_962_LC_9_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_962_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_962_LC_9_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_962_LC_9_19_5  (
            .in0(N__22574),
            .in1(N__22529),
            .in2(N__25984),
            .in3(N__20541),
            .lcout(\c0.n2092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i140_LC_9_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i140_LC_9_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i140_LC_9_19_6 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i140_LC_9_19_6  (
            .in0(N__22530),
            .in1(N__33270),
            .in2(N__21135),
            .in3(N__32173),
            .lcout(\c0.data_in_field_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37527),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i20_LC_9_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i20_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i20_LC_9_19_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i20_LC_9_19_7  (
            .in0(N__33269),
            .in1(N__22582),
            .in2(N__21111),
            .in3(N__32126),
            .lcout(\c0.data_in_field_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37527),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i48_LC_9_20_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i48_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i48_LC_9_20_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i48_LC_9_20_0  (
            .in0(N__35904),
            .in1(N__21081),
            .in2(_gnd_net_),
            .in3(N__27181),
            .lcout(data_in_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37539),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i46_LC_9_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i46_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i46_LC_9_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i46_LC_9_20_1  (
            .in0(N__35901),
            .in1(N__21044),
            .in2(_gnd_net_),
            .in3(N__22501),
            .lcout(data_in_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37539),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i45_LC_9_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i45_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i45_LC_9_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i45_LC_9_20_2  (
            .in0(N__23396),
            .in1(N__35902),
            .in2(_gnd_net_),
            .in3(N__27343),
            .lcout(data_in_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37539),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_957_LC_9_20_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_957_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_957_LC_9_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_957_LC_9_20_3  (
            .in0(N__22091),
            .in1(N__31102),
            .in2(N__22278),
            .in3(N__21478),
            .lcout(\c0.n25_adj_1948 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_911_LC_9_20_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_911_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_911_LC_9_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_911_LC_9_20_4  (
            .in0(N__21002),
            .in1(N__20951),
            .in2(_gnd_net_),
            .in3(N__20923),
            .lcout(\c0.n5545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_979_LC_9_20_6 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_979_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_979_LC_9_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_979_LC_9_20_6  (
            .in0(N__21273),
            .in1(N__22725),
            .in2(N__30734),
            .in3(N__23655),
            .lcout(\c0.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_907_LC_9_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_907_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_907_LC_9_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_907_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__20858),
            .in2(_gnd_net_),
            .in3(N__20810),
            .lcout(\c0.n5427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_LC_9_21_0 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_LC_9_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_3_lut_4_lut_LC_9_21_0  (
            .in0(N__21809),
            .in1(N__21539),
            .in2(N__25455),
            .in3(N__28114),
            .lcout(\c0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i94_LC_9_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i94_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i94_LC_9_21_1 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i94_LC_9_21_1  (
            .in0(N__25104),
            .in1(N__32006),
            .in2(N__27021),
            .in3(N__32895),
            .lcout(\c0.data_in_field_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37549),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i118_LC_9_21_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i118_LC_9_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i118_LC_9_21_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i118_LC_9_21_2  (
            .in0(N__31297),
            .in1(N__35903),
            .in2(_gnd_net_),
            .in3(N__21308),
            .lcout(data_in_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37549),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_rep_100_2_lut_3_lut_LC_9_21_3 .C_ON=1'b0;
    defparam \c0.i1_rep_100_2_lut_3_lut_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_rep_100_2_lut_3_lut_LC_9_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_rep_100_2_lut_3_lut_LC_9_21_3  (
            .in0(N__21209),
            .in1(N__26642),
            .in2(_gnd_net_),
            .in3(N__21179),
            .lcout(\c0.n6414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_853_LC_9_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_853_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_853_LC_9_21_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_853_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__21808),
            .in2(_gnd_net_),
            .in3(N__21538),
            .lcout(\c0.n5563 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i46_LC_9_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i46_LC_9_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i46_LC_9_21_5 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i46_LC_9_21_5  (
            .in0(N__21210),
            .in1(N__32894),
            .in2(N__22506),
            .in3(N__32007),
            .lcout(\c0.data_in_field_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37549),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i90_LC_9_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i90_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i90_LC_9_21_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i90_LC_9_21_6  (
            .in0(N__32005),
            .in1(N__33227),
            .in2(N__21258),
            .in3(N__23338),
            .lcout(\c0.data_in_field_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37549),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_952_LC_9_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_952_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_952_LC_9_22_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_952_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__21211),
            .in2(_gnd_net_),
            .in3(N__26643),
            .lcout(),
            .ltout(\c0.n2149_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_9_22_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_9_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_LC_9_22_1  (
            .in0(N__21183),
            .in1(N__21156),
            .in2(N__21150),
            .in3(N__22608),
            .lcout(\c0.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i27_LC_9_22_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i27_LC_9_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i27_LC_9_22_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i27_LC_9_22_3  (
            .in0(N__36054),
            .in1(N__21413),
            .in2(_gnd_net_),
            .in3(N__21471),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37559),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_899_LC_9_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_899_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_899_LC_9_22_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_899_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__25094),
            .in2(_gnd_net_),
            .in3(N__23221),
            .lcout(\c0.n1955 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i35_LC_9_22_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i35_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i35_LC_9_22_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i35_LC_9_22_5  (
            .in0(N__36055),
            .in1(N__21412),
            .in2(_gnd_net_),
            .in3(N__25628),
            .lcout(data_in_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37559),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i142_LC_9_22_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i142_LC_9_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i142_LC_9_22_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i142_LC_9_22_7  (
            .in0(N__36053),
            .in1(N__21340),
            .in2(_gnd_net_),
            .in3(N__21395),
            .lcout(data_in_17_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37559),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i0_LC_9_23_0 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i0_LC_9_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i0_LC_9_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i0_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__23549),
            .in2(N__36792),
            .in3(_gnd_net_),
            .lcout(\c0.delay_counter_0 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\c0.n4754 ),
            .clk(N__37569),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i1_LC_9_23_1 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i1_LC_9_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i1_LC_9_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i1_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__21597),
            .in2(_gnd_net_),
            .in3(N__21324),
            .lcout(\c0.delay_counter_1 ),
            .ltout(),
            .carryin(\c0.n4754 ),
            .carryout(\c0.n4755 ),
            .clk(N__37569),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i2_LC_9_23_2 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i2_LC_9_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i2_LC_9_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i2_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__23562),
            .in2(_gnd_net_),
            .in3(N__21321),
            .lcout(\c0.delay_counter_2 ),
            .ltout(),
            .carryin(\c0.n4755 ),
            .carryout(\c0.n4756 ),
            .clk(N__37569),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i3_LC_9_23_3 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i3_LC_9_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i3_LC_9_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i3_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__26099),
            .in2(_gnd_net_),
            .in3(N__21318),
            .lcout(\c0.delay_counter_3 ),
            .ltout(),
            .carryin(\c0.n4756 ),
            .carryout(\c0.n4757 ),
            .clk(N__37569),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i4_LC_9_23_4 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i4_LC_9_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i4_LC_9_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i4_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__26021),
            .in2(_gnd_net_),
            .in3(N__21315),
            .lcout(\c0.delay_counter_4 ),
            .ltout(),
            .carryin(\c0.n4757 ),
            .carryout(\c0.n4758 ),
            .clk(N__37569),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i5_LC_9_23_5 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i5_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i5_LC_9_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i5_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__21585),
            .in2(_gnd_net_),
            .in3(N__21312),
            .lcout(\c0.delay_counter_5 ),
            .ltout(),
            .carryin(\c0.n4758 ),
            .carryout(\c0.n4759 ),
            .clk(N__37569),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i6_LC_9_23_6 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i6_LC_9_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i6_LC_9_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i6_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__26081),
            .in2(_gnd_net_),
            .in3(N__21612),
            .lcout(\c0.delay_counter_6 ),
            .ltout(),
            .carryin(\c0.n4759 ),
            .carryout(\c0.n4760 ),
            .clk(N__37569),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i7_LC_9_23_7 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i7_LC_9_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i7_LC_9_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i7_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__23535),
            .in2(_gnd_net_),
            .in3(N__21609),
            .lcout(\c0.delay_counter_7 ),
            .ltout(),
            .carryin(\c0.n4760 ),
            .carryout(\c0.n4761 ),
            .clk(N__37569),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i8_LC_9_24_0 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i8_LC_9_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i8_LC_9_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i8_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__26039),
            .in2(_gnd_net_),
            .in3(N__21606),
            .lcout(\c0.delay_counter_8 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\c0.n4762 ),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i9_LC_9_24_1 .C_ON=1'b1;
    defparam \c0.delay_counter_528__i9_LC_9_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i9_LC_9_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_528__i9_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__23574),
            .in2(_gnd_net_),
            .in3(N__21603),
            .lcout(\c0.delay_counter_9 ),
            .ltout(),
            .carryin(\c0.n4762 ),
            .carryout(\c0.n4763 ),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_528__i10_LC_9_24_2 .C_ON=1'b0;
    defparam \c0.delay_counter_528__i10_LC_9_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_528__i10_LC_9_24_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.delay_counter_528__i10_LC_9_24_2  (
            .in0(N__26063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21600),
            .lcout(\c0.delay_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37577),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_LC_9_24_3 .C_ON=1'b0;
    defparam \c0.i5_2_lut_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_LC_9_24_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i5_2_lut_LC_9_24_3  (
            .in0(N__21596),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21584),
            .lcout(\c0.n16_adj_1921 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5799_LC_9_24_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5799_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5799_LC_9_24_5 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5799_LC_9_24_5  (
            .in0(N__27703),
            .in1(N__21573),
            .in2(N__30173),
            .in3(N__21543),
            .lcout(),
            .ltout(\c0.n6171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6171_bdd_4_lut_LC_9_24_6 .C_ON=1'b0;
    defparam \c0.n6171_bdd_4_lut_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.n6171_bdd_4_lut_LC_9_24_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6171_bdd_4_lut_LC_9_24_6  (
            .in0(N__30113),
            .in1(N__30260),
            .in2(N__21504),
            .in3(N__24869),
            .lcout(\c0.n5731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6189_bdd_4_lut_LC_9_25_0 .C_ON=1'b0;
    defparam \c0.n6189_bdd_4_lut_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.n6189_bdd_4_lut_LC_9_25_0 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n6189_bdd_4_lut_LC_9_25_0  (
            .in0(N__30100),
            .in1(N__21813),
            .in2(N__21657),
            .in3(N__21770),
            .lcout(\c0.n5722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i3388_2_lut_LC_9_25_1 .C_ON=1'b0;
    defparam \c0.tx.i3388_2_lut_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i3388_2_lut_LC_9_25_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i3388_2_lut_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__29017),
            .in2(_gnd_net_),
            .in3(N__29092),
            .lcout(),
            .ltout(\c0.tx.n3631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5592_3_lut_4_lut_LC_9_25_2 .C_ON=1'b0;
    defparam \c0.tx.i5592_3_lut_4_lut_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5592_3_lut_4_lut_LC_9_25_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.tx.i5592_3_lut_4_lut_LC_9_25_2  (
            .in0(N__28609),
            .in1(N__29173),
            .in2(N__21702),
            .in3(N__23807),
            .lcout(\c0.tx.n5883 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_9_25_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_9_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_9_25_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_9_25_3  (
            .in0(N__23727),
            .in1(N__33605),
            .in2(_gnd_net_),
            .in3(N__21624),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i17_LC_9_25_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i17_LC_9_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i17_LC_9_25_7 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \c0.data_out_0___i17_LC_9_25_7  (
            .in0(N__28725),
            .in1(N__23847),
            .in2(N__36183),
            .in3(N__37727),
            .lcout(data_out_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37583),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5819_LC_9_26_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5819_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5819_LC_9_26_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5819_LC_9_26_1  (
            .in0(N__27612),
            .in1(N__28238),
            .in2(N__30174),
            .in3(N__21697),
            .lcout(\c0.n6189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5604_2_lut_3_lut_LC_9_26_4 .C_ON=1'b0;
    defparam \c0.tx.i5604_2_lut_3_lut_LC_9_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5604_2_lut_3_lut_LC_9_26_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.tx.i5604_2_lut_3_lut_LC_9_26_4  (
            .in0(N__28477),
            .in1(_gnd_net_),
            .in2(N__29253),
            .in3(N__33888),
            .lcout(),
            .ltout(\c0.tx.n5812_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i28_4_lut_LC_9_26_5 .C_ON=1'b0;
    defparam \c0.tx.i28_4_lut_LC_9_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i28_4_lut_LC_9_26_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \c0.tx.i28_4_lut_LC_9_26_5  (
            .in0(N__28613),
            .in1(N__29089),
            .in2(N__21648),
            .in3(N__29326),
            .lcout(),
            .ltout(\c0.tx.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_9_26_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_9_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_9_26_6 .LUT_INIT=16'b0001000100110000;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_9_26_6  (
            .in0(N__28478),
            .in1(N__29016),
            .in2(N__21645),
            .in3(N__29175),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37592),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_26_7 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_26_7 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx.r_Bit_Index_0__bdd_4_lut_LC_9_26_7  (
            .in0(N__21642),
            .in1(N__21623),
            .in2(N__33893),
            .in3(N__29325),
            .lcout(\c0.tx.n6285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_2_lut_LC_9_27_0 .C_ON=1'b1;
    defparam \c0.tx.add_59_2_lut_LC_9_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_2_lut_LC_9_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_2_lut_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__26499),
            .in2(_gnd_net_),
            .in3(N__21840),
            .lcout(n321),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\c0.tx.n4764 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_3_lut_LC_9_27_1 .C_ON=1'b1;
    defparam \c0.tx.add_59_3_lut_LC_9_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_3_lut_LC_9_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_3_lut_LC_9_27_1  (
            .in0(_gnd_net_),
            .in1(N__26421),
            .in2(_gnd_net_),
            .in3(N__21837),
            .lcout(n320),
            .ltout(),
            .carryin(\c0.tx.n4764 ),
            .carryout(\c0.tx.n4765 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_4_lut_LC_9_27_2 .C_ON=1'b1;
    defparam \c0.tx.add_59_4_lut_LC_9_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_4_lut_LC_9_27_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_4_lut_LC_9_27_2  (
            .in0(N__22134),
            .in1(N__23977),
            .in2(_gnd_net_),
            .in3(N__21834),
            .lcout(\c0.tx.n5885 ),
            .ltout(),
            .carryin(\c0.tx.n4765 ),
            .carryout(\c0.tx.n4766 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_5_lut_LC_9_27_3 .C_ON=1'b1;
    defparam \c0.tx.add_59_5_lut_LC_9_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_5_lut_LC_9_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_5_lut_LC_9_27_3  (
            .in0(_gnd_net_),
            .in1(N__26538),
            .in2(_gnd_net_),
            .in3(N__21831),
            .lcout(n318),
            .ltout(),
            .carryin(\c0.tx.n4766 ),
            .carryout(\c0.tx.n4767 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_6_lut_LC_9_27_4 .C_ON=1'b1;
    defparam \c0.tx.add_59_6_lut_LC_9_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_6_lut_LC_9_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_6_lut_LC_9_27_4  (
            .in0(_gnd_net_),
            .in1(N__24068),
            .in2(_gnd_net_),
            .in3(N__21828),
            .lcout(n317),
            .ltout(),
            .carryin(\c0.tx.n4767 ),
            .carryout(\c0.tx.n4768 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_7_lut_LC_9_27_5 .C_ON=1'b1;
    defparam \c0.tx.add_59_7_lut_LC_9_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_7_lut_LC_9_27_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_7_lut_LC_9_27_5  (
            .in0(N__23997),
            .in1(N__23781),
            .in2(_gnd_net_),
            .in3(N__21825),
            .lcout(\c0.tx.n5821 ),
            .ltout(),
            .carryin(\c0.tx.n4768 ),
            .carryout(\c0.tx.n4769 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_8_lut_LC_9_27_6 .C_ON=1'b1;
    defparam \c0.tx.add_59_8_lut_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_8_lut_LC_9_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_8_lut_LC_9_27_6  (
            .in0(_gnd_net_),
            .in1(N__24099),
            .in2(_gnd_net_),
            .in3(N__21822),
            .lcout(n315),
            .ltout(),
            .carryin(\c0.tx.n4769 ),
            .carryout(\c0.tx.n4770 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_9_lut_LC_9_27_7 .C_ON=1'b1;
    defparam \c0.tx.add_59_9_lut_LC_9_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_9_lut_LC_9_27_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_9_lut_LC_9_27_7  (
            .in0(N__22133),
            .in1(N__24037),
            .in2(_gnd_net_),
            .in3(N__21819),
            .lcout(\c0.tx.n5884 ),
            .ltout(),
            .carryin(\c0.tx.n4770 ),
            .carryout(\c0.tx.n4771 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_10_lut_LC_9_28_0 .C_ON=1'b0;
    defparam \c0.tx.add_59_10_lut_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_10_lut_LC_9_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx.add_59_10_lut_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(N__23930),
            .in2(_gnd_net_),
            .in3(N__21816),
            .lcout(n313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i2_LC_9_28_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i2_LC_9_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_9_28_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_9_28_3  (
            .in0(N__23979),
            .in1(N__29010),
            .in2(_gnd_net_),
            .in3(N__22140),
            .lcout(\c0.tx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37603),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i33_3_lut_LC_9_28_4 .C_ON=1'b0;
    defparam \c0.tx.i33_3_lut_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i33_3_lut_LC_9_28_4 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \c0.tx.i33_3_lut_LC_9_28_4  (
            .in0(N__29009),
            .in1(N__23978),
            .in2(_gnd_net_),
            .in3(N__23996),
            .lcout(\c0.tx.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i7_LC_9_28_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i7_LC_9_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_9_28_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_9_28_5  (
            .in0(N__24038),
            .in1(N__29011),
            .in2(_gnd_net_),
            .in3(N__22122),
            .lcout(\c0.tx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37603),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i28_LC_10_15_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i28_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i28_LC_10_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i28_LC_10_15_3  (
            .in0(N__35630),
            .in1(N__22115),
            .in2(_gnd_net_),
            .in3(N__22077),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37529),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i11_LC_10_16_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i11_LC_10_16_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i11_LC_10_16_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i11_LC_10_16_4  (
            .in0(N__35978),
            .in1(N__22006),
            .in2(_gnd_net_),
            .in3(N__22056),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37518),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_977_LC_10_16_6 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_977_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_977_LC_10_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_977_LC_10_16_6  (
            .in0(N__26890),
            .in1(N__29503),
            .in2(N__23157),
            .in3(N__21983),
            .lcout(),
            .ltout(\c0.n42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_LC_10_16_7 .C_ON=1'b0;
    defparam \c0.i21_4_lut_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_LC_10_16_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i21_4_lut_LC_10_16_7  (
            .in0(N__24555),
            .in1(N__25835),
            .in2(N__21936),
            .in3(N__22589),
            .lcout(\c0.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i145_LC_10_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i145_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i145_LC_10_17_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i145_LC_10_17_0  (
            .in0(N__35688),
            .in1(N__24168),
            .in2(_gnd_net_),
            .in3(N__21914),
            .lcout(data_in_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i128_LC_10_17_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i128_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i128_LC_10_17_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i128_LC_10_17_1  (
            .in0(N__22415),
            .in1(N__35689),
            .in2(_gnd_net_),
            .in3(N__21853),
            .lcout(data_in_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i136_LC_10_17_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i136_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i136_LC_10_17_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i136_LC_10_17_2  (
            .in0(N__35687),
            .in1(N__22414),
            .in2(_gnd_net_),
            .in3(N__23102),
            .lcout(data_in_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_826_LC_10_17_3 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_826_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_826_LC_10_17_3 .LUT_INIT=16'b1111111101101001;
    LogicCell40 \c0.i6_4_lut_adj_826_LC_10_17_3  (
            .in0(N__22401),
            .in1(N__24390),
            .in2(N__22395),
            .in3(N__24246),
            .lcout(\c0.n22_adj_1890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_855_LC_10_17_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_855_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_855_LC_10_17_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_855_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__24528),
            .in2(_gnd_net_),
            .in3(N__22365),
            .lcout(\c0.n5384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i26_LC_10_17_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i26_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i26_LC_10_17_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i26_LC_10_17_6  (
            .in0(N__23180),
            .in1(_gnd_net_),
            .in2(N__35876),
            .in3(N__22300),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37508),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i1_LC_10_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i1_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i1_LC_10_18_0 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i1_LC_10_18_0  (
            .in0(N__22274),
            .in1(N__31997),
            .in2(N__33228),
            .in3(N__22228),
            .lcout(\c0.data_in_field_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i78_LC_10_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i78_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i78_LC_10_18_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i78_LC_10_18_1  (
            .in0(N__31996),
            .in1(N__33098),
            .in2(N__28824),
            .in3(N__25983),
            .lcout(\c0.data_in_field_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37519),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_LC_10_18_2 .C_ON=1'b0;
    defparam \c0.i4_3_lut_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_LC_10_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i4_3_lut_LC_10_18_2  (
            .in0(N__22188),
            .in1(N__23654),
            .in2(_gnd_net_),
            .in3(N__22166),
            .lcout(),
            .ltout(\c0.n12_adj_1898_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_830_LC_10_18_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_830_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_830_LC_10_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_830_LC_10_18_3  (
            .in0(N__22604),
            .in1(N__22155),
            .in2(N__22143),
            .in3(N__24135),
            .lcout(),
            .ltout(\c0.n5567_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_834_LC_10_18_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_834_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_834_LC_10_18_4 .LUT_INIT=16'b1001111101101111;
    LogicCell40 \c0.i1_4_lut_adj_834_LC_10_18_4  (
            .in0(N__22872),
            .in1(N__22860),
            .in2(N__22848),
            .in3(N__22845),
            .lcout(\c0.n17_adj_1902 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6219_bdd_4_lut_LC_10_18_5 .C_ON=1'b0;
    defparam \c0.n6219_bdd_4_lut_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.n6219_bdd_4_lut_LC_10_18_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n6219_bdd_4_lut_LC_10_18_5  (
            .in0(N__30200),
            .in1(N__25025),
            .in2(N__22839),
            .in3(N__22824),
            .lcout(\c0.n5707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_948_LC_10_19_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_948_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_948_LC_10_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_948_LC_10_19_0  (
            .in0(N__22794),
            .in1(N__22770),
            .in2(N__24999),
            .in3(N__22749),
            .lcout(\c0.n5506 ),
            .ltout(\c0.n5506_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_831_LC_10_19_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_831_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_831_LC_10_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_831_LC_10_19_1  (
            .in0(N__24477),
            .in1(N__22719),
            .in2(N__22698),
            .in3(N__22695),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1010_LC_10_19_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1010_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1010_LC_10_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1010_LC_10_19_2  (
            .in0(N__22673),
            .in1(N__28338),
            .in2(N__26859),
            .in3(N__22638),
            .lcout(\c0.n5500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_890_LC_10_19_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_890_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_890_LC_10_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_890_LC_10_19_3  (
            .in0(N__25982),
            .in1(N__22575),
            .in2(_gnd_net_),
            .in3(N__22531),
            .lcout(\c0.n5372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i38_LC_10_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i38_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i38_LC_10_19_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i38_LC_10_19_4  (
            .in0(N__35981),
            .in1(N__25583),
            .in2(_gnd_net_),
            .in3(N__22502),
            .lcout(data_in_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37530),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i42_LC_10_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i42_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i42_LC_10_19_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i42_LC_10_19_5  (
            .in0(N__22438),
            .in1(N__35983),
            .in2(_gnd_net_),
            .in3(N__22485),
            .lcout(data_in_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37530),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i34_LC_10_19_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i34_LC_10_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i34_LC_10_19_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i34_LC_10_19_7  (
            .in0(N__22439),
            .in1(N__35982),
            .in2(_gnd_net_),
            .in3(N__23173),
            .lcout(data_in_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37530),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i144_LC_10_20_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i144_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i144_LC_10_20_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i144_LC_10_20_0  (
            .in0(N__36052),
            .in1(N__23095),
            .in2(_gnd_net_),
            .in3(N__23149),
            .lcout(data_in_17_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37540),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_964_LC_10_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_964_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_964_LC_10_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_964_LC_10_20_1  (
            .in0(N__23675),
            .in1(N__25934),
            .in2(N__25454),
            .in3(N__25017),
            .lcout(\c0.n6_adj_1918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i13_LC_10_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i13_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i13_LC_10_20_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i13_LC_10_20_2  (
            .in0(N__31103),
            .in1(_gnd_net_),
            .in2(N__36073),
            .in3(N__23047),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37540),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_891_LC_10_20_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_891_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_891_LC_10_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_891_LC_10_20_3  (
            .in0(N__23676),
            .in1(N__25935),
            .in2(_gnd_net_),
            .in3(N__25018),
            .lcout(),
            .ltout(\c0.n2043_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_992_LC_10_20_4 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_992_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_992_LC_10_20_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_adj_992_LC_10_20_4  (
            .in0(N__23021),
            .in1(N__22977),
            .in2(N__22971),
            .in3(N__22967),
            .lcout(\c0.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i70_LC_10_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i70_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i70_LC_10_20_5 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i70_LC_10_20_5  (
            .in0(N__26580),
            .in1(N__33108),
            .in2(N__32171),
            .in3(N__25936),
            .lcout(\c0.data_in_field_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37540),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i111_LC_10_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i111_LC_10_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i111_LC_10_20_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0___i111_LC_10_20_6  (
            .in0(N__31994),
            .in1(N__23677),
            .in2(N__33229),
            .in3(N__22923),
            .lcout(\c0.data_in_field_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37540),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i102_LC_10_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i102_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i102_LC_10_20_7 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i102_LC_10_20_7  (
            .in0(N__25441),
            .in1(N__33107),
            .in2(N__34461),
            .in3(N__31995),
            .lcout(\c0.data_in_field_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37540),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_973_LC_10_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_973_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_973_LC_10_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_973_LC_10_21_0  (
            .in0(N__23298),
            .in1(N__26877),
            .in2(N__24521),
            .in3(N__26951),
            .lcout(\c0.n5443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i49_LC_10_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i49_LC_10_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i49_LC_10_21_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i49_LC_10_21_1  (
            .in0(N__26878),
            .in1(N__28800),
            .in2(N__32170),
            .in3(N__33241),
            .lcout(\c0.data_in_field_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i91_LC_10_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i91_LC_10_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i91_LC_10_21_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i91_LC_10_21_2  (
            .in0(N__23299),
            .in1(N__33005),
            .in2(N__31260),
            .in3(N__32004),
            .lcout(\c0.data_in_field_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_951_LC_10_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_951_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_951_LC_10_21_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_951_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__23331),
            .in2(_gnd_net_),
            .in3(N__23297),
            .lcout(\c0.n1866 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i64_LC_10_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i64_LC_10_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i64_LC_10_21_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i64_LC_10_21_4  (
            .in0(N__33238),
            .in1(N__32000),
            .in2(N__23277),
            .in3(N__26952),
            .lcout(\c0.data_in_field_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i63_LC_10_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i63_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i63_LC_10_21_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i63_LC_10_21_5  (
            .in0(N__31999),
            .in1(N__33240),
            .in2(N__24529),
            .in3(N__24240),
            .lcout(\c0.data_in_field_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i85_LC_10_21_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i85_LC_10_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i85_LC_10_21_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i85_LC_10_21_6  (
            .in0(N__36048),
            .in1(N__24959),
            .in2(_gnd_net_),
            .in3(N__30406),
            .lcout(data_in_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i29_LC_10_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i29_LC_10_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i29_LC_10_21_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i29_LC_10_21_7  (
            .in0(N__31998),
            .in1(N__33239),
            .in2(N__31137),
            .in3(N__28224),
            .lcout(\c0.data_in_field_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37550),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i38_LC_10_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i38_LC_10_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i38_LC_10_22_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i38_LC_10_22_1  (
            .in0(N__33125),
            .in1(N__32244),
            .in2(N__25599),
            .in3(N__23227),
            .lcout(\c0.data_in_field_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37560),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i145_LC_10_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i145_LC_10_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i145_LC_10_22_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0___i145_LC_10_22_3  (
            .in0(N__23195),
            .in1(N__24176),
            .in2(N__33232),
            .in3(N__32245),
            .lcout(\c0.data_in_frame_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37560),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_943_LC_10_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_943_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_943_LC_10_22_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_943_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__27986),
            .in2(_gnd_net_),
            .in3(N__24781),
            .lcout(\c0.n2077 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6195_bdd_4_lut_LC_10_22_6 .C_ON=1'b0;
    defparam \c0.n6195_bdd_4_lut_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.n6195_bdd_4_lut_LC_10_22_6 .LUT_INIT=16'b1111110000001010;
    LogicCell40 \c0.n6195_bdd_4_lut_LC_10_22_6  (
            .in0(N__23610),
            .in1(N__23598),
            .in2(N__25413),
            .in3(N__25158),
            .lcout(\c0.n6198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_852_LC_10_23_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_852_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_852_LC_10_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_852_LC_10_23_0  (
            .in0(N__23573),
            .in1(N__23561),
            .in2(N__23550),
            .in3(N__23534),
            .lcout(\c0.n18_adj_1919 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i41_LC_10_23_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i41_LC_10_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i41_LC_10_23_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i41_LC_10_23_1  (
            .in0(N__35816),
            .in1(N__28799),
            .in2(_gnd_net_),
            .in3(N__23509),
            .lcout(data_in_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i33_LC_10_23_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i33_LC_10_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i33_LC_10_23_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i33_LC_10_23_2  (
            .in0(N__23510),
            .in1(N__35819),
            .in2(_gnd_net_),
            .in3(N__23473),
            .lcout(data_in_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i61_LC_10_23_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i61_LC_10_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i61_LC_10_23_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i61_LC_10_23_3  (
            .in0(N__35818),
            .in1(N__23413),
            .in2(_gnd_net_),
            .in3(N__23456),
            .lcout(data_in_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i51_LC_10_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i51_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i51_LC_10_23_4 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i51_LC_10_23_4  (
            .in0(N__33231),
            .in1(N__32243),
            .in2(N__25662),
            .in3(N__24792),
            .lcout(\c0.data_in_field_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i53_LC_10_23_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i53_LC_10_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i53_LC_10_23_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i53_LC_10_23_5  (
            .in0(N__35817),
            .in1(N__23414),
            .in2(_gnd_net_),
            .in3(N__23383),
            .lcout(data_in_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i47_LC_10_23_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i47_LC_10_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i47_LC_10_23_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i47_LC_10_23_6  (
            .in0(N__33230),
            .in1(N__32242),
            .in2(N__23367),
            .in3(N__27994),
            .lcout(\c0.data_in_field_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37570),
            .ce(),
            .sr(_gnd_net_));
    defparam i5299_4_lut_LC_10_24_0.C_ON=1'b0;
    defparam i5299_4_lut_LC_10_24_0.SEQ_MODE=4'b0000;
    defparam i5299_4_lut_LC_10_24_0.LUT_INIT=16'b1011101100100000;
    LogicCell40 i5299_4_lut_LC_10_24_0 (
            .in0(N__34808),
            .in1(N__36230),
            .in2(N__36261),
            .in3(N__34835),
            .lcout(n5645),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5300_4_lut_LC_10_24_1.C_ON=1'b0;
    defparam i5300_4_lut_LC_10_24_1.SEQ_MODE=4'b0000;
    defparam i5300_4_lut_LC_10_24_1.LUT_INIT=16'b1110101011101100;
    LogicCell40 i5300_4_lut_LC_10_24_1 (
            .in0(N__34836),
            .in1(N__36260),
            .in2(N__36234),
            .in3(N__34809),
            .lcout(),
            .ltout(n5646_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5301_3_lut_LC_10_24_2.C_ON=1'b0;
    defparam i5301_3_lut_LC_10_24_2.SEQ_MODE=4'b0000;
    defparam i5301_3_lut_LC_10_24_2.LUT_INIT=16'b0000101001011111;
    LogicCell40 i5301_3_lut_LC_10_24_2 (
            .in0(N__36204),
            .in1(_gnd_net_),
            .in2(N__23721),
            .in3(N__23718),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i32_LC_10_24_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i32_LC_10_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i32_LC_10_24_4 .LUT_INIT=16'b1110101101000001;
    LogicCell40 \c0.data_out_0___i32_LC_10_24_4  (
            .in0(N__37717),
            .in1(N__28560),
            .in2(N__28713),
            .in3(N__26247),
            .lcout(data_out_19_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37578),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i23_LC_10_24_5 .C_ON=1'b0;
    defparam \c0.data_out_0___i23_LC_10_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i23_LC_10_24_5 .LUT_INIT=16'b1111000010011001;
    LogicCell40 \c0.data_out_0___i23_LC_10_24_5  (
            .in0(N__33669),
            .in1(N__34602),
            .in2(N__23637),
            .in3(N__37715),
            .lcout(data_out_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37578),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i25_LC_10_24_6 .C_ON=1'b0;
    defparam \c0.data_out_0___i25_LC_10_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i25_LC_10_24_6 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \c0.data_out_0___i25_LC_10_24_6  (
            .in0(N__37716),
            .in1(N__23831),
            .in2(N__33504),
            .in3(N__28758),
            .lcout(data_out_19_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37578),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_906_LC_10_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_906_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_906_LC_10_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_906_LC_10_24_7  (
            .in0(N__27987),
            .in1(N__24782),
            .in2(_gnd_net_),
            .in3(N__23684),
            .lcout(\c0.n5533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_931_LC_10_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_931_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_931_LC_10_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_931_LC_10_25_0  (
            .in0(N__35040),
            .in1(N__34970),
            .in2(_gnd_net_),
            .in3(N__34707),
            .lcout(n4_adj_1975),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i17_3_lut_LC_10_25_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i17_3_lut_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i17_3_lut_LC_10_25_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i17_3_lut_LC_10_25_1  (
            .in0(N__34326),
            .in1(N__28548),
            .in2(_gnd_net_),
            .in3(N__23633),
            .lcout(),
            .ltout(\c0.n17_adj_1913_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5575_3_lut_LC_10_25_2 .C_ON=1'b0;
    defparam \c0.i5575_3_lut_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5575_3_lut_LC_10_25_2 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \c0.i5575_3_lut_LC_10_25_2  (
            .in0(N__33781),
            .in1(_gnd_net_),
            .in2(N__23751),
            .in3(N__34072),
            .lcout(\c0.n5830 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_894_LC_10_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_894_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_894_LC_10_25_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_894_LC_10_25_3  (
            .in0(N__33665),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35038),
            .lcout(n4_adj_1982),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i957_4_lut_LC_10_25_4 .C_ON=1'b0;
    defparam \c0.i957_4_lut_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i957_4_lut_LC_10_25_4 .LUT_INIT=16'b1001000111000100;
    LogicCell40 \c0.i957_4_lut_LC_10_25_4  (
            .in0(N__34211),
            .in1(N__34070),
            .in2(N__28770),
            .in3(N__34325),
            .lcout(\c0.n1198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_10_25_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_10_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_10_25_5 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_10_25_5  (
            .in0(N__29282),
            .in1(N__23748),
            .in2(N__33612),
            .in3(N__23808),
            .lcout(\c0.tx.r_Tx_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37584),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_904_LC_10_25_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_904_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_904_LC_10_25_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_904_LC_10_25_6  (
            .in0(N__35039),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34971),
            .lcout(n1991),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5563_3_lut_LC_10_25_7 .C_ON=1'b0;
    defparam \c0.i5563_3_lut_LC_10_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5563_3_lut_LC_10_25_7 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \c0.i5563_3_lut_LC_10_25_7  (
            .in0(N__34071),
            .in1(N__33780),
            .in2(_gnd_net_),
            .in3(N__26235),
            .lcout(\c0.n5827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i746_2_lut_LC_10_26_0 .C_ON=1'b0;
    defparam \c0.i746_2_lut_LC_10_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i746_2_lut_LC_10_26_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i746_2_lut_LC_10_26_0  (
            .in0(_gnd_net_),
            .in1(N__34132),
            .in2(_gnd_net_),
            .in3(N__34079),
            .lcout(\c0.n1253 ),
            .ltout(\c0.n1253_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_10_26_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_10_26_1 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i31_4_lut_LC_10_26_1  (
            .in0(N__33633),
            .in1(N__26169),
            .in2(N__23742),
            .in3(N__33738),
            .lcout(tx_data_2_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_841_LC_10_26_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_841_LC_10_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_841_LC_10_26_3 .LUT_INIT=16'b0011111100100010;
    LogicCell40 \c0.i1_4_lut_adj_841_LC_10_26_3  (
            .in0(N__34328),
            .in1(N__34212),
            .in2(N__33396),
            .in3(N__34080),
            .lcout(),
            .ltout(\c0.n22_adj_1914_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_10_26_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_10_26_4 .LUT_INIT=16'b1101110110001101;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i31_4_lut_LC_10_26_4  (
            .in0(N__33739),
            .in1(N__23739),
            .in2(N__23730),
            .in3(N__34134),
            .lcout(tx_data_6_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_10_26_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_10_26_5 .LUT_INIT=16'b1100110010101111;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i31_4_lut_LC_10_26_5  (
            .in0(N__26295),
            .in1(N__23877),
            .in2(N__23871),
            .in3(N__33740),
            .lcout(tx_data_7_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5588_4_lut_LC_10_26_6 .C_ON=1'b0;
    defparam \c0.i5588_4_lut_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5588_4_lut_LC_10_26_6 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \c0.i5588_4_lut_LC_10_26_6  (
            .in0(N__23846),
            .in1(N__26200),
            .in2(N__23835),
            .in3(N__34327),
            .lcout(),
            .ltout(\c0.n5810_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_10_26_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_10_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_10_26_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i31_4_lut_LC_10_26_7  (
            .in0(N__34133),
            .in1(N__23817),
            .in2(N__23811),
            .in3(N__33737),
            .lcout(\c0.tx_data_0_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5281_4_lut_LC_10_27_0 .C_ON=1'b0;
    defparam \c0.tx.i5281_4_lut_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5281_4_lut_LC_10_27_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i5281_4_lut_LC_10_27_0  (
            .in0(N__24096),
            .in1(N__23929),
            .in2(N__24069),
            .in3(N__23778),
            .lcout(\c0.tx.n5627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i6_4_lut_LC_10_27_1 .C_ON=1'b0;
    defparam \c0.tx.i6_4_lut_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i6_4_lut_LC_10_27_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i6_4_lut_LC_10_27_1  (
            .in0(N__24066),
            .in1(N__24097),
            .in2(N__23984),
            .in3(N__24033),
            .lcout(),
            .ltout(\c0.tx.n14_adj_1869_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i7_4_lut_LC_10_27_2 .C_ON=1'b0;
    defparam \c0.tx.i7_4_lut_LC_10_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i7_4_lut_LC_10_27_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i7_4_lut_LC_10_27_2  (
            .in0(N__24045),
            .in1(N__26280),
            .in2(N__23796),
            .in3(N__23779),
            .lcout(\c0.tx.r_SM_Main_2_N_1767_1 ),
            .ltout(\c0.tx.r_SM_Main_2_N_1767_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_10_27_3 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_10_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_10_27_3 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_10_27_3  (
            .in0(N__28976),
            .in1(N__29174),
            .in2(N__23793),
            .in3(N__29090),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37598),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i5_LC_10_27_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i5_LC_10_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_10_27_4 .LUT_INIT=16'b1100110000001010;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_10_27_4  (
            .in0(N__23790),
            .in1(N__23780),
            .in2(N__23985),
            .in3(N__28978),
            .lcout(\c0.tx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37598),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i6_LC_10_27_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i6_LC_10_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_10_27_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_10_27_5  (
            .in0(N__28975),
            .in1(N__26458),
            .in2(N__23763),
            .in3(N__24098),
            .lcout(r_Clock_Count_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37598),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i4_LC_10_27_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i4_LC_10_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_10_27_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_10_27_6  (
            .in0(N__26457),
            .in1(N__28977),
            .in2(N__24081),
            .in3(N__24067),
            .lcout(r_Clock_Count_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37598),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_LC_10_27_7 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_LC_10_27_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.tx.i2_2_lut_LC_10_27_7  (
            .in0(N__23928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26533),
            .lcout(\c0.tx.n10_adj_1868 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5283_3_lut_4_lut_LC_10_28_0 .C_ON=1'b0;
    defparam \c0.tx.i5283_3_lut_4_lut_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5283_3_lut_4_lut_LC_10_28_0 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \c0.tx.i5283_3_lut_4_lut_LC_10_28_0  (
            .in0(N__26532),
            .in1(N__26493),
            .in2(N__24039),
            .in3(N__26412),
            .lcout(\c0.tx.n5629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_10_28_2.C_ON=1'b0;
    defparam i1_2_lut_LC_10_28_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_10_28_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_LC_10_28_2 (
            .in0(_gnd_net_),
            .in1(N__29198),
            .in2(_gnd_net_),
            .in3(N__29070),
            .lcout(n11_adj_1979),
            .ltout(n11_adj_1979_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_adj_805_LC_10_28_3 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_adj_805_LC_10_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_adj_805_LC_10_28_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx.i2_4_lut_adj_805_LC_10_28_3  (
            .in0(N__28956),
            .in1(N__24012),
            .in2(N__24006),
            .in3(N__24003),
            .lcout(\c0.tx.n3120 ),
            .ltout(\c0.tx.n3120_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_3_lut_LC_10_28_4 .C_ON=1'b0;
    defparam \c0.tx.i1_3_lut_LC_10_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_3_lut_LC_10_28_4 .LUT_INIT=16'b0000000010101111;
    LogicCell40 \c0.tx.i1_3_lut_LC_10_28_4  (
            .in0(N__23980),
            .in1(_gnd_net_),
            .in2(N__23946),
            .in3(N__28957),
            .lcout(n782),
            .ltout(n782_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i8_LC_10_28_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_10_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_10_28_5 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_10_28_5  (
            .in0(N__28958),
            .in1(N__23943),
            .in2(N__23934),
            .in3(N__23931),
            .lcout(r_Clock_Count_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37604),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i75_LC_11_15_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i75_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i75_LC_11_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i75_LC_11_15_3  (
            .in0(N__35631),
            .in1(N__23890),
            .in2(_gnd_net_),
            .in3(N__30671),
            .lcout(data_in_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37541),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_819_LC_11_17_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_819_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_819_LC_11_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_819_LC_11_17_0  (
            .in0(N__24453),
            .in1(N__24447),
            .in2(N__24426),
            .in3(N__24411),
            .lcout(\c0.n24_adj_1885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_11_17_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_11_17_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_LC_11_17_1  (
            .in0(N__25555),
            .in1(N__26739),
            .in2(N__25901),
            .in3(N__24384),
            .lcout(),
            .ltout(\c0.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_822_LC_11_17_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_822_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_822_LC_11_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_822_LC_11_17_2  (
            .in0(N__24366),
            .in1(N__24324),
            .in2(N__24273),
            .in3(N__24270),
            .lcout(\c0.n5519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i17_LC_11_17_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i17_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i17_LC_11_17_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i17_LC_11_17_3  (
            .in0(N__28419),
            .in1(N__35685),
            .in2(_gnd_net_),
            .in3(N__27861),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37517),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i55_LC_11_17_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i55_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i55_LC_11_17_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i55_LC_11_17_5  (
            .in0(N__24202),
            .in1(N__35686),
            .in2(_gnd_net_),
            .in3(N__24239),
            .lcout(data_in_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37517),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i45_LC_11_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i45_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i45_LC_11_18_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i45_LC_11_18_0  (
            .in0(N__32128),
            .in1(N__24890),
            .in2(N__27363),
            .in3(N__33103),
            .lcout(\c0.data_in_field_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37531),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i137_LC_11_18_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i137_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i137_LC_11_18_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i137_LC_11_18_2  (
            .in0(N__30694),
            .in1(_gnd_net_),
            .in2(N__36063),
            .in3(N__24169),
            .lcout(data_in_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37531),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i101_LC_11_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i101_LC_11_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i101_LC_11_18_3 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i101_LC_11_18_3  (
            .in0(N__24845),
            .in1(N__33102),
            .in2(N__24990),
            .in3(N__32129),
            .lcout(\c0.data_in_field_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37531),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_998_LC_11_18_4 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_998_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_998_LC_11_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_998_LC_11_18_4  (
            .in0(N__24144),
            .in1(N__24134),
            .in2(N__24120),
            .in3(N__24914),
            .lcout(\c0.n35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_856_LC_11_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_856_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_856_LC_11_18_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_856_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__24886),
            .in2(_gnd_net_),
            .in3(N__24832),
            .lcout(\c0.n4_adj_1920 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_996_LC_11_18_6 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_996_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_996_LC_11_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_996_LC_11_18_6  (
            .in0(N__24802),
            .in1(N__24750),
            .in2(N__24732),
            .in3(N__24714),
            .lcout(),
            .ltout(\c0.n31_adj_1900_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_833_LC_11_18_7 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_833_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_833_LC_11_18_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i19_4_lut_adj_833_LC_11_18_7  (
            .in0(N__26586),
            .in1(N__25068),
            .in2(N__24693),
            .in3(N__24690),
            .lcout(\c0.n5582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i3_LC_11_19_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i3_LC_11_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i3_LC_11_19_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0___i3_LC_11_19_0  (
            .in0(N__33104),
            .in1(N__27241),
            .in2(N__24684),
            .in3(N__32131),
            .lcout(\c0.data_in_field_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37542),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_838_LC_11_19_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_838_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_838_LC_11_19_3 .LUT_INIT=16'b1111111111101101;
    LogicCell40 \c0.i9_4_lut_adj_838_LC_11_19_3  (
            .in0(N__24651),
            .in1(N__24645),
            .in2(N__24639),
            .in3(N__24627),
            .lcout(\c0.n25_adj_1907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_858_LC_11_19_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_858_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_858_LC_11_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_858_LC_11_19_4  (
            .in0(N__30243),
            .in1(N__24612),
            .in2(N__27242),
            .in3(N__24604),
            .lcout(\c0.n5593 ),
            .ltout(\c0.n5593_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_974_LC_11_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_974_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_974_LC_11_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_974_LC_11_19_5  (
            .in0(N__24527),
            .in1(N__26897),
            .in2(N__24480),
            .in3(N__26960),
            .lcout(\c0.n5430 ),
            .ltout(\c0.n5430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_999_LC_11_19_6 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_999_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_999_LC_11_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i17_4_lut_adj_999_LC_11_19_6  (
            .in0(N__27032),
            .in1(N__24471),
            .in2(N__24465),
            .in3(N__24462),
            .lcout(\c0.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i14_LC_11_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i14_LC_11_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i14_LC_11_20_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0___i14_LC_11_20_0  (
            .in0(N__33106),
            .in1(N__25062),
            .in2(N__25026),
            .in3(N__32127),
            .lcout(\c0.data_in_field_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_LC_11_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_LC_11_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_LC_11_20_1  (
            .in0(N__25789),
            .in1(N__30569),
            .in2(N__30935),
            .in3(N__30534),
            .lcout(\c0.n6_adj_1939 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i101_LC_11_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i101_LC_11_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i101_LC_11_20_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_in_0___i101_LC_11_20_2  (
            .in0(N__24982),
            .in1(_gnd_net_),
            .in2(N__30291),
            .in3(N__35906),
            .lcout(data_in_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i89_LC_11_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i89_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i89_LC_11_20_3 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i89_LC_11_20_3  (
            .in0(N__28339),
            .in1(N__32130),
            .in2(N__30483),
            .in3(N__33105),
            .lcout(\c0.data_in_field_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i65_LC_11_20_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i65_LC_11_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i65_LC_11_20_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i65_LC_11_20_4  (
            .in0(N__25869),
            .in1(N__35907),
            .in2(_gnd_net_),
            .in3(N__31045),
            .lcout(data_in_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i93_LC_11_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i93_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i93_LC_11_20_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i93_LC_11_20_5  (
            .in0(N__35905),
            .in1(N__24958),
            .in2(_gnd_net_),
            .in3(N__24983),
            .lcout(data_in_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37551),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_942_LC_11_20_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_942_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_942_LC_11_20_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_942_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(N__30926),
            .in2(_gnd_net_),
            .in3(N__25788),
            .lcout(\c0.n2089 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_868_LC_11_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_868_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_868_LC_11_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_868_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__27443),
            .in2(_gnd_net_),
            .in3(N__24927),
            .lcout(\c0.n5581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i88_LC_11_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i88_LC_11_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i88_LC_11_21_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i88_LC_11_21_1  (
            .in0(N__32992),
            .in1(N__32164),
            .in2(N__28121),
            .in3(N__31367),
            .lcout(\c0.data_in_field_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37561),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i73_LC_11_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i73_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i73_LC_11_21_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i73_LC_11_21_2  (
            .in0(N__32161),
            .in1(N__32994),
            .in2(N__25868),
            .in3(N__25793),
            .lcout(\c0.data_in_field_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37561),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i129_LC_11_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i129_LC_11_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i129_LC_11_21_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i129_LC_11_21_3  (
            .in0(N__32991),
            .in1(N__32163),
            .in2(N__35103),
            .in3(N__28045),
            .lcout(\c0.data_in_field_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37561),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i121_LC_11_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i121_LC_11_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i121_LC_11_21_5 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i121_LC_11_21_5  (
            .in0(N__32990),
            .in1(N__32162),
            .in2(N__35073),
            .in3(N__25543),
            .lcout(\c0.data_in_field_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37561),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i43_LC_11_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i43_LC_11_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i43_LC_11_21_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i43_LC_11_21_6  (
            .in0(N__32160),
            .in1(N__32993),
            .in2(N__25629),
            .in3(N__25828),
            .lcout(\c0.data_in_field_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37561),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_969_LC_11_21_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_969_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_969_LC_11_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_969_LC_11_21_7  (
            .in0(N__28277),
            .in1(N__25542),
            .in2(_gnd_net_),
            .in3(N__28044),
            .lcout(\c0.n2107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i155_LC_11_22_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i155_LC_11_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i155_LC_11_22_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i155_LC_11_22_0  (
            .in0(N__25894),
            .in1(N__25500),
            .in2(_gnd_net_),
            .in3(N__35918),
            .lcout(data_in_19_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37571),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6201_bdd_4_lut_LC_11_22_1 .C_ON=1'b0;
    defparam \c0.n6201_bdd_4_lut_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.n6201_bdd_4_lut_LC_11_22_1 .LUT_INIT=16'b1010110110101000;
    LogicCell40 \c0.n6201_bdd_4_lut_LC_11_22_1  (
            .in0(N__25479),
            .in1(N__26646),
            .in2(N__30206),
            .in3(N__25462),
            .lcout(),
            .ltout(\c0.n5716_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5844_LC_11_22_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5844_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_5844_LC_11_22_2 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_5844_LC_11_22_2  (
            .in0(N__25409),
            .in1(N__25259),
            .in2(N__25161),
            .in3(N__25914),
            .lcout(\c0.n6195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5829_LC_11_22_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5829_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5829_LC_11_22_3 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5829_LC_11_22_3  (
            .in0(N__27743),
            .in1(N__25152),
            .in2(N__30205),
            .in3(N__25113),
            .lcout(),
            .ltout(\c0.n6207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6207_bdd_4_lut_LC_11_22_4 .C_ON=1'b0;
    defparam \c0.n6207_bdd_4_lut_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.n6207_bdd_4_lut_LC_11_22_4 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n6207_bdd_4_lut_LC_11_22_4  (
            .in0(N__25994),
            .in1(N__30180),
            .in2(N__25950),
            .in3(N__25946),
            .lcout(\c0.n5713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i147_LC_11_22_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i147_LC_11_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i147_LC_11_22_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_in_0___i147_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__25893),
            .in2(N__36022),
            .in3(N__25714),
            .lcout(data_in_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37571),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i73_LC_11_22_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i73_LC_11_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i73_LC_11_22_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i73_LC_11_22_6  (
            .in0(N__30453),
            .in1(N__25861),
            .in2(_gnd_net_),
            .in3(N__35919),
            .lcout(data_in_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37571),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_875_LC_11_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_875_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_875_LC_11_22_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_875_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__25821),
            .in2(_gnd_net_),
            .in3(N__25787),
            .lcout(\c0.n2068 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i89_LC_11_23_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i89_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i89_LC_11_23_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i89_LC_11_23_0  (
            .in0(N__35821),
            .in1(N__25764),
            .in2(_gnd_net_),
            .in3(N__30469),
            .lcout(data_in_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37579),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i139_LC_11_23_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i139_LC_11_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i139_LC_11_23_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i139_LC_11_23_1  (
            .in0(N__25715),
            .in1(N__25673),
            .in2(_gnd_net_),
            .in3(N__35822),
            .lcout(data_in_17_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37579),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i43_LC_11_23_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i43_LC_11_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i43_LC_11_23_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i43_LC_11_23_2  (
            .in0(N__25661),
            .in1(N__35823),
            .in2(_gnd_net_),
            .in3(N__25615),
            .lcout(data_in_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37579),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i30_LC_11_23_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i30_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i30_LC_11_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i30_LC_11_23_4  (
            .in0(N__35820),
            .in1(N__25595),
            .in2(_gnd_net_),
            .in3(N__27889),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37579),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i88_LC_11_23_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i88_LC_11_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i88_LC_11_23_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i88_LC_11_23_5  (
            .in0(N__35824),
            .in1(N__26162),
            .in2(_gnd_net_),
            .in3(N__31357),
            .lcout(data_in_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37579),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i6_LC_11_23_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i6_LC_11_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i6_LC_11_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter__i6_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(N__33457),
            .in2(_gnd_net_),
            .in3(N__33336),
            .lcout(\c0.byte_transmit_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37579),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_11_24_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i17_3_lut_LC_11_24_1  (
            .in0(N__26123),
            .in1(N__26111),
            .in2(_gnd_net_),
            .in3(N__34332),
            .lcout(\c0.n17_adj_1908 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_968_LC_11_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_968_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_968_LC_11_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_968_LC_11_24_2  (
            .in0(N__36518),
            .in1(N__34657),
            .in2(_gnd_net_),
            .in3(N__35013),
            .lcout(),
            .ltout(n5448_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i29_LC_11_24_3 .C_ON=1'b0;
    defparam \c0.data_out_0___i29_LC_11_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i29_LC_11_24_3 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \c0.data_out_0___i29_LC_11_24_3  (
            .in0(N__37708),
            .in1(N__26124),
            .in2(N__26136),
            .in3(N__26133),
            .lcout(data_out_19_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37585),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i21_LC_11_24_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i21_LC_11_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i21_LC_11_24_4 .LUT_INIT=16'b1011100010001011;
    LogicCell40 \c0.data_out_0___i21_LC_11_24_4  (
            .in0(N__26112),
            .in1(N__37707),
            .in2(N__33516),
            .in3(N__28692),
            .lcout(data_out_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37585),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_859_LC_11_24_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_859_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_859_LC_11_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i9_4_lut_adj_859_LC_11_24_5  (
            .in0(N__26103),
            .in1(N__26085),
            .in2(N__26067),
            .in3(N__26049),
            .lcout(),
            .ltout(\c0.n20_adj_1922_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_862_LC_11_24_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_862_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_862_LC_11_24_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_862_LC_11_24_6  (
            .in0(N__26043),
            .in1(N__26025),
            .in2(N__26007),
            .in3(N__26004),
            .lcout(n21_adj_1977),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5571_4_lut_LC_11_25_0 .C_ON=1'b0;
    defparam \c0.i5571_4_lut_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5571_4_lut_LC_11_25_0 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \c0.i5571_4_lut_LC_11_25_0  (
            .in0(N__34324),
            .in1(N__26475),
            .in2(N__28533),
            .in3(N__26201),
            .lcout(\c0.n5833 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_865_LC_11_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_865_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_865_LC_11_25_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.i1_2_lut_adj_865_LC_11_25_1  (
            .in0(_gnd_net_),
            .in1(N__36731),
            .in2(_gnd_net_),
            .in3(N__36825),
            .lcout(n4334),
            .ltout(n4334_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i28_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.data_out_0___i28_LC_11_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i28_LC_11_25_2 .LUT_INIT=16'b1100101011000101;
    LogicCell40 \c0.data_out_0___i28_LC_11_25_2  (
            .in0(N__28517),
            .in1(N__33926),
            .in2(N__26256),
            .in3(N__26253),
            .lcout(data_out_19_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37593),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_11_25_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_11_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_11_25_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i17_3_lut_LC_11_25_3  (
            .in0(N__26246),
            .in1(N__26213),
            .in2(_gnd_net_),
            .in3(N__34323),
            .lcout(\c0.n17_adj_1950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i27_LC_11_25_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i27_LC_11_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i27_LC_11_25_4 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \c0.data_out_0___i27_LC_11_25_4  (
            .in0(N__26186),
            .in1(N__26229),
            .in2(N__28518),
            .in3(N__37702),
            .lcout(data_out_19_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37593),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_11_25_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_11_25_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i31_4_lut_LC_11_25_5  (
            .in0(N__26202),
            .in1(N__33678),
            .in2(N__26223),
            .in3(N__33722),
            .lcout(tx_data_4_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i24_LC_11_25_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i24_LC_11_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i24_LC_11_25_7 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_out_0___i24_LC_11_25_7  (
            .in0(N__26214),
            .in1(N__36732),
            .in2(N__28674),
            .in3(N__36826),
            .lcout(data_out_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37593),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_997_LC_11_26_0 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_997_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_997_LC_11_26_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_997_LC_11_26_0  (
            .in0(N__34204),
            .in1(N__34130),
            .in2(_gnd_net_),
            .in3(N__34067),
            .lcout(\c0.n1508 ),
            .ltout(\c0.n1508_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5587_4_lut_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.i5587_4_lut_LC_11_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5587_4_lut_LC_11_26_1 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \c0.i5587_4_lut_LC_11_26_1  (
            .in0(N__26187),
            .in1(N__26303),
            .in2(N__26172),
            .in3(N__34331),
            .lcout(\c0.n5840 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_11_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_11_26_2 .LUT_INIT=16'b0110010011101100;
    LogicCell40 \c0.byte_transmit_counter_2__bdd_4_lut_4_lut_LC_11_26_2  (
            .in0(N__34206),
            .in1(N__34131),
            .in2(N__28650),
            .in3(N__34068),
            .lcout(),
            .ltout(\c0.n6309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6309_bdd_4_lut_4_lut_LC_11_26_3 .C_ON=1'b0;
    defparam \c0.n6309_bdd_4_lut_4_lut_LC_11_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.n6309_bdd_4_lut_4_lut_LC_11_26_3 .LUT_INIT=16'b1110000111100011;
    LogicCell40 \c0.n6309_bdd_4_lut_4_lut_LC_11_26_3  (
            .in0(N__34069),
            .in1(N__34207),
            .in2(N__26307),
            .in3(N__34330),
            .lcout(\c0.n6312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i19_LC_11_26_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i19_LC_11_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i19_LC_11_26_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.data_out_0___i19_LC_11_26_4  (
            .in0(N__26304),
            .in1(N__37706),
            .in2(N__36591),
            .in3(N__36440),
            .lcout(data_out_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37599),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1006_4_lut_LC_11_26_5 .C_ON=1'b0;
    defparam \c0.i1006_4_lut_LC_11_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1006_4_lut_LC_11_26_5 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \c0.i1006_4_lut_LC_11_26_5  (
            .in0(N__34531),
            .in1(N__34205),
            .in2(N__36519),
            .in3(N__34329),
            .lcout(\c0.n1249 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_11_26_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_11_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_11_26_6 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_11_26_6  (
            .in0(N__28452),
            .in1(N__29091),
            .in2(_gnd_net_),
            .in3(N__29321),
            .lcout(\c0.tx.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37599),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_857_LC_11_26_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_857_LC_11_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_857_LC_11_26_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_857_LC_11_26_7  (
            .in0(N__36176),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34658),
            .lcout(n1768),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_11_27_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_11_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_11_27_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_11_27_0  (
            .in0(N__33598),
            .in1(N__33833),
            .in2(_gnd_net_),
            .in3(N__26289),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37605),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i3401_2_lut_LC_11_27_1 .C_ON=1'b0;
    defparam \c0.tx.i3401_2_lut_LC_11_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i3401_2_lut_LC_11_27_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx.i3401_2_lut_LC_11_27_1  (
            .in0(_gnd_net_),
            .in1(N__26494),
            .in2(_gnd_net_),
            .in3(N__26413),
            .lcout(\c0.tx.n3644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5566_2_lut_3_lut_LC_11_27_2 .C_ON=1'b0;
    defparam \c0.tx.i5566_2_lut_3_lut_LC_11_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5566_2_lut_3_lut_LC_11_27_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i5566_2_lut_3_lut_LC_11_27_2  (
            .in0(N__29204),
            .in1(N__29087),
            .in2(_gnd_net_),
            .in3(N__28485),
            .lcout(),
            .ltout(n5818_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Done_44_LC_11_27_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Done_44_LC_11_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Done_44_LC_11_27_3 .LUT_INIT=16'b1011101111111000;
    LogicCell40 \c0.tx.r_Tx_Done_44_LC_11_27_3  (
            .in0(N__26265),
            .in1(N__26274),
            .in2(N__26268),
            .in3(N__28973),
            .lcout(n4155),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37605),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i3_LC_11_27_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i3_LC_11_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_11_27_4 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_11_27_4  (
            .in0(N__28968),
            .in1(N__26460),
            .in2(N__26550),
            .in3(N__26537),
            .lcout(r_Clock_Count_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37605),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_11_27_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i0_LC_11_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_11_27_5 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_11_27_5  (
            .in0(N__26459),
            .in1(N__28969),
            .in2(N__26511),
            .in3(N__26495),
            .lcout(r_Clock_Count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37605),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_11_27_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_11_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_11_27_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_11_27_6  (
            .in0(N__29205),
            .in1(N__29088),
            .in2(N__29004),
            .in3(N__28486),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37605),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i22_LC_11_27_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i22_LC_11_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i22_LC_11_27_7 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \c0.data_out_0___i22_LC_11_27_7  (
            .in0(N__33624),
            .in1(N__26474),
            .in2(N__37757),
            .in3(N__37726),
            .lcout(data_out_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37605),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i1_LC_11_28_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i1_LC_11_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_11_28_1 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_11_28_1  (
            .in0(N__28974),
            .in1(N__26456),
            .in2(N__26436),
            .in3(N__26417),
            .lcout(r_Clock_Count_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37609),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i154_LC_11_29_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i154_LC_11_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i154_LC_11_29_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i154_LC_11_29_7  (
            .in0(N__35760),
            .in1(N__26391),
            .in2(_gnd_net_),
            .in3(N__26700),
            .lcout(data_in_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37614),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i108_LC_12_17_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i108_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i108_LC_12_17_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i108_LC_12_17_1  (
            .in0(N__35693),
            .in1(N__26366),
            .in2(_gnd_net_),
            .in3(N__26321),
            .lcout(data_in_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37528),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i129_LC_12_17_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i129_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i129_LC_12_17_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i129_LC_12_17_6  (
            .in0(N__35719),
            .in1(N__30695),
            .in2(_gnd_net_),
            .in3(N__35086),
            .lcout(data_in_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37528),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i86_LC_12_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i86_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i86_LC_12_18_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i86_LC_12_18_1  (
            .in0(N__36020),
            .in1(N__27014),
            .in2(_gnd_net_),
            .in3(N__28840),
            .lcout(data_in_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37543),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i109_LC_12_18_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i109_LC_12_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i109_LC_12_18_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i109_LC_12_18_2  (
            .in0(N__26918),
            .in1(N__36021),
            .in2(_gnd_net_),
            .in3(N__30280),
            .lcout(data_in_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37543),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5661_LC_12_18_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5661_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5661_LC_12_18_4 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5661_LC_12_18_4  (
            .in0(N__26991),
            .in1(N__27754),
            .in2(N__30209),
            .in3(N__26964),
            .lcout(\c0.n5997 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i117_LC_12_18_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i117_LC_12_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i117_LC_12_18_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i117_LC_12_18_5  (
            .in0(N__36019),
            .in1(N__26917),
            .in2(_gnd_net_),
            .in3(N__30308),
            .lcout(data_in_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37543),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5685_LC_12_18_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5685_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5685_LC_12_18_6 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5685_LC_12_18_6  (
            .in0(N__30198),
            .in1(N__27755),
            .in2(N__26904),
            .in3(N__29460),
            .lcout(),
            .ltout(\c0.n6033_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n6033_bdd_4_lut_LC_12_18_7 .C_ON=1'b0;
    defparam \c0.n6033_bdd_4_lut_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.n6033_bdd_4_lut_LC_12_18_7 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n6033_bdd_4_lut_LC_12_18_7  (
            .in0(N__26858),
            .in1(N__26805),
            .in2(N__26754),
            .in3(N__30199),
            .lcout(\c0.n5791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_889_LC_12_19_1 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_889_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_889_LC_12_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_889_LC_12_19_1  (
            .in0(N__27909),
            .in1(N__29361),
            .in2(N__28143),
            .in3(N__30903),
            .lcout(\c0.n1814 ),
            .ltout(\c0.n1814_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_993_LC_12_19_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_993_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_993_LC_12_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_993_LC_12_19_2  (
            .in0(N__26710),
            .in1(N__26676),
            .in2(N__26649),
            .in3(N__26644),
            .lcout(\c0.n32_adj_1901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i85_LC_12_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i85_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i85_LC_12_19_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i85_LC_12_19_3  (
            .in0(N__33070),
            .in1(N__32230),
            .in2(N__30423),
            .in3(N__29542),
            .lcout(\c0.data_in_field_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37552),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i70_LC_12_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i70_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i70_LC_12_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i70_LC_12_19_4  (
            .in0(N__35878),
            .in1(N__28817),
            .in2(_gnd_net_),
            .in3(N__26579),
            .lcout(data_in_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37552),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i133_LC_12_19_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i133_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i133_LC_12_19_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i133_LC_12_19_5  (
            .in0(N__35499),
            .in1(N__27399),
            .in2(_gnd_net_),
            .in3(N__30340),
            .lcout(data_in_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37552),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i37_LC_12_19_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i37_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i37_LC_12_19_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i37_LC_12_19_6  (
            .in0(N__35877),
            .in1(N__31210),
            .in2(_gnd_net_),
            .in3(N__27356),
            .lcout(data_in_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37552),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i25_LC_12_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i25_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i25_LC_12_19_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \c0.data_in_frame_0___i25_LC_12_19_7  (
            .in0(N__27856),
            .in1(N__32229),
            .in2(N__33218),
            .in3(N__27442),
            .lcout(\c0.data_in_field_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37552),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_913_LC_12_20_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_913_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_913_LC_12_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_913_LC_12_20_0  (
            .in0(N__27435),
            .in1(N__30593),
            .in2(N__31407),
            .in3(N__30561),
            .lcout(\c0.n5560 ),
            .ltout(\c0.n5560_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_LC_12_20_1 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_LC_12_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_LC_12_20_1  (
            .in0(N__27300),
            .in1(N__27234),
            .in2(N__27213),
            .in3(N__30230),
            .lcout(\c0.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i40_LC_12_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i40_LC_12_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i40_LC_12_20_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i40_LC_12_20_2  (
            .in0(N__35923),
            .in1(N__31432),
            .in2(_gnd_net_),
            .in3(N__27188),
            .lcout(data_in_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37562),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_947_LC_12_20_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_947_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_947_LC_12_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_947_LC_12_20_3  (
            .in0(N__27164),
            .in1(N__27138),
            .in2(N__30606),
            .in3(N__27099),
            .lcout(\c0.n5378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i94_LC_12_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i94_LC_12_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i94_LC_12_20_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i94_LC_12_20_5  (
            .in0(N__35925),
            .in1(N__27007),
            .in2(_gnd_net_),
            .in3(N__34457),
            .lcout(data_in_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37562),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i99_LC_12_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i99_LC_12_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i99_LC_12_21_0 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0___i99_LC_12_21_0  (
            .in0(N__33234),
            .in1(N__28281),
            .in2(N__32241),
            .in3(N__31277),
            .lcout(\c0.data_in_field_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37572),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i17_LC_12_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i17_LC_12_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i17_LC_12_21_2 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0___i17_LC_12_21_2  (
            .in0(N__32165),
            .in1(N__28433),
            .in2(N__33272),
            .in3(N__30934),
            .lcout(\c0.data_in_field_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37572),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i99_LC_12_21_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i99_LC_12_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i99_LC_12_21_3 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \c0.data_in_0___i99_LC_12_21_3  (
            .in0(N__35924),
            .in1(N__28391),
            .in2(N__31281),
            .in3(_gnd_net_),
            .lcout(data_in_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37572),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_3_lut_4_lut_adj_1001_LC_12_21_5 .C_ON=1'b0;
    defparam \c0.i8_3_lut_4_lut_adj_1001_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_3_lut_4_lut_adj_1001_LC_12_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_3_lut_4_lut_adj_1001_LC_12_21_5  (
            .in0(N__28332),
            .in1(N__28270),
            .in2(N__28234),
            .in3(N__28197),
            .lcout(\c0.n23_adj_1935 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_878_LC_12_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_878_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_878_LC_12_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_878_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__28096),
            .in2(_gnd_net_),
            .in3(N__28043),
            .lcout(),
            .ltout(\c0.n1965_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_887_LC_12_21_7 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_887_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_887_LC_12_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_887_LC_12_21_7  (
            .in0(N__28016),
            .in1(N__28001),
            .in2(N__27960),
            .in3(N__27953),
            .lcout(\c0.n24_adj_1930 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_876_LC_12_22_3 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_876_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_876_LC_12_22_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i12_4_lut_adj_876_LC_12_22_3  (
            .in0(N__27882),
            .in1(N__27857),
            .in2(N__31130),
            .in3(N__27814),
            .lcout(\c0.n28_adj_1925 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5704_LC_12_22_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5704_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_5704_LC_12_22_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_5704_LC_12_22_6  (
            .in0(N__27744),
            .in1(N__27444),
            .in2(N__30194),
            .in3(N__30933),
            .lcout(\c0.n6039 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i16_3_lut_4_lut_4_lut_LC_12_23_0 .C_ON=1'b0;
    defparam \c0.tx.i16_3_lut_4_lut_4_lut_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i16_3_lut_4_lut_4_lut_LC_12_23_0 .LUT_INIT=16'b1001100000010000;
    LogicCell40 \c0.tx.i16_3_lut_4_lut_4_lut_LC_12_23_0  (
            .in0(N__29202),
            .in1(N__29113),
            .in2(N__28608),
            .in3(N__28497),
            .lcout(),
            .ltout(n5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_12_23_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_12_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_12_23_1 .LUT_INIT=16'b1000101010111010;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_12_23_1  (
            .in0(N__28637),
            .in1(N__29015),
            .in2(N__28506),
            .in3(N__29114),
            .lcout(tx_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_809_LC_12_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_809_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_809_LC_12_23_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i1_2_lut_adj_809_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__28503),
            .in2(_gnd_net_),
            .in3(N__28636),
            .lcout(\c0.n50_adj_1875 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_prev_1793_LC_12_23_3 .C_ON=1'b0;
    defparam \c0.tx_active_prev_1793_LC_12_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx_active_prev_1793_LC_12_23_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.tx_active_prev_1793_LC_12_23_3  (
            .in0(N__28638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.tx_active_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_4_lut_adj_804_LC_12_23_4 .C_ON=1'b0;
    defparam \c0.tx.i2_4_lut_adj_804_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_4_lut_adj_804_LC_12_23_4 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \c0.tx.i2_4_lut_adj_804_LC_12_23_4  (
            .in0(N__29201),
            .in1(N__29112),
            .in2(N__29021),
            .in3(N__28496),
            .lcout(\c0.tx.n2177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_12_23_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_12_23_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_LC_12_23_5  (
            .in0(N__33356),
            .in1(N__33332),
            .in2(_gnd_net_),
            .in3(N__33302),
            .lcout(\c0.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i5_LC_12_23_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i5_LC_12_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i5_LC_12_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter__i5_LC_12_23_6  (
            .in0(_gnd_net_),
            .in1(N__33456),
            .in2(_gnd_net_),
            .in3(N__33357),
            .lcout(\c0.byte_transmit_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37586),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5640_3_lut_4_lut_LC_12_24_0 .C_ON=1'b0;
    defparam \c0.i5640_3_lut_4_lut_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5640_3_lut_4_lut_LC_12_24_0 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \c0.i5640_3_lut_4_lut_LC_12_24_0  (
            .in0(N__33488),
            .in1(N__28639),
            .in2(N__28597),
            .in3(N__33524),
            .lcout(n4333),
            .ltout(n4333_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i10_LC_12_24_1 .C_ON=1'b0;
    defparam \c0.data_out_0___i10_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i10_LC_12_24_1 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_out_0___i10_LC_12_24_1  (
            .in0(N__36828),
            .in1(N__36303),
            .in2(N__28443),
            .in3(N__35008),
            .lcout(data_out_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37594),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_12_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_12_24_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_12_24_2  (
            .in0(N__28583),
            .in1(N__28640),
            .in2(_gnd_net_),
            .in3(N__36827),
            .lcout(\c0.n81_adj_1872 ),
            .ltout(\c0.n81_adj_1872_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i4_LC_12_24_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i4_LC_12_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i4_LC_12_24_3 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \c0.byte_transmit_counter__i4_LC_12_24_3  (
            .in0(N__33282),
            .in1(N__33437),
            .in2(N__28440),
            .in3(N__33489),
            .lcout(\c0.byte_transmit_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37594),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_1794_LC_12_24_4 .C_ON=1'b0;
    defparam \c0.tx_transmit_1794_LC_12_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_1794_LC_12_24_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \c0.tx_transmit_1794_LC_12_24_4  (
            .in0(N__33490),
            .in1(N__28641),
            .in2(N__28598),
            .in3(N__33525),
            .lcout(\c0.tx_transmit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37594),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_975_LC_12_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_975_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_975_LC_12_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_975_LC_12_24_5  (
            .in0(N__36954),
            .in1(N__33972),
            .in2(_gnd_net_),
            .in3(N__36408),
            .lcout(n135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_873_LC_12_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_873_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_873_LC_12_24_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_873_LC_12_24_6  (
            .in0(N__35007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36681),
            .lcout(n5482),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_994_LC_12_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_994_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_994_LC_12_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_994_LC_12_24_7  (
            .in0(N__34431),
            .in1(N__36683),
            .in2(_gnd_net_),
            .in3(N__36635),
            .lcout(n5433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_813_LC_12_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_813_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_813_LC_12_25_0 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_813_LC_12_25_0  (
            .in0(N__36554),
            .in1(_gnd_net_),
            .in2(N__35018),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n4_adj_1986_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i31_LC_12_25_1 .C_ON=1'b0;
    defparam \c0.data_out_0___i31_LC_12_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i31_LC_12_25_1 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \c0.data_out_0___i31_LC_12_25_1  (
            .in0(N__37705),
            .in1(N__28746),
            .in2(N__28551),
            .in3(N__28547),
            .lcout(data_out_19_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37600),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i30_LC_12_25_2 .C_ON=1'b0;
    defparam \c0.data_out_0___i30_LC_12_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i30_LC_12_25_2 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \c0.data_out_0___i30_LC_12_25_2  (
            .in0(N__34917),
            .in1(N__37704),
            .in2(N__33798),
            .in3(N__28532),
            .lcout(data_out_19_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37600),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i18_LC_12_25_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i18_LC_12_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i18_LC_12_25_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.data_out_0___i18_LC_12_25_4  (
            .in0(N__33950),
            .in1(N__37703),
            .in2(N__34905),
            .in3(N__33971),
            .lcout(data_out_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37600),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_930_LC_12_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_930_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_930_LC_12_25_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_930_LC_12_25_5  (
            .in0(N__34659),
            .in1(N__34430),
            .in2(N__36508),
            .in3(N__35012),
            .lcout(n5440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_12_25_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_12_25_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i9_3_lut_LC_12_25_6  (
            .in0(N__34279),
            .in1(_gnd_net_),
            .in2(N__36564),
            .in3(N__34380),
            .lcout(\c0.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_LC_12_25_7 .C_ON=1'b0;
    defparam \c0.i3_3_lut_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_LC_12_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i3_3_lut_LC_12_25_7  (
            .in0(N__36495),
            .in1(N__28745),
            .in2(_gnd_net_),
            .in3(N__36687),
            .lcout(n8_adj_1987),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_963_LC_12_26_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_963_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_963_LC_12_26_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_963_LC_12_26_1  (
            .in0(N__33967),
            .in1(N__36413),
            .in2(N__36965),
            .in3(N__34381),
            .lcout(n5400),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_12_26_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_12_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_12_26_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_12_26_3  (
            .in0(N__33611),
            .in1(N__28734),
            .in2(_gnd_net_),
            .in3(N__29346),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37606),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_987_LC_12_26_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_987_LC_12_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_987_LC_12_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_987_LC_12_26_5  (
            .in0(N__36430),
            .in1(N__36412),
            .in2(N__36966),
            .in3(N__34382),
            .lcout(n5364),
            .ltout(n5364_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5552_4_lut_LC_12_26_6.C_ON=1'b0;
    defparam i5552_4_lut_LC_12_26_6.SEQ_MODE=4'b0000;
    defparam i5552_4_lut_LC_12_26_6.LUT_INIT=16'b0110100110010110;
    LogicCell40 i5552_4_lut_LC_12_26_6 (
            .in0(N__28709),
            .in1(N__28688),
            .in2(N__28677),
            .in3(N__34429),
            .lcout(n5871),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_12_26_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_12_26_7 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i31_4_lut_LC_12_26_7  (
            .in0(N__28665),
            .in1(N__33912),
            .in2(N__33782),
            .in3(N__33736),
            .lcout(tx_data_3_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_12_27_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_12_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_12_27_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_12_27_0  (
            .in0(N__29355),
            .in1(_gnd_net_),
            .in2(N__28659),
            .in3(N__33610),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37610),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5572_4_lut_LC_12_27_2 .C_ON=1'b0;
    defparam \c0.i5572_4_lut_LC_12_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5572_4_lut_LC_12_27_2 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \c0.i5572_4_lut_LC_12_27_2  (
            .in0(N__36614),
            .in1(N__34066),
            .in2(N__36414),
            .in3(N__34319),
            .lcout(\c0.n5853 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_5889_LC_12_27_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_5889_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_Bit_Index_0__bdd_4_lut_5889_LC_12_27_6 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx.r_Bit_Index_0__bdd_4_lut_5889_LC_12_27_6  (
            .in0(N__29354),
            .in1(N__29345),
            .in2(N__33894),
            .in3(N__29317),
            .lcout(),
            .ltout(\c0.tx.n6051_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n6051_bdd_4_lut_LC_12_27_7 .C_ON=1'b0;
    defparam \c0.tx.n6051_bdd_4_lut_LC_12_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n6051_bdd_4_lut_LC_12_27_7 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.tx.n6051_bdd_4_lut_LC_12_27_7  (
            .in0(N__29264),
            .in1(N__29286),
            .in2(N__29268),
            .in3(N__33892),
            .lcout(\c0.tx.n6054 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_12_28_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_12_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_12_28_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_12_28_0  (
            .in0(N__33571),
            .in1(N__29265),
            .in2(_gnd_net_),
            .in3(N__33687),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37615),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i367827_i1_3_lut_LC_12_28_4 .C_ON=1'b0;
    defparam \c0.tx.i367827_i1_3_lut_LC_12_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i367827_i1_3_lut_LC_12_28_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.i367827_i1_3_lut_LC_12_28_4  (
            .in0(N__29252),
            .in1(N__29211),
            .in2(_gnd_net_),
            .in3(N__33804),
            .lcout(),
            .ltout(\c0.tx.o_Tx_Serial_N_1798_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i26_3_lut_LC_12_28_5 .C_ON=1'b0;
    defparam \c0.tx.i26_3_lut_LC_12_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i26_3_lut_LC_12_28_5 .LUT_INIT=16'b0000001111001100;
    LogicCell40 \c0.tx.i26_3_lut_LC_12_28_5  (
            .in0(_gnd_net_),
            .in1(N__29199),
            .in2(N__29124),
            .in3(N__29117),
            .lcout(),
            .ltout(\c0.tx.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_12_28_6 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_12_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_12_28_6 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_12_28_6  (
            .in0(_gnd_net_),
            .in1(N__28868),
            .in2(N__29025),
            .in3(N__28979),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37615),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i78_LC_13_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i78_LC_13_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i78_LC_13_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i78_LC_13_18_0  (
            .in0(N__35880),
            .in1(N__28841),
            .in2(_gnd_net_),
            .in3(N__28816),
            .lcout(data_in_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37553),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i49_LC_13_18_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i49_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i49_LC_13_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i49_LC_13_18_4  (
            .in0(N__35879),
            .in1(N__31031),
            .in2(_gnd_net_),
            .in3(N__28781),
            .lcout(data_in_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37553),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i77_LC_13_18_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i77_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i77_LC_13_18_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i77_LC_13_18_5  (
            .in0(N__35899),
            .in1(N__30367),
            .in2(_gnd_net_),
            .in3(N__30419),
            .lcout(data_in_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37553),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i125_LC_13_19_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i125_LC_13_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i125_LC_13_19_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i125_LC_13_19_0  (
            .in0(N__30307),
            .in1(N__35980),
            .in2(_gnd_net_),
            .in3(N__30341),
            .lcout(data_in_15_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i109_LC_13_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i109_LC_13_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i109_LC_13_19_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i109_LC_13_19_1  (
            .in0(N__33074),
            .in1(N__32133),
            .in2(N__30290),
            .in3(N__30250),
            .lcout(\c0.data_in_field_108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i71_LC_13_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i71_LC_13_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i71_LC_13_19_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i71_LC_13_19_2  (
            .in0(N__29484),
            .in1(N__33076),
            .in2(N__31169),
            .in3(N__32232),
            .lcout(\c0.data_in_field_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5997_bdd_4_lut_LC_13_19_3 .C_ON=1'b0;
    defparam \c0.n5997_bdd_4_lut_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.n5997_bdd_4_lut_LC_13_19_3 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.n5997_bdd_4_lut_LC_13_19_3  (
            .in0(N__30210),
            .in1(N__31411),
            .in2(N__29625),
            .in3(N__29586),
            .lcout(\c0.n6000 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i57_LC_13_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i57_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i57_LC_13_19_4 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0___i57_LC_13_19_4  (
            .in0(N__29459),
            .in1(N__33075),
            .in2(N__31032),
            .in3(N__32231),
            .lcout(\c0.data_in_field_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_880_LC_13_19_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_880_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_880_LC_13_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_880_LC_13_19_5  (
            .in0(N__29535),
            .in1(N__29483),
            .in2(_gnd_net_),
            .in3(N__29458),
            .lcout(\c0.n5494 ),
            .ltout(\c0.n5494_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_884_LC_13_19_6 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_884_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_884_LC_13_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_884_LC_13_19_6  (
            .in0(N__29429),
            .in1(N__29412),
            .in2(N__29385),
            .in3(N__29378),
            .lcout(\c0.n26_adj_1927 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i57_LC_13_19_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i57_LC_13_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i57_LC_13_19_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i57_LC_13_19_7  (
            .in0(N__35979),
            .in1(N__31027),
            .in2(_gnd_net_),
            .in3(N__31058),
            .lcout(data_in_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37563),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_888_LC_13_20_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_888_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_888_LC_13_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_888_LC_13_20_0  (
            .in0(N__31013),
            .in1(N__30974),
            .in2(N__30936),
            .in3(N__30489),
            .lcout(\c0.n25_adj_1931 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_965_LC_13_20_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_965_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_965_LC_13_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_965_LC_13_20_2  (
            .in0(N__31400),
            .in1(N__30897),
            .in2(N__30846),
            .in3(N__30780),
            .lcout(\c0.n5542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i137_LC_13_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i137_LC_13_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i137_LC_13_20_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i137_LC_13_20_3  (
            .in0(N__33153),
            .in1(N__32134),
            .in2(N__30705),
            .in3(N__30568),
            .lcout(\c0.data_in_field_136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i83_LC_13_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i83_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i83_LC_13_20_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i83_LC_13_20_6  (
            .in0(N__36074),
            .in1(N__31253),
            .in2(_gnd_net_),
            .in3(N__30658),
            .lcout(data_in_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i39_LC_13_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i39_LC_13_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i39_LC_13_20_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0___i39_LC_13_20_7  (
            .in0(N__33154),
            .in1(N__32135),
            .in2(N__30642),
            .in3(N__30605),
            .lcout(\c0.data_in_field_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37573),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i7_LC_13_21_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i7_LC_13_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i7_LC_13_21_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.byte_transmit_counter__i7_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__33466),
            .in2(_gnd_net_),
            .in3(N__33306),
            .lcout(\c0.byte_transmit_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_941_LC_13_21_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_941_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_941_LC_13_21_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_941_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__30560),
            .in2(_gnd_net_),
            .in3(N__30530),
            .lcout(\c0.n2113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i81_LC_13_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i81_LC_13_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i81_LC_13_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i81_LC_13_21_4  (
            .in0(N__36015),
            .in1(N__30482),
            .in2(_gnd_net_),
            .in3(N__30439),
            .lcout(data_in_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i40_LC_13_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i40_LC_13_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i40_LC_13_21_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0___i40_LC_13_21_5  (
            .in0(N__32989),
            .in1(N__32169),
            .in2(N__31412),
            .in3(N__31436),
            .lcout(\c0.data_in_field_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i80_LC_13_21_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i80_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i80_LC_13_21_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i80_LC_13_21_6  (
            .in0(N__36014),
            .in1(N__31322),
            .in2(_gnd_net_),
            .in3(N__31368),
            .lcout(data_in_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i110_LC_13_21_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i110_LC_13_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i110_LC_13_21_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i110_LC_13_21_7  (
            .in0(N__35900),
            .in1(N__31310),
            .in2(_gnd_net_),
            .in3(N__34477),
            .lcout(data_in_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37580),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i91_LC_13_22_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i91_LC_13_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i91_LC_13_22_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i91_LC_13_22_0  (
            .in0(N__36058),
            .in1(N__31246),
            .in2(_gnd_net_),
            .in3(N__31276),
            .lcout(data_in_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i29_LC_13_22_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i29_LC_13_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i29_LC_13_22_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i29_LC_13_22_2  (
            .in0(N__36057),
            .in1(N__31223),
            .in2(_gnd_net_),
            .in3(N__31125),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i71_LC_13_22_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i71_LC_13_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i71_LC_13_22_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i71_LC_13_22_3  (
            .in0(N__36062),
            .in1(N__31197),
            .in2(_gnd_net_),
            .in3(N__31153),
            .lcout(data_in_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i21_LC_13_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i21_LC_13_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i21_LC_13_22_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i21_LC_13_22_4  (
            .in0(N__36056),
            .in1(N__31089),
            .in2(_gnd_net_),
            .in3(N__31126),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37587),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i0_LC_13_23_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter__i0_LC_13_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i0_LC_13_23_0 .LUT_INIT=16'b1001011000000000;
    LogicCell40 \c0.byte_transmit_counter__i0_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__31068),
            .in2(N__34278),
            .in3(N__37734),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\c0.n4703 ),
            .clk(N__37595),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i1_LC_13_23_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter__i1_LC_13_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i1_LC_13_23_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.byte_transmit_counter__i1_LC_13_23_1  (
            .in0(N__37735),
            .in1(N__34017),
            .in2(_gnd_net_),
            .in3(N__33375),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(\c0.n4703 ),
            .carryout(\c0.n4704 ),
            .clk(N__37595),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_4_lut_LC_13_23_2 .C_ON=1'b1;
    defparam \c0.add_1824_4_lut_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_4_lut_LC_13_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_4_lut_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__34108),
            .in2(_gnd_net_),
            .in3(N__33372),
            .lcout(\c0.tx_transmit_N_568_2 ),
            .ltout(),
            .carryin(\c0.n4704 ),
            .carryout(\c0.n4705 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_5_lut_LC_13_23_3 .C_ON=1'b1;
    defparam \c0.add_1824_5_lut_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_5_lut_LC_13_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_5_lut_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34187),
            .in3(N__33369),
            .lcout(\c0.tx_transmit_N_568_3 ),
            .ltout(),
            .carryin(\c0.n4705 ),
            .carryout(\c0.n4706 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_6_lut_LC_13_23_4 .C_ON=1'b1;
    defparam \c0.add_1824_6_lut_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_6_lut_LC_13_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_6_lut_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__33713),
            .in2(_gnd_net_),
            .in3(N__33366),
            .lcout(\c0.tx_transmit_N_568_4 ),
            .ltout(),
            .carryin(\c0.n4706 ),
            .carryout(\c0.n4707 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_7_lut_LC_13_23_5 .C_ON=1'b1;
    defparam \c0.add_1824_7_lut_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_7_lut_LC_13_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_7_lut_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__33363),
            .in2(_gnd_net_),
            .in3(N__33348),
            .lcout(\c0.tx_transmit_N_568_5 ),
            .ltout(),
            .carryin(\c0.n4707 ),
            .carryout(\c0.n4708 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_8_lut_LC_13_23_6 .C_ON=1'b1;
    defparam \c0.add_1824_8_lut_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_8_lut_LC_13_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_1824_8_lut_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__33345),
            .in2(_gnd_net_),
            .in3(N__33321),
            .lcout(\c0.tx_transmit_N_568_6 ),
            .ltout(),
            .carryin(\c0.n4708 ),
            .carryout(\c0.n4709 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_1824_9_lut_LC_13_23_7 .C_ON=1'b0;
    defparam \c0.add_1824_9_lut_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_1824_9_lut_LC_13_23_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.add_1824_9_lut_LC_13_23_7  (
            .in0(N__33318),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33309),
            .lcout(\c0.tx_transmit_N_568_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i3_LC_13_24_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i3_LC_13_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i3_LC_13_24_0 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \c0.byte_transmit_counter__i3_LC_13_24_0  (
            .in0(N__33291),
            .in1(N__33436),
            .in2(N__33471),
            .in3(N__33492),
            .lcout(\c0.byte_transmit_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_842_LC_13_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_842_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_842_LC_13_24_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_842_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__33416),
            .in2(_gnd_net_),
            .in3(N__33290),
            .lcout(\c0.n95 ),
            .ltout(\c0.n95_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i120_2_lut_LC_13_24_2 .C_ON=1'b0;
    defparam \c0.i120_2_lut_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i120_2_lut_LC_13_24_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i120_2_lut_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33528),
            .in3(N__33432),
            .lcout(\c0.n106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_995_LC_13_24_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_995_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_995_LC_13_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_995_LC_13_24_3  (
            .in0(N__34533),
            .in1(N__33664),
            .in2(N__34383),
            .in3(N__36120),
            .lcout(n4_adj_1981),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_13_24_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_13_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_13_24_4  (
            .in0(N__36175),
            .in1(N__36641),
            .in2(_gnd_net_),
            .in3(N__34650),
            .lcout(n7_adj_1988),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i2_LC_13_24_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i2_LC_13_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i2_LC_13_24_5 .LUT_INIT=16'b1100110100000000;
    LogicCell40 \c0.byte_transmit_counter__i2_LC_13_24_5  (
            .in0(N__33491),
            .in1(N__33467),
            .in2(N__33438),
            .in3(N__33417),
            .lcout(\c0.byte_transmit_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i13_LC_13_24_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i13_LC_13_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i13_LC_13_24_7 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i13_LC_13_24_7  (
            .in0(N__34962),
            .in1(N__36892),
            .in2(N__37110),
            .in3(N__36752),
            .lcout(data_out_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37601),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_13_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_13_25_0 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i31_4_lut_LC_13_25_0  (
            .in0(N__33381),
            .in1(N__33723),
            .in2(N__33408),
            .in3(N__34116),
            .lcout(tx_data_5_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1000_LC_13_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1000_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1000_LC_13_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1000_LC_13_25_1  (
            .in0(N__33656),
            .in1(N__36173),
            .in2(_gnd_net_),
            .in3(N__34375),
            .lcout(n5424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i35_3_lut_LC_13_25_2 .C_ON=1'b0;
    defparam \c0.i35_3_lut_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i35_3_lut_LC_13_25_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i35_3_lut_LC_13_25_2  (
            .in0(N__34649),
            .in1(N__36119),
            .in2(_gnd_net_),
            .in3(N__34302),
            .lcout(\c0.n31_adj_1912 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i748_4_lut_LC_13_25_3 .C_ON=1'b0;
    defparam \c0.i748_4_lut_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i748_4_lut_LC_13_25_3 .LUT_INIT=16'b1101000100100010;
    LogicCell40 \c0.i748_4_lut_LC_13_25_3  (
            .in0(N__34303),
            .in1(N__34173),
            .in2(N__34395),
            .in3(N__34058),
            .lcout(\c0.n989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_13_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_13_25_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i9_3_lut_LC_13_25_4  (
            .in0(N__34945),
            .in1(N__33655),
            .in2(_gnd_net_),
            .in3(N__34301),
            .lcout(),
            .ltout(\c0.n9_adj_1906_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i15_4_lut_LC_13_25_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i15_4_lut_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i15_4_lut_LC_13_25_5 .LUT_INIT=16'b1100100001110111;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i15_4_lut_LC_13_25_5  (
            .in0(N__34115),
            .in1(N__34172),
            .in2(N__33681),
            .in3(N__34057),
            .lcout(\c0.n15_adj_1909 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i951_2_lut_LC_13_25_6 .C_ON=1'b0;
    defparam \c0.i951_2_lut_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i951_2_lut_LC_13_25_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i951_2_lut_LC_13_25_6  (
            .in0(N__34171),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34114),
            .lcout(\c0.n1251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i5_LC_13_25_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i5_LC_13_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i5_LC_13_25_7 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i5_LC_13_25_7  (
            .in0(N__33657),
            .in1(N__36897),
            .in2(N__37866),
            .in3(N__36748),
            .lcout(data_out_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37607),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2044_4_lut_LC_13_26_1 .C_ON=1'b0;
    defparam \c0.i2044_4_lut_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2044_4_lut_LC_13_26_1 .LUT_INIT=16'b1100000010111011;
    LogicCell40 \c0.i2044_4_lut_LC_13_26_1  (
            .in0(N__36169),
            .in1(N__34197),
            .in2(N__36964),
            .in3(N__34320),
            .lcout(\c0.n2293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i16_LC_13_26_2 .C_ON=1'b0;
    defparam \c0.data_out_0___i16_LC_13_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i16_LC_13_26_2 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i16_LC_13_26_2  (
            .in0(N__34521),
            .in1(N__36898),
            .in2(N__37044),
            .in3(N__36783),
            .lcout(data_out_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37611),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_933_LC_13_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_933_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_933_LC_13_26_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_933_LC_13_26_3  (
            .in0(N__34695),
            .in1(N__34518),
            .in2(N__34969),
            .in3(N__36111),
            .lcout(n5479),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_844_LC_13_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_844_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_844_LC_13_26_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_844_LC_13_26_4  (
            .in0(N__34520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36499),
            .lcout(n4_adj_1996),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_13_26_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_13_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_13_26_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_13_26_6  (
            .in0(N__33609),
            .in1(N__33906),
            .in2(_gnd_net_),
            .in3(N__33534),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37611),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1005_LC_13_26_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1005_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1005_LC_13_26_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1005_LC_13_26_7  (
            .in0(N__34696),
            .in1(N__34519),
            .in2(N__34968),
            .in3(N__36112),
            .lcout(n5421),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i8_LC_13_27_0 .C_ON=1'b0;
    defparam \c0.data_out_0___i8_LC_13_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i8_LC_13_27_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.data_out_0___i8_LC_13_27_0  (
            .in0(N__36785),
            .in1(N__37791),
            .in2(N__36500),
            .in3(N__36894),
            .lcout(data_out_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37616),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5595_4_lut_LC_13_27_1 .C_ON=1'b0;
    defparam \c0.i5595_4_lut_LC_13_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5595_4_lut_LC_13_27_1 .LUT_INIT=16'b1111001110111011;
    LogicCell40 \c0.i5595_4_lut_LC_13_27_1  (
            .in0(N__33951),
            .in1(N__34060),
            .in2(N__36348),
            .in3(N__34322),
            .lcout(\c0.n5845 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i4_LC_13_27_2 .C_ON=1'b0;
    defparam \c0.data_out_0___i4_LC_13_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i4_LC_13_27_2 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0___i4_LC_13_27_2  (
            .in0(N__36784),
            .in1(N__36639),
            .in2(N__37887),
            .in3(N__36893),
            .lcout(data_out_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37616),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5582_4_lut_LC_13_27_3 .C_ON=1'b0;
    defparam \c0.i5582_4_lut_LC_13_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5582_4_lut_LC_13_27_3 .LUT_INIT=16'b1111001110111011;
    LogicCell40 \c0.i5582_4_lut_LC_13_27_3  (
            .in0(N__37641),
            .in1(N__34059),
            .in2(N__33936),
            .in3(N__34321),
            .lcout(\c0.n5837 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.n6285_bdd_4_lut_LC_13_27_4 .C_ON=1'b0;
    defparam \c0.tx.n6285_bdd_4_lut_LC_13_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.n6285_bdd_4_lut_LC_13_27_4 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.tx.n6285_bdd_4_lut_LC_13_27_4  (
            .in0(N__33905),
            .in1(N__33883),
            .in2(N__33834),
            .in3(N__33816),
            .lcout(\c0.tx.n6288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i9_LC_13_27_6 .C_ON=1'b0;
    defparam \c0.data_out_0___i9_LC_13_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i9_LC_13_27_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0___i9_LC_13_27_6  (
            .in0(N__36786),
            .in1(N__36550),
            .in2(N__36327),
            .in3(N__36895),
            .lcout(data_out_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37616),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_897_LC_13_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_897_LC_13_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_897_LC_13_28_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_897_LC_13_28_1  (
            .in0(N__34706),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36109),
            .lcout(n5415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_13_28_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_13_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_13_28_4 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i31_4_lut_LC_13_28_4  (
            .in0(N__33984),
            .in1(N__33783),
            .in2(N__33753),
            .in3(N__33744),
            .lcout(tx_data_1_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_937_LC_13_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_937_LC_13_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_937_LC_13_28_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_937_LC_13_28_5  (
            .in0(N__34705),
            .in1(N__36108),
            .in2(_gnd_net_),
            .in3(N__34532),
            .lcout(n1579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i102_LC_14_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i102_LC_14_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i102_LC_14_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i102_LC_14_21_4  (
            .in0(N__35999),
            .in1(N__34478),
            .in2(_gnd_net_),
            .in3(N__34444),
            .lcout(data_in_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37588),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i6_LC_14_23_0 .C_ON=1'b0;
    defparam \c0.data_out_0___i6_LC_14_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i6_LC_14_23_0 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i6_LC_14_23_0  (
            .in0(N__34419),
            .in1(N__36900),
            .in2(N__37842),
            .in3(N__36791),
            .lcout(data_out_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37602),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_14_23_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_14_23_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i9_3_lut_LC_14_23_6  (
            .in0(N__34682),
            .in1(N__34411),
            .in2(_gnd_net_),
            .in3(N__34269),
            .lcout(\c0.n9_adj_1911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i1_LC_14_24_0 .C_ON=1'b0;
    defparam \c0.data_out_0___i1_LC_14_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i1_LC_14_24_0 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.data_out_0___i1_LC_14_24_0  (
            .in0(N__34379),
            .in1(N__37023),
            .in2(N__36912),
            .in3(N__36769),
            .lcout(data_out_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37608),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_14_24_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_14_24_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i9_3_lut_LC_14_24_1  (
            .in0(N__35014),
            .in1(N__36666),
            .in2(_gnd_net_),
            .in3(N__34270),
            .lcout(),
            .ltout(\c0.n9_adj_1891_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_LC_14_24_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_LC_14_24_2 .LUT_INIT=16'b0110010010011001;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i15_4_lut_LC_14_24_2  (
            .in0(N__34186),
            .in1(N__34117),
            .in2(N__34083),
            .in3(N__34036),
            .lcout(\c0.n15_adj_1893 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i7_LC_14_24_4 .C_ON=1'b0;
    defparam \c0.data_out_0___i7_LC_14_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i7_LC_14_24_4 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i7_LC_14_24_4  (
            .in0(N__34642),
            .in1(N__36902),
            .in2(N__37818),
            .in3(N__36771),
            .lcout(data_out_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37608),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i2_LC_14_24_5 .C_ON=1'b0;
    defparam \c0.data_out_0___i2_LC_14_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i2_LC_14_24_5 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \c0.data_out_0___i2_LC_14_24_5  (
            .in0(N__36770),
            .in1(N__37005),
            .in2(N__36911),
            .in3(N__36667),
            .lcout(data_out_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37608),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i14_LC_14_24_6 .C_ON=1'b0;
    defparam \c0.data_out_0___i14_LC_14_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i14_LC_14_24_6 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i14_LC_14_24_6  (
            .in0(N__34694),
            .in1(N__36901),
            .in2(N__37086),
            .in3(N__36768),
            .lcout(data_out_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37608),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_959_LC_14_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_959_LC_14_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_959_LC_14_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_959_LC_14_24_7  (
            .in0(N__36174),
            .in1(N__34641),
            .in2(_gnd_net_),
            .in3(N__36566),
            .lcout(n4_adj_1976),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i0_LC_14_25_0.C_ON=1'b1;
    defparam blink_counter_523__i0_LC_14_25_0.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i0_LC_14_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i0_LC_14_25_0 (
            .in0(_gnd_net_),
            .in1(N__34593),
            .in2(_gnd_net_),
            .in3(N__34587),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(n4710),
            .clk(N__37612),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i1_LC_14_25_1.C_ON=1'b1;
    defparam blink_counter_523__i1_LC_14_25_1.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i1_LC_14_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i1_LC_14_25_1 (
            .in0(_gnd_net_),
            .in1(N__34584),
            .in2(_gnd_net_),
            .in3(N__34578),
            .lcout(n25),
            .ltout(),
            .carryin(n4710),
            .carryout(n4711),
            .clk(N__37612),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i2_LC_14_25_2.C_ON=1'b1;
    defparam blink_counter_523__i2_LC_14_25_2.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i2_LC_14_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i2_LC_14_25_2 (
            .in0(_gnd_net_),
            .in1(N__34575),
            .in2(_gnd_net_),
            .in3(N__34569),
            .lcout(n24),
            .ltout(),
            .carryin(n4711),
            .carryout(n4712),
            .clk(N__37612),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i3_LC_14_25_3.C_ON=1'b1;
    defparam blink_counter_523__i3_LC_14_25_3.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i3_LC_14_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i3_LC_14_25_3 (
            .in0(_gnd_net_),
            .in1(N__34566),
            .in2(_gnd_net_),
            .in3(N__34560),
            .lcout(n23),
            .ltout(),
            .carryin(n4712),
            .carryout(n4713),
            .clk(N__37612),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i4_LC_14_25_4.C_ON=1'b1;
    defparam blink_counter_523__i4_LC_14_25_4.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i4_LC_14_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i4_LC_14_25_4 (
            .in0(_gnd_net_),
            .in1(N__34557),
            .in2(_gnd_net_),
            .in3(N__34551),
            .lcout(n22),
            .ltout(),
            .carryin(n4713),
            .carryout(n4714),
            .clk(N__37612),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i5_LC_14_25_5.C_ON=1'b1;
    defparam blink_counter_523__i5_LC_14_25_5.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i5_LC_14_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i5_LC_14_25_5 (
            .in0(_gnd_net_),
            .in1(N__34548),
            .in2(_gnd_net_),
            .in3(N__34542),
            .lcout(n21),
            .ltout(),
            .carryin(n4714),
            .carryout(n4715),
            .clk(N__37612),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i6_LC_14_25_6.C_ON=1'b1;
    defparam blink_counter_523__i6_LC_14_25_6.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i6_LC_14_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i6_LC_14_25_6 (
            .in0(_gnd_net_),
            .in1(N__34539),
            .in2(_gnd_net_),
            .in3(N__34782),
            .lcout(n20),
            .ltout(),
            .carryin(n4715),
            .carryout(n4716),
            .clk(N__37612),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i7_LC_14_25_7.C_ON=1'b1;
    defparam blink_counter_523__i7_LC_14_25_7.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i7_LC_14_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i7_LC_14_25_7 (
            .in0(_gnd_net_),
            .in1(N__34779),
            .in2(_gnd_net_),
            .in3(N__34773),
            .lcout(n19),
            .ltout(),
            .carryin(n4716),
            .carryout(n4717),
            .clk(N__37612),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i8_LC_14_26_0.C_ON=1'b1;
    defparam blink_counter_523__i8_LC_14_26_0.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i8_LC_14_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i8_LC_14_26_0 (
            .in0(_gnd_net_),
            .in1(N__34770),
            .in2(_gnd_net_),
            .in3(N__34764),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(n4718),
            .clk(N__37617),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i9_LC_14_26_1.C_ON=1'b1;
    defparam blink_counter_523__i9_LC_14_26_1.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i9_LC_14_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i9_LC_14_26_1 (
            .in0(_gnd_net_),
            .in1(N__34761),
            .in2(_gnd_net_),
            .in3(N__34755),
            .lcout(n17),
            .ltout(),
            .carryin(n4718),
            .carryout(n4719),
            .clk(N__37617),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i10_LC_14_26_2.C_ON=1'b1;
    defparam blink_counter_523__i10_LC_14_26_2.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i10_LC_14_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i10_LC_14_26_2 (
            .in0(_gnd_net_),
            .in1(N__34752),
            .in2(_gnd_net_),
            .in3(N__34746),
            .lcout(n16),
            .ltout(),
            .carryin(n4719),
            .carryout(n4720),
            .clk(N__37617),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i11_LC_14_26_3.C_ON=1'b1;
    defparam blink_counter_523__i11_LC_14_26_3.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i11_LC_14_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i11_LC_14_26_3 (
            .in0(_gnd_net_),
            .in1(N__34743),
            .in2(_gnd_net_),
            .in3(N__34737),
            .lcout(n15),
            .ltout(),
            .carryin(n4720),
            .carryout(n4721),
            .clk(N__37617),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i12_LC_14_26_4.C_ON=1'b1;
    defparam blink_counter_523__i12_LC_14_26_4.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i12_LC_14_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i12_LC_14_26_4 (
            .in0(_gnd_net_),
            .in1(N__34734),
            .in2(_gnd_net_),
            .in3(N__34728),
            .lcout(n14),
            .ltout(),
            .carryin(n4721),
            .carryout(n4722),
            .clk(N__37617),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i13_LC_14_26_5.C_ON=1'b1;
    defparam blink_counter_523__i13_LC_14_26_5.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i13_LC_14_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i13_LC_14_26_5 (
            .in0(_gnd_net_),
            .in1(N__34725),
            .in2(_gnd_net_),
            .in3(N__34719),
            .lcout(n13),
            .ltout(),
            .carryin(n4722),
            .carryout(n4723),
            .clk(N__37617),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i14_LC_14_26_6.C_ON=1'b1;
    defparam blink_counter_523__i14_LC_14_26_6.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i14_LC_14_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i14_LC_14_26_6 (
            .in0(_gnd_net_),
            .in1(N__34716),
            .in2(_gnd_net_),
            .in3(N__34710),
            .lcout(n12),
            .ltout(),
            .carryin(n4723),
            .carryout(n4724),
            .clk(N__37617),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i15_LC_14_26_7.C_ON=1'b1;
    defparam blink_counter_523__i15_LC_14_26_7.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i15_LC_14_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i15_LC_14_26_7 (
            .in0(_gnd_net_),
            .in1(N__34890),
            .in2(_gnd_net_),
            .in3(N__34884),
            .lcout(n11),
            .ltout(),
            .carryin(n4724),
            .carryout(n4725),
            .clk(N__37617),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i16_LC_14_27_0.C_ON=1'b1;
    defparam blink_counter_523__i16_LC_14_27_0.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i16_LC_14_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i16_LC_14_27_0 (
            .in0(_gnd_net_),
            .in1(N__34881),
            .in2(_gnd_net_),
            .in3(N__34875),
            .lcout(n10),
            .ltout(),
            .carryin(bfn_14_27_0_),
            .carryout(n4726),
            .clk(N__37619),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i17_LC_14_27_1.C_ON=1'b1;
    defparam blink_counter_523__i17_LC_14_27_1.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i17_LC_14_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i17_LC_14_27_1 (
            .in0(_gnd_net_),
            .in1(N__34872),
            .in2(_gnd_net_),
            .in3(N__34866),
            .lcout(n9),
            .ltout(),
            .carryin(n4726),
            .carryout(n4727),
            .clk(N__37619),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i18_LC_14_27_2.C_ON=1'b1;
    defparam blink_counter_523__i18_LC_14_27_2.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i18_LC_14_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i18_LC_14_27_2 (
            .in0(_gnd_net_),
            .in1(N__34863),
            .in2(_gnd_net_),
            .in3(N__34857),
            .lcout(n8),
            .ltout(),
            .carryin(n4727),
            .carryout(n4728),
            .clk(N__37619),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i19_LC_14_27_3.C_ON=1'b1;
    defparam blink_counter_523__i19_LC_14_27_3.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i19_LC_14_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i19_LC_14_27_3 (
            .in0(_gnd_net_),
            .in1(N__34854),
            .in2(_gnd_net_),
            .in3(N__34848),
            .lcout(n7),
            .ltout(),
            .carryin(n4728),
            .carryout(n4729),
            .clk(N__37619),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i20_LC_14_27_4.C_ON=1'b1;
    defparam blink_counter_523__i20_LC_14_27_4.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i20_LC_14_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i20_LC_14_27_4 (
            .in0(_gnd_net_),
            .in1(N__34845),
            .in2(_gnd_net_),
            .in3(N__34839),
            .lcout(n6),
            .ltout(),
            .carryin(n4729),
            .carryout(n4730),
            .clk(N__37619),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i21_LC_14_27_5.C_ON=1'b1;
    defparam blink_counter_523__i21_LC_14_27_5.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i21_LC_14_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i21_LC_14_27_5 (
            .in0(_gnd_net_),
            .in1(N__34823),
            .in2(_gnd_net_),
            .in3(N__34812),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n4730),
            .carryout(n4731),
            .clk(N__37619),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i22_LC_14_27_6.C_ON=1'b1;
    defparam blink_counter_523__i22_LC_14_27_6.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i22_LC_14_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i22_LC_14_27_6 (
            .in0(_gnd_net_),
            .in1(N__34796),
            .in2(_gnd_net_),
            .in3(N__34785),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n4731),
            .carryout(n4732),
            .clk(N__37619),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i23_LC_14_27_7.C_ON=1'b1;
    defparam blink_counter_523__i23_LC_14_27_7.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i23_LC_14_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i23_LC_14_27_7 (
            .in0(_gnd_net_),
            .in1(N__36248),
            .in2(_gnd_net_),
            .in3(N__36237),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n4732),
            .carryout(n4733),
            .clk(N__37619),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i24_LC_14_28_0.C_ON=1'b1;
    defparam blink_counter_523__i24_LC_14_28_0.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i24_LC_14_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i24_LC_14_28_0 (
            .in0(_gnd_net_),
            .in1(N__36221),
            .in2(_gnd_net_),
            .in3(N__36210),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_14_28_0_),
            .carryout(n4734),
            .clk(N__37621),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_523__i25_LC_14_28_1.C_ON=1'b0;
    defparam blink_counter_523__i25_LC_14_28_1.SEQ_MODE=4'b1000;
    defparam blink_counter_523__i25_LC_14_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_523__i25_LC_14_28_1 (
            .in0(_gnd_net_),
            .in1(N__36194),
            .in2(_gnd_net_),
            .in3(N__36207),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37621),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i3_LC_14_28_6 .C_ON=1'b0;
    defparam \c0.data_out_0___i3_LC_14_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i3_LC_14_28_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_out_0___i3_LC_14_28_6  (
            .in0(N__36788),
            .in1(N__36150),
            .in2(N__36984),
            .in3(N__36896),
            .lcout(data_out_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37621),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i15_LC_14_28_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i15_LC_14_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i15_LC_14_28_7 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_out_0___i15_LC_14_28_7  (
            .in0(N__36110),
            .in1(N__36787),
            .in2(N__37065),
            .in3(N__36899),
            .lcout(data_out_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37621),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i121_LC_15_21_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i121_LC_15_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i121_LC_15_21_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i121_LC_15_21_3  (
            .in0(N__36000),
            .in1(N__35051),
            .in2(_gnd_net_),
            .in3(N__35099),
            .lcout(data_in_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37596),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_978_LC_15_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_978_LC_15_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_978_LC_15_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_978_LC_15_24_0  (
            .in0(N__36935),
            .in1(N__36390),
            .in2(_gnd_net_),
            .in3(N__36565),
            .lcout(\c0.n5409 ),
            .ltout(\c0.n5409_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_15_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_15_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_15_24_1  (
            .in0(N__36507),
            .in1(N__35019),
            .in2(N__34974),
            .in3(N__34961),
            .lcout(n4_adj_1978),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_990_LC_15_24_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_990_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_990_LC_15_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_990_LC_15_24_4  (
            .in0(N__36682),
            .in1(N__36391),
            .in2(_gnd_net_),
            .in3(N__36640),
            .lcout(n4_adj_1983),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i11_LC_15_24_5 .C_ON=1'b0;
    defparam \c0.data_out_0___i11_LC_15_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i11_LC_15_24_5 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i11_LC_15_24_5  (
            .in0(N__36945),
            .in1(N__36909),
            .in2(N__36282),
            .in3(N__36789),
            .lcout(data_out_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37613),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i12_LC_15_24_7 .C_ON=1'b0;
    defparam \c0.data_out_0___i12_LC_15_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i12_LC_15_24_7 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \c0.data_out_0___i12_LC_15_24_7  (
            .in0(N__36392),
            .in1(N__36910),
            .in2(N__37131),
            .in3(N__36790),
            .lcout(data_out_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37613),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_LC_15_25_2 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_LC_15_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_LC_15_25_2  (
            .in0(N__36680),
            .in1(N__36642),
            .in2(N__36587),
            .in3(N__36567),
            .lcout(n8_adj_1984),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_981_LC_15_25_4 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_981_LC_15_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_981_LC_15_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_981_LC_15_25_4  (
            .in0(N__36506),
            .in1(N__36441),
            .in2(_gnd_net_),
            .in3(N__36399),
            .lcout(),
            .ltout(n7_adj_1985_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i26_LC_15_25_5 .C_ON=1'b0;
    defparam \c0.data_out_0___i26_LC_15_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i26_LC_15_25_5 .LUT_INIT=16'b1010101011000011;
    LogicCell40 \c0.data_out_0___i26_LC_15_25_5  (
            .in0(N__36341),
            .in1(N__36357),
            .in2(N__36351),
            .in3(N__37736),
            .lcout(data_out_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37618),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i0_LC_15_26_0 .C_ON=1'b1;
    defparam \c0.data_527__i0_LC_15_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i0_LC_15_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i0_LC_15_26_0  (
            .in0(_gnd_net_),
            .in1(N__36317),
            .in2(_gnd_net_),
            .in3(N__36306),
            .lcout(data_0),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(\c0.n4739 ),
            .clk(N__37620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i1_LC_15_26_1 .C_ON=1'b1;
    defparam \c0.data_527__i1_LC_15_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i1_LC_15_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i1_LC_15_26_1  (
            .in0(_gnd_net_),
            .in1(N__36296),
            .in2(_gnd_net_),
            .in3(N__36285),
            .lcout(data_1),
            .ltout(),
            .carryin(\c0.n4739 ),
            .carryout(\c0.n4740 ),
            .clk(N__37620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i2_LC_15_26_2 .C_ON=1'b1;
    defparam \c0.data_527__i2_LC_15_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i2_LC_15_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i2_LC_15_26_2  (
            .in0(_gnd_net_),
            .in1(N__36275),
            .in2(_gnd_net_),
            .in3(N__36264),
            .lcout(data_2),
            .ltout(),
            .carryin(\c0.n4740 ),
            .carryout(\c0.n4741 ),
            .clk(N__37620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i3_LC_15_26_3 .C_ON=1'b1;
    defparam \c0.data_527__i3_LC_15_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i3_LC_15_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i3_LC_15_26_3  (
            .in0(_gnd_net_),
            .in1(N__37124),
            .in2(_gnd_net_),
            .in3(N__37113),
            .lcout(data_3),
            .ltout(),
            .carryin(\c0.n4741 ),
            .carryout(\c0.n4742 ),
            .clk(N__37620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i4_LC_15_26_4 .C_ON=1'b1;
    defparam \c0.data_527__i4_LC_15_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i4_LC_15_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i4_LC_15_26_4  (
            .in0(_gnd_net_),
            .in1(N__37100),
            .in2(_gnd_net_),
            .in3(N__37089),
            .lcout(data_4),
            .ltout(),
            .carryin(\c0.n4742 ),
            .carryout(\c0.n4743 ),
            .clk(N__37620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i5_LC_15_26_5 .C_ON=1'b1;
    defparam \c0.data_527__i5_LC_15_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i5_LC_15_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i5_LC_15_26_5  (
            .in0(_gnd_net_),
            .in1(N__37079),
            .in2(_gnd_net_),
            .in3(N__37068),
            .lcout(data_5),
            .ltout(),
            .carryin(\c0.n4743 ),
            .carryout(\c0.n4744 ),
            .clk(N__37620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i6_LC_15_26_6 .C_ON=1'b1;
    defparam \c0.data_527__i6_LC_15_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i6_LC_15_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i6_LC_15_26_6  (
            .in0(_gnd_net_),
            .in1(N__37058),
            .in2(_gnd_net_),
            .in3(N__37047),
            .lcout(data_6),
            .ltout(),
            .carryin(\c0.n4744 ),
            .carryout(\c0.n4745 ),
            .clk(N__37620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i7_LC_15_26_7 .C_ON=1'b1;
    defparam \c0.data_527__i7_LC_15_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i7_LC_15_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i7_LC_15_26_7  (
            .in0(_gnd_net_),
            .in1(N__37037),
            .in2(_gnd_net_),
            .in3(N__37026),
            .lcout(data_7),
            .ltout(),
            .carryin(\c0.n4745 ),
            .carryout(\c0.n4746 ),
            .clk(N__37620),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i8_LC_15_27_0 .C_ON=1'b1;
    defparam \c0.data_527__i8_LC_15_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i8_LC_15_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i8_LC_15_27_0  (
            .in0(_gnd_net_),
            .in1(N__37019),
            .in2(_gnd_net_),
            .in3(N__37008),
            .lcout(data_8),
            .ltout(),
            .carryin(bfn_15_27_0_),
            .carryout(\c0.n4747 ),
            .clk(N__37622),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i9_LC_15_27_1 .C_ON=1'b1;
    defparam \c0.data_527__i9_LC_15_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i9_LC_15_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i9_LC_15_27_1  (
            .in0(_gnd_net_),
            .in1(N__36998),
            .in2(_gnd_net_),
            .in3(N__36987),
            .lcout(data_9),
            .ltout(),
            .carryin(\c0.n4747 ),
            .carryout(\c0.n4748 ),
            .clk(N__37622),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i10_LC_15_27_2 .C_ON=1'b1;
    defparam \c0.data_527__i10_LC_15_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i10_LC_15_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i10_LC_15_27_2  (
            .in0(_gnd_net_),
            .in1(N__36980),
            .in2(_gnd_net_),
            .in3(N__36969),
            .lcout(data_10),
            .ltout(),
            .carryin(\c0.n4748 ),
            .carryout(\c0.n4749 ),
            .clk(N__37622),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i11_LC_15_27_3 .C_ON=1'b1;
    defparam \c0.data_527__i11_LC_15_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i11_LC_15_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i11_LC_15_27_3  (
            .in0(_gnd_net_),
            .in1(N__37880),
            .in2(_gnd_net_),
            .in3(N__37869),
            .lcout(data_11),
            .ltout(),
            .carryin(\c0.n4749 ),
            .carryout(\c0.n4750 ),
            .clk(N__37622),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i12_LC_15_27_4 .C_ON=1'b1;
    defparam \c0.data_527__i12_LC_15_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i12_LC_15_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i12_LC_15_27_4  (
            .in0(_gnd_net_),
            .in1(N__37856),
            .in2(_gnd_net_),
            .in3(N__37845),
            .lcout(data_12),
            .ltout(),
            .carryin(\c0.n4750 ),
            .carryout(\c0.n4751 ),
            .clk(N__37622),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i13_LC_15_27_5 .C_ON=1'b1;
    defparam \c0.data_527__i13_LC_15_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i13_LC_15_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i13_LC_15_27_5  (
            .in0(_gnd_net_),
            .in1(N__37832),
            .in2(_gnd_net_),
            .in3(N__37821),
            .lcout(data_13),
            .ltout(),
            .carryin(\c0.n4751 ),
            .carryout(\c0.n4752 ),
            .clk(N__37622),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i14_LC_15_27_6 .C_ON=1'b1;
    defparam \c0.data_527__i14_LC_15_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i14_LC_15_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i14_LC_15_27_6  (
            .in0(_gnd_net_),
            .in1(N__37808),
            .in2(_gnd_net_),
            .in3(N__37797),
            .lcout(data_14),
            .ltout(),
            .carryin(\c0.n4752 ),
            .carryout(\c0.n4753 ),
            .clk(N__37622),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_527__i15_LC_15_27_7 .C_ON=1'b0;
    defparam \c0.data_527__i15_LC_15_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_527__i15_LC_15_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_527__i15_LC_15_27_7  (
            .in0(_gnd_net_),
            .in1(N__37790),
            .in2(_gnd_net_),
            .in3(N__37794),
            .lcout(data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37622),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0___i20_LC_15_29_6 .C_ON=1'b0;
    defparam \c0.data_out_0___i20_LC_15_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0___i20_LC_15_29_6 .LUT_INIT=16'b1100110010100101;
    LogicCell40 \c0.data_out_0___i20_LC_15_29_6  (
            .in0(N__37776),
            .in1(N__37637),
            .in2(N__37764),
            .in3(N__37737),
            .lcout(data_out_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37623),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
